

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AFl2kw3wjuupeEJWAVRMjvI4n2F9ZwKYCyTdtTbrj99jYEYTJx3fm7Ch7UNHIYnYCZk+hug4a3M6
XIrSFOf3lw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kJIX1i40eaci6RDbcVVzg1fYaa68r2QTZ19EbYvWyiO0MSVCOi3GfcyJJxOR52/mcv4FD0GrKyok
p1d2616K9ikEjuEHDsOkFkQxSSfEgbSNAEkwJoywFb1NEza/LgnXq4wCMserYGd0Ho12V4osIEdI
exWoz7u39lGc9ZiaBS4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2kMqoMFPLn7FsBBTsV6uCri7uN+peyfxKN5B0t+cAsrbL+lDiZoUrv6niJBSapyempvdNVVmTzxI
0OOKA0SUZL7oQT5S7r5QAMg9q0wHtWdtsxsKxFyZXOcUUs3IkLwLNJ9fExPXmVlCDUNWWyZ/Qtik
1q9ZynUcX4DCv1pUeRs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uW1nShxn5xYxSfsiNvMbC6cL7GFjn45B3GrJxFfTPdqHxW6l/7kPGVqMN4yc97bwWb5swAmg1/ia
P9L6G5Lmjygww+NIedzfhB4znXCEs1F+LwtP/Eo4UZuH4rQ55XUhLKrRNEqAJ5lTqYxfdIa1JIeg
6YgrU98QHKeOeZUeearBuTROZ6q9d2QFGZhc5MxjU8pwV5JQ++j3EkUIuMZJi3DVdwnYj2d1DzSG
tEt9nWmDzn5rqjvrP0c2GlNBg1tCMJxGfC7y54n+J8H6ETagMe97uL4QvKLTEhjArVfHkKedz6Hw
BLtL2VPOf8fCVrM+AsqxA6SscLteiE3Y/tcuqg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IV462y1jHGYFO6K2VU9zTKlfXJZ4kSNvewSr8uczSbz2qRhu1urkppbYmZyNPMNjUUiJfr+4xl1K
sPX+MN8CN040mI1y/WRE8sMEH4yPflkbYjeDH/AX8AZf0f51eUS3cIc3p5KYvECdG8h6xmZ6jH0F
7BqDcSAL8OaSnIetqzLPr2v1rtYXH+RRlVWmvCK2nFZ02kt8pCYkp8L5RKceyNIKFWCdOT5JdjZY
4tvHtPn6P1gVHsYV30mBGWhvJczj5zrLjwFlzuRt1FBD773q8FliSEnvM5VLjXeYVAshW6krIgcC
JRjJFfG2fLeH0eKFVJ7kqIzwNNYB0nt3Mho0og==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gxKMu2AB/FASbqvyKO7D61/XUsdMsjazR7APgUWhLu8z6ePEw4il1OmWHsQOCjylECfctRxhrNKA
ZkqobGwUpbLybNlM8OLmxSq7gFftkFYAAbUlTfr+gHIvTw0OHQ1EytNPCAXJ3C16VMRZRtIOMhuu
qWzd7JSTNzsFNMOGqUkbAJ25aM5fSFIBT9RqdtK6aDtxz+XRgnizFyeXsqGdP7bY03KX5HgTMa9w
sW64LQcPjQEuBBRxSfYreUKE1jQbO9XuIjtoOmZGDsEtv2KkhTAdFbwHWRiiIzAO+Bx945pksp3X
TfC9rKLaXHs75mi0HkNR/3vshocjTDFwp+bJaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 122928)
`protect data_block
QYoIrrfrQHHs0/IDKowIIOJdF7GDREW8cAkn5W2857GJvsoBifsi+xiQFzb4W/Kb2Rk4AUZeTWM7
2KLzwEVFDhWATiIbnX0qyAdlyuZwIyk+rBaagWYdZWmLy2ZJYIe+f0R100fCo5mFYJ6aXFA+Krvj
W3gObwr56CFZlOZu4h8IGAzKdDmVEbNFfyLF3lB9q5Rlx0TIBCV2ciMApx2MRo3ZmpUf0tF+jtjf
406nvWqFK+nOVgMeqahnehSOJl5LNinmcnkekKd7lrsTEvNkIkNY+JQkFoRox59WGaqn2ttrmpht
Uf8OoRvx3mi9Bh/bdy+8ajyXoWOdC/SLyU2qlvuVAx3AeMzElbp60rYCjKQ34Pol0lv6DXxGdmpH
sne6bzVJJ9cg77sA3X4U4itmZNOkxN1PuKY02TqFfk9gqu9QnwOhFhd0qTQJt+xRkMf2ovwNWQTc
ON8K8E+1iL35gD+LWD5ph2+wAi3UTFOwvHqhGLCqycPgXl9Kx1CVARn3cGAISKVLxsJn8EYczRLZ
CAZllithENvGwt/Yq2e/PqQCVaOgfIZGkH0r4O6Be3R74WgsOzDb2spGbSj3r2Y8NLguKgLOO8Ed
Pacteut9YtLsclRmIjJtS4UhvHiC4T+GDDPVx5yVzU2NCL21IOsLlQUVlr/vOgu9tXZKYslzOICs
Wg1bBwLwlTH5XwqCWTc29/ME+h/pr0K5lyqrsnIe9w42GpmnHmul7qk8KsmER2LXUx8RbbFxxxc3
NcyYg3z5BkuslCbqmPHZ922FKZtGXXin66rn+iOap6vrDakYXvNVKGluVCtQWVc6UrfEEAExDyfP
IIVmwGAxYFa9kbBp5itZLRiKBl5GmFhrRPfd5RBuMSzE4YohbMKy1xZ3Z2V24N+X7ARpsk4gvYNk
AwU58cmD8afFhGW85E9PgaWplY0hrqmaz85w+VDG2ZDOXTdYjt2Rs9Gf0pdoXP35IoZfLXTcXkci
FxeGqt01a8HfFHgOyrW6hZ1LWM0irkkmVOR9qsp6IhNNUaTJf4Gil7IUTQXEAPHVhsE+rYQx4hhr
woTlFCHVi1SF+3oCw4ecA5+pnHo6SMigXdua5iwxC0AZq9IwPGze0kY7qQLwkv4Gs627JQUhkCpB
88p5A0zTFD2bkUUv5TrOh1V1Z0HV4Dgt9O17nCJcauaG6bCWvjf2swFjqbeJWQCMsxGeGqFhYenk
B7KbZW0duVSn0BCDxVq4erUeYFBAf+hENSNEVDsUHEs6b/5e/jacicRjqGsd+5Z3Aj/6SIng1qkx
kIBMLPZcvrjyv0P3krB9Pakm72Q1xL2mjTetV6jKq7w8HtGMqViwtPrME1I4hIhicGlRmKOv8+sn
73nQI7plqt40FYaQrimWuCbhYatKaKNiJXQgVCd0NIoUIx80FB5/pvkcSvBk1NwaElT8uvljdDi/
LhW3bPbq9S7/c2uhYJJNzKuf61QtDJ0ZX4lxh8U1bEosHn7zNCHzGnb3y2PFx4L0yWFNpGPBxgij
d54Vy4t6GBF/XPHoUVvulcEYBaDLKyM78So36YAWFfgP9y/COX7g6/kA52Pxqj85Swaa45raK9Nv
tTFjA/HZ7ffvTUHcPIPvuHS9syhBJTlTtEyY/hvhCAcUmD9yBUBPtwg9B/7FoSnUOyIamscmklij
5gJ6LrSvCoqh1kVaSvS3NOvGq7ziPC44sr7K3fitqABjNde1wtZvs1hrfkiKZ5oagOwGHdL9QQBW
xXffHgAH7r+ffhtFBFr8qUnofhNNBaAr84VUEEl15yKVRjeHMJBSKgV1B2XSNSKxDcAds+hx5rCU
9SWqVoX8JTNkrfkFG5BcEG2WF8RBBue1sNKMvQmanbtA4zsVWog8yaIlE6pSDtFzxuBRcdeA6UYQ
/cF8cT6gk81y9kPIwxk2ZusrhyqbRCUff15guh/Z0Ea/vIHZ1GtUi8zN72ga78lmbsITfmI7DA6I
XD2cb/vuZpzUUUafSXVnt37SOlJ4jfhrnJdIMzVl7uVfleLsxGEq8EWKwL5aEU59g5AiwXxjUoZe
RO+NVC4WERlPt0F0LD8FwnXQPtgg7d7yYZQRjVeQESG03mXIEdpqq/CZ/xdB4vsSIdfs8bhHNJ6M
HfDRXoYnF5v2XUYvXoSqpqSfmo+0gO5wfInaUJaR/gc2tjDL9+dnZ9cUArtcwK7bTszBdlY4//9k
Jgtno1nRkIoFtf+gzAvVABMtVXmmVNwbLJWxdxsoOMI+Oz5I1ti1PrjVDBURYKvWqcWsmBpLkkr0
x2ZhQmQv96s0abx7tTGwHVTZ3aahu1wkJuJssoBiod5YZyLY337tMJYdh6KAMAMZj1NArUQCet2y
PFI+h2nQNgYJ7RUAFCZr2hnxokikF1zOUOurw+FC6MT52CCQProge6C4/Zn2FkyKcCTjLk2VAvv8
qa7RcjtExHXy7piD6FlJvTd1247vEd2k5HNUOIggqA/wXUK8NrzYUskHKCLTQwCuNYGuieLr4mqv
syJe/wOBmzHgiuNFrYd4XrssCZy7DLjSvAKPNoC0qoi5dXGF/U9acGdZkui+OV4gDQ34WUmYQx6c
G++wDElkHtlkrobpREXb4oL+HpeCLiRU1hr2bETn4I40nbFTQQLWQslBk9FPH9wf+il5dL9bO7t5
oME8M/bls2fIRrwYSlZH6W+ZfXv41agKQndaCXCt10HjmQbaBisBZtZSupJxM8X2gCma/U3LQNaR
a3SO7SZi8Bs7BjEsduvA81gx0ZFnkTBwU/oP7vArIClMHfPCWnAXc5fT1SnvmBwqS2lyiGp7DBD2
/jRrygi0utJyEoKs/37jcXelKoZ8L67hnZqaO7FB4UYP1EdRma6PElEMp/z3187BftNIvbKSKbck
jw8wMqUeyOI34ngY4j7L1XHRjyiz/7JTzJ8BX1zKZUThHsfVufx3de4he57BzDh8iz/LkCDMu5I7
5TrNRIPNdopiI//7aCZa8ag+HGxYVcO/lMV5iFxiWwKlhOU6KQw6AuRHszxyE6WqZ61yx4tYLeib
U/FflgjTC/0Qt//LJiV9RKJedf6Yl62r5ndCQaaf2FGW6RRWn3aBp+HtahGaQmJEoTDGORnTwZGp
l9xvc9UayhwXn81oKDTbI7fPPQCqoFRMPjxYAgfwyxtzD4WQtwViosGbYHZnCXukmzAljD0lgMUM
hmqhrAfJMxFIDP8X1ZgnfCbhznJF7WrjP2TPwGm0OyU7aWqA8dVOCh5pcKRPBCd3haqZCGL59j7i
F+Q7zVPTiS6yTKSY1aNChSvpMT/WceGcwhqS2wWNPCMkILYloB+8c3IV5fqk0Pn+qfeiVt6g+/C+
alBB3rjEEL5+5NfmbVxZaLyHWh4sONlHEk+/Dw6M+o7uo143+xfoWz97EDBbfxuT3DpNqFBkMjan
rtHI7I7X60Tt0f5BQ5ql24Ty98zqV63tTn09BF6EAKYNC4VQzFQHRPIYFJzuJCksjWnQbEnuuYF3
kVVRjrk6DKYyufpCdDp9JTDLc0WT/xbs/AXkdsIIY2Xe8lLG0mZ3l3HBURlO0MkN/lIb3HZZKXXO
Z31/daDFRQo3n51WZmXzn9/V3RQ/euhnSb714a1qPu54RlQ+TRrWZsrylxuOEK3ViYuLLriH8F5V
3UO+SCzvkF0NtVCX+Nn4T3wApemStq4RmoRIt42wZNBYyuL0RKC1G9VrHleUl+9fMCB7mqkhawR8
PWFtiKHAd7FwgJI4l2z+Q7d5xyOzKkryOggWeRrasgt7/mDTbMR/VEXHKkf+buRe6gRcyMgMF3xc
r7U43lapzGssON+aREt3RY1ymR+VaLW4r0iJf2h/66eCzVkLqX4OBH7IFKgKDvfMj00bYHNrbPFa
8k4KLtsrQ757E9EhsgWaqitT/KBW/YAiTDhec3QK3ZEn1Ch5QjbKCD9NyNoPhD6I43VrKu0py7+k
onZjspb9ijqZhxsqwTRAJ5m6sU1pQwJTCPFGc8VQnOMGbDr/7WPt7dqVihPyZ35HjXWpsBDa2/62
q1A0OK3iltZwdmrEgRP4Pp4Tdq6bz51Gj9LkX2lLeiNqgLMemoSDFdbcR+PjrAvWw0U9tQBKcn8U
c2X6BlGqtTQdus3yQEuAelO0Vr9gAvWQfQopve9zaMoxJkNbwyXADow9YVpn6LRMiqkErcu9bKC7
r5+ts5OTKzCxq6J3ekfHyh1DRPeEg3XH26FSsSEOGIbmdSUKsgvOqKDyGpmwgEFxIj0Cb+Jzk3TF
0LvWsE/1LKtX9uGKDIqUxTkJVqaSHob+lN3UuKa23Ph7mc2RKvo1vQUXjAQJOs/H5T4hwX+ocmyj
Ia2KbH/DMmGJAOHUKASdFXwpCi/brMq9hmtZqoA9YEi1w3FWti7SxR9AztavdbA/2aQHRSjORcJX
XRCBrHG8n4lYZiPJv1asrjYxeXF+1lwpyIc0me7oNGYKC6EvrbL3BU/NTJ/p+hRBFSky1o0QSVv/
DpBmaoFsMd/85UM+H4XS1ZCHE/fMwFaJOB8FmNnCv7aFi+5gEj5RTfkVBmW9y8JRygpipo5bcmuO
zmnQ+oU21ClkJwPnFcJo180sTXM2r4Pb4zrVQlmQDA9d5lm7gUT9zyS+GCgVEQuaVLQnTj2DgQ7Q
BhqNK988QVzbSHV+RDfnIrCjh53giwl+D0MIDnc5TfV8Cx2ZZA8Jphcx1HRBASCf7HsoQTEtG0om
CyXdGobZRqg9c163d2EFaJxRLTML81Zsxg/RczyemJi0dISyJn0VzXjUxJPwyNIizqDpBAYdv6JA
+71jfK+jUdosPT2qy4G4A+Z036A6YJML7Of54X1XQperlWz25J5cb+vXZuOfF4oFuwYs8CKstuwE
RizWijUNUQeQc+R8gndLsbl94N4T1fFfn7o4/ZsB99N4vpql3/4sB/PydL5oRLs0fXU/S3OkIHTs
7W8pTiRv2SPRtR3hxbI982PKmHJNcw5PubKj++nra6c0QV2vqjOkapE2DyD5ki/1Ds4/yRoZkvcm
ypSBL0ncsm62/SSRifCBNCeL2FG78+ZY8KS0d7cG7aXhpwFu+AX7irDsOsr2BUoXVdzo5WQ7ej4u
0v2nq2rAikdKvr3DhJC5V+tJdcEaPF6YRH9cMmOoZal2PVd59HZ1Prvfu+wwFfjyd0mqH+/lEOAO
YTI9EF2J67iwxk+9qc5vPa0F7E5cKLngMTkQq6XnG50gb69/WHT0AX9w9YHKHvXmffxh0U0t054K
OWHDRqZn7naK2wqG8zUG/N0zCY6fqryrpYmw5G+hIUNPen++J3KUsOxtM/JwHH9vhooVIysKhwad
FJd2UXiKPd8/GC3kkNm0gOfE4I4+CBnPt7sLL0WzEFGHhMg6eS/M7GdF4aAqZXJvpNZVBoVZ8X9A
fruiV00RrCWOs8H9SS0kD+MOEh1m77xQjnxM1wYmZFxSEr4//nAE3UKpIBTnvSeFsBkygEdNOavU
8LBl1zJ7k6cvGOd6aCdQQZ83HaCm5bWiUHz9vuiNsZlvtCYJWy9E8eeMk5nQf0GgKjfFoTGMqjbU
AV0GHTHuYNDHXcvbzq6uhGA/+Sn3nGya5/s48sC099VXqtNxjzHSUGRXwyYqG+1G9/c5m+lypddY
GBgB3bh7Mjwk2MrMjWn/2iuFuytPSrSOtc5crho7zQSEA4rlPjIsBsGj0P+Fci9VfgNGRGtJN+tH
G+T81UtQy7txOPNB807Drkf6CnmMagQklrtr5SAPxDs8/q8Ol3uoM5ZeSj9KyyuZE6GyB4qCrvbf
ygl2OEn3a087zkNlZysK85pRmi+HPLYrx5ziBL3BVPK/7iUY2uFLrBqSsIUu4CZfR4/c/GdXWN7A
/xF+9/mqLZkEMzz14/4rX2gL1jQsqF8/VaZN6iIw9A7hI2zz3vinRjlsWf8j8/hGn2Ppfv+48mqH
MuLdMX8SeEl3qqTX4VcRj27YSF6OTV1dC1Qa4Mb2NZov/uU6UZYWeiX4hNQPTOPfhqR6QCh2JMq3
1B/rGlfqyrmfX9+IHAruMDV2sKXmTD62pQMwUglCPhARrDXWool87f1PGIV0buDY9j7buehCjLpy
SE7ZTq5f+ObToaldwDfmrryTq1VbtzuihNsXV4cgWFy3JfNlqKllo0howfx774Rvp4cWFIXg9YpY
DPzLDwogj/+PDNX/eoO7B/ou1RKUyxeFjQ0Px4y9daRtwfL+Bnl0mZr+Uex18+zPcOUc77Z+7w43
kCkvbCupaZeP7COz0am2HzM8ijFgJzw9EOfxLNtHFEGfhkzNGZh/Rlp7cvmkOMRlVkEd64vR20kN
YqAekRg7BoRGAy0OWkCr8amP/qcmy3oPhGAIrLtf8yj232v06hUT6eG3ZM+mw1Uaq2uNPvDmXLpl
zR+BY4GKy0XGPp34bYMHLlc8DcFL2LiBWCQn/cMq4+nzvBFVZPHva/rlr+dMX6xi/bwKpGRq3wX3
JVLZ4RFM1bJLUeROndew9vvO1rMLxNMpCmoWfXkhGXZncDRiJVZq/POaWBPTuuU+nSZB1m2EFt3e
5PtaBMwsRBEgoz2teE8/HNu/rP8Q7/FqU5CMQsR7ELTCpKkqwb9J9AIEvi9T/VSrqZagkAuP5MH+
iDp4616TWG/Mw1NTiRCOoQl5NRS0aQVSKgnyihq71cxtL8xSgA0ChBb47YUL3sh2Qp3RMqmWLq7s
LtGo28uwIMLiRHN/O6nS8CgM97WemORLluuAQHaYNtygiAWJE6SduB2q1p5qhX9P4wGgG7sbsa0+
10dX7zeBpsPp3P1waUczw6mis7Wax3NJSw8p9BNsBLmg0BlPTgegHhG7u7sxSZmtqfUVsg7g14kD
i1wIohYOtjnMfk4FsqfJDNBUBWfGnP/kLwZymhjZAVBiX126JqAilunOD9INlaLjjeDkuKVsuaPP
nEEhokY1aaIh9LYAfcUxewmmapKvq1hjq4nJgLDLXjMoHBTLbqxqNfWlJrUKoTi7H1v/zeM1lT0P
fkKUT8C0CRIVCKs/JubGUGefr3618f9r35lvbaUTBCnNRfwNk1UysHUSxiWEkGhI6LZSyLhpt0qM
9oJfK7aPoVgjlIsHXKH/ID7x+dzCd9ZAJ2ogQ+CmnU+MUQbSbJk71kAmJxcB7ViBICQhOhY7T0PJ
LdbAdHdSl/TlO0CSNeLYJgib0FphI0iKkToPvtmcdVhGgrW7O+5udaUnygWsnC94pAic3nTdRRN6
lQ7VLl1TPLHGvPpvYYX3kLHUV1DIDGUdCRZNY9bVfu6Gt9pJU85pUHPqCWtrf7I4Rr2xNOl+Hs6G
gs20YZwA58XwjrjGaIcmxHr8N8OcpzYNOWDIHaIlNXAhHOkzB1LpTJtmkHQsxQu/Wh1wrLZeDI8C
Ts+lCSO8EAOaxsSe8gn6Nu0oXDo06QZF6QUUxLKC5VMSz9YO3trTkcapWqIiHWo2E0iuuLQIC8Z+
n5uDH/F5hELkv0OB8F4ejrtZs7K8G7LNjI0ZBmBWCzqKZy+vBC34CU6Al+keSTKe0Hpan/mxi0SU
0dtSYqv5vLhOfFQa2s5knWPcq/8Dzfm180RfcJQjcMwxbHfnEX/Z56Oq6CpZ0+R2huL1+Ezi8nep
/tKdKuUo65/1lzxVhSWA34w9/75gIGOy/md7NQ6Tn0mWsoxaX+Yg1KphyBc77sZEC52Sp2E/lZjd
pDu9BYY1rBhoJkmdIF6yP6hViIVlSSW39rAbKMnCIKoYOvlRgsV0+wVdM4CDygA1ZLIwQDD35RzF
PCJaTRYKYWqLv/GgK7PSslX50g88BpVnSDGQKHnZyHjAUNIyvTXTCb+edTtmu+18ecTOIPKsMjhn
Su+hlYcWjOaQo1cDMt9KtRBeAM/WKlJEM9jp+JFbiwd1Z+MJooTtacE7UtTenfG+wU3ScpSPBygK
PMHXQ70gzRl2IgSazndjgYUq3UGxYNjS/yUQXXQfo4d4ry3s+uf5FN7DB8HcCu5Z7e6ibO4hRz1B
RY4nIJA2gZZkHROn586pEqGjSjpgpxEpxlpYzmolL93tL8kM8hDuaQI3t44rm+afCR3ykHjdySns
NGvi2QpqG8m7J1/kCQj0ZKalOg2KtWcdB0L/TisjH59CpSFGJLM0qxnsmPcbMMTgTvNIyldcTKXK
6fO1TsEXl0KLRQLV7xDNPW37gyp4R4BcOvVTIHMkmT6apFOL9ZxxwGL9qGxDpYIxA2XFCneDqHvK
mUGn4Hc+HkFiTybdiJfOuDXIbsbhshW625RogmeR6etng1xpWSmeQe5X6680VZKQqUyKHglqjsxN
N1ewmxrnzcRBG5HKteZRd8mc7AJysC5Qw7P0dGnUNHlXMLDEa4R4O56Z1HPy3k72tG+NFiyTJorO
MpUs2XuAQuOa9s5skR/ku97Pqw/nrWp7SI9hHUrfY0X4qN1W/THkc7Zw041LpcvY7jIuRPF+izHU
ZJWeyjJ6e36Gg1heurEVc6q91xDQtMhQcFKxc543G1Dva1NhGQ4rVv86IaaTcamtmT62cHjYfXzs
yeR7pyjykvJGh9WPJXDjDr/k+83sqNA2nfwVD0OPNFf5M+IVUdK9zHeqLo8gjK9eptDujpgTBuGf
5hlUfamNkgkBh0EY7TA7gzBXKCgXkWcBvMdbQ6pWO8JV9obsjrWiED0eEQZokpgRMZv3ANUyfljz
YeAE/pVhvwqhNJsNIcc3CbzZ1Uf5QFR7P1P9xubfk8zeu4Vz15ysWcLkkZNjZzoj0JyFuN6mwjiR
4X5SrS1A0lfKm03ve/a2Ea2MsdAkOgybUz8uGbSQkKTVsau5kS33U53e/++FTijSvVlfLubIofCE
dVXU4sLn5KnD/AuX2h1eONSF1l4UyP6OPlHDPqKYa5v+p4DtrFEhkGipqRdIEYpxkX7AXRv6KSu/
+ieFtCoxD5zriRpFiGKsiA+AVdMIgMFL5S6WLWgU8/HOJYvwu3dw/BJtQRrS3L3Y4EO0LsN1NNwb
hdOPJmFu0rmL8sAtuML2UZ77xI9vtHThvHzjayCUfmu8H+Bx8W0ebTHjHn3gADobZ83njZdLg5HH
46A5KBScwROeoirgPX04GIEsNGnOrSa+uq1buIT3GQ+FuWJMAHmH0FqCstvZJFUUfqCBDeTPaItq
JObBSs2bSWx7CNxqhhf9Ps7siIwx6h+VVw9rJJPZyYKOrsEgTg1g6+Lu5N+rtSB4SzCGyxmkHH3Q
wlATuOCFQcqDF+DjCWQW5LKacpoMYo+/t9zA22KuxU+xdWhEnirMRb5nSRJagCDWg652sZEzhb5j
qVGZ1m8sY/4Yp0gdDIqsFa6J5ffI7MZbgflCgP6f5FOvkyjOmJsboS+0ob3kkM9DrfYE40Yo00IC
7l2axxqZBDDj70YdMS8tXv+67fMUNdWzOmBlJJmiY+FNEs4N2jMm6sUiKK/lbhWUkeo8ZjN+iCGC
qS/deaxLwlTINJozZ4qbcLjQVf/GfS4JrkKz2ggEoaNr7E85e+LzeSImHX2KiSN7qxKH0R7Al/0R
riEwnWuc2xcN29fBAC1Zp6Dm75xF1ko/oAtZBuOKLjuMe/xBYf3OUugdCk66YAz9XWPb+PBn25Jv
1py2tLoO7hDvurrXPM096kdPKP1BdyUmlXPa3xiYA7Op1hz1zy89QcEsyeBsJ+/Hd6j8hc+PhgUS
mgcxlKoxxpyt5Lbi9FI9UcN4UZp6UBGtk7FED9vp1sZw987hzIcTc6TtjoXXgiX2S/U+u6/2vw3u
nI67FvUvQQsKGPJk7S2i8xHiP8BMO/Un5T1FQYdki9MAbnb4INXYjQsAJGGw/dVGD0U4Y0UdG/Kh
fXRIo3U57rpKMNYZNa17f8cej3bgReeTG82ZCGSsuRXnFpBs0MhHk+x6pf4AxRZlid/ucoD3yX25
XwJv24Vs3j5W0W10jfMcPO3Yy5BHY5wUJ7vpSeUKdWA5483lFNpneIhbTzkmoiMxba1owcusIqHn
tDjRJF/3tcpyGy8J8kc3JQypA8vmKZc1zo1+ENLW4r3jYZjQKDnnCb+Y0BMfBCtFHEUK+57EqTCJ
7c+Gi1OxJnn9yr88Dpiv0umx88Ig+rVlXFckQBXJdTPPBySLwr5VxrIk2lv+iuBvYOBGCgfjQ99U
XnuiFG3n+ii1BC+8sC5h6eDCnFvYqxCGCmkdbpkcKCXKRZpzAgMrktwkISx/8Wkc82qfRKgp9tKO
l6uEQu/3GWPF4Sh1ZSOEjJviPHtGlyXQChXZ1ThaE3gp06h2YxffOdwDqhFVOcyYSVOveHXvsQ+q
uofaTLo6PgtS3CgCT2MybtpFqBIobXfRg55roHtVMBPYOWVb/PdHtwQR0064+7oh/vu8g0SHbtJN
GStHxJ/AYyyqnpKzwMbANx0+LRwocYPejNhVFyw+Yf61oFjReyPNTb9lLQ4r6BP+yGPTbZM2yuP2
LZCwanBju5V2INP9QhhohIY49XNXbEQgc8hfQmfST3x/xSFShNnkVZq6xG1TaMkZPEVU5bE2f/sf
k1cjWUu/4FO97eQcYEUOi5D0iWDEAgpG/0IAVVNxoZgNWDSksvQph4S2uBCQ+pqHuMdmq6EbcX8d
814lslU/Xaa9pxAaw1ix4RaeanKIpjXKF2wRyw77t8FAooxFTUv7J0H5ZoeCRAMoE/lkdtM0/xZa
y0+XQyQokzp9d6YTv3le6m74nAZC/Exofd7GiPYluoLkQbTpKuD4q7AWAptkG1fEW6/CjTCQPSje
L4hFq0BT5ymhQ/w0eSoh/kou3B6f2WFqtYZJMtYmUQfa0es6jJDGhyu3PtoxIC9JICUgH3h7otLt
ina9ZX8X2+a7IcAfhTLPNfAas1MAjPKMrOioa5/93lvoTE7UVHt8oIBloeGnlv7nZRZGgkGNehpt
QhjQr+63fVhnYatYghkjYA2cdR0KxBbCTUcvQgMRPKDCwCZw4eZ5lJeNH/uqLX7qVcYhvDVeuazM
AQvaYWCIxCTIzb8wFvTRhoF4ddCtH+C6TEyDL+CxYLpWwLzUPPTCLLW3m3SnWEAaXayvixo3+rlr
2UJE+W5kwbfK1aXkH3pCTLQBs8ZnxZaEsdKm6PDpaBD+WDJs8X0X8lwwyLuY5IecT0mSyRr/wGKG
ZuhVQGXY2L5MHwW3FpKoJJ62iFT2dWa0WRYfzrltGmHnoDh7reCXoI6tKqvU/ExqrR5t3GfrS1vY
ZqR622A7InVDQDYStRPrxX8H5+Ldl6NjbeDfvuAWWNhgp/WkFohHbQhAnIJdWgZTHvzC/u3qfx82
wx2bNjdRwxdMZRUVafIg7zY0Okzfn4fH7sNWmMkSlnfNU36LMqD68t3sh68ssZmGMp++u76QKodA
jYYTOLUHGByk/K9OLlyAvQ+s9Kpc2y4Qhlq9IYFec3wkUduxpv7tY7hO+HznSPV+oC9BSkTd7Ndf
WOXIWf7s4MYd+wDBXXZU+NR6qw+yYZVRIsypw2/9ZM8jT23pWir6ogeWL5wGP2lWwu2JXMh3GlrI
2/9L7zwYPMjD1T1L3Q13p7sy+hM2CByj+TvVEyAoPUe/q4R2Q43e4tntTi/w+cSDlljdfNIdiz96
F3A1upgEHIxQGBNvPH8USN5fasXlJChLGzM66ZQL4CAluNkV9yTRGwqwabn548YH96J4w8BJBhpn
OSW+PMFuqakDRRZAuVAksDNHZe7xRC7vLSDG+Nir3zU7sBLuE+UAJxyadgbObEQO/s/zbqrVfjPY
flGPpaXWlL0jrhMLDB4KryOY7YrcGSw8ugUpJ1XJJWrClprl7H2h+YFSnAo7XXaYDb1n6IxfFNIj
Xi5exv2FnHGRe+8xONrbLO+5urkfXrCM7MDe/kNjzs/EdHooeJFRAwaa+jJa2eVJ1INyBZvrYrg1
GNOuBJestIAhBO4FcSxYpq3akzM+SNsp5oSGLmR4hq0yoNjIXtdOMJ/yBd+iYaIH/t6gKY7Y7Jbz
gwKPBpIMf2LsdeVCr8yz9bde1dmvmKXgSsBJ+i2TR6fNneeZuW+NjteRgs52DIfK2ylW/oIMvhtg
Nan/jveGTAQofdA3gxAV/wrCSuFE826gC/7kz/hGCtzmSzB6YHwlgxvcfgupKu1ujH3mFyXSbV+T
ZaNRYrskBzW61Yjr5z9mlD1hE/kXyIYqw7gDAnuKklIR9abVT3anvNQoIfAhXlrrPizG24D0Ksbh
xTURbSE38ka0ifIlSuEk3M5IAxHyXssGDq+I0C7VAEH8pYyMVjX0RO2Tc730Z37mTNeE4rgDSUKd
peDeuRjhdXtED0jU5u9nm6p2qGXW2slVV7vKdpRDGXspnYHDc2COwmOmYH25o1g0Kfol8Ad74b4Z
dujDTqcpfJfuQw+LY3dD0XruevuKjM2xp90lK4YVkCbGRfSwhfgysUVsyB9LBVZh4sYx3OzpXEPA
6fHxVtLILgxpb/EpJ+zAMCEi4ZDN5v8sUGAYVCluN+gdJy3JgPb9x7JzAfTAC8/ChwSueiPBFSl3
tY8FCIeiaFFp3w8TGkyB3LF6zZIbWelLvFi6AP0dtSciYOP/ynQulzm6oCU1ZGL2oWu+9Eys/YOm
mr1ZWeaRATVc8UELer18st/gJ9go1awzX237olQzB/Zp0LEQuEBtvvtOQcx5nqaHV51pjr4vYLuL
8VR0nmga94xNypJFSiGZ8/YwvMjCpaLKm13eOZvDnYubhSszTXfVAHUyWezitzQtYEATGnOSWngZ
da+g7O6kna3LU+K029hmRXBXWbNnSxJgO1k1ph31/bc8UMg8MqNRUwYvA9xFDDqdxdorav49+KLF
MHpaYfGoFhrqmIM7fGWY9Y/xD/juLzXkY2/utUEaYUufsD+QuKJQiml9CjXusYAaTxn2+aS30cAs
G4CkQDLNSSRxw1uNa66QYp9unapnSeu7mGL6NsIiWzkjjG8uyjZ0K9WUfK/PhHW+TpzRc99+4vD1
rOjbpzFdq9xqh70lJhMSn5MyrTLDLq5RqQcz5VflCozccFTO1I8pfGpBCoCvc/cm/E/aDMDUcli2
MR5Sh8KneeI/iAzFCenLOID/hUOJljlqOheG8Eg05gkb5P8eN22LMltZHPRpHbUKjhfP1tWT7m2P
L/sF1DRbRNNM12PEnonnDoJ29Rsn+O/byrJqyMxS45fyATPzJcG53bk0x0Z6WFItFWz5fJUSJPhG
pL4mLh0qdZ09quKYHWP2hLz60WptLbwRzCVnuQmbiBVQwimKENl15L+L9F33tEiG2qqIyHGaKqzF
vwAc4T2xsJzRcFzt14tpo/3Iz4gJi2+i/8XwGHACqfmlU8TBdzG/5NYaMJ1quPYMAfSxjTk/oHvh
P3GEwBCeYipUYY+mIQXINbVi0ssWc2RAqC+gi7GyoaKmImpptkgYZl0Z1ZcteVyUvWyxLKpLofWY
9dO2YNfliK5pm6rIzZ88rwU68Qe0EdImDJ+coU79NqyEkrnM0SgSfKXBZyLTrpIT9iAKjYeKa8Zs
4wqPEbsrPw8NT0kOXVqz6upEamsS9R5n1oSGdc1jmOk5sTBSYFQlxYPIXwdO72IvkfJNgEHnzmGj
smpDyd2MvLHxen4ea7c2nvpiat1bHR53nvjCA7ldu+f7/gM5fzutpoOjDHaWpWstvLVXo15x9suA
yMfpIKWdwmw6Z5rXbdsbBoQ4HwDEtgPP8IJ29A6Nd6ciYuUqZEjq2K/myW1LKCICYWZXVRQsp9Vz
Fv6IoOfVW69hdcLCmuGwA07CVYizaUQbFESrDeIIuKiDSqPkvYydJ7kkntVwDKdB7ka6A5GCOqI0
7RGzCDS/8S6eFu+9yquWUIswj524Nh31co0AdDZKVMIEKOduFoEIS0kTZiMfMaemvi3YIVm6Lljq
G+nEsYkl0vzjyD/UCUYNRZcR5sq76VNgflOjWFlSqwf6fxj7CGQx+ozgGpqzxhuBwV8wgjDnhKiV
q8nxl4+H5jYMEMevostUuQxT8Hf9lRdnIvq7O9nHFyg01Cpd+EVNDyGNutSvSyrRaREoW8eZHvDi
25KhM2BThx/Dv6vQKKk8Ayj1OoRNVgFaFqOkpXm618RcH3ONo8e1Nnh/PNDg0xCbzfASAD5lBYX1
grjpuHFjw7H7MTSqbE+u/eVq70lC3tYEGScZG6LOWBLbva13/6gTDHXMJLlEz48fuf742DbcHMpD
fiJo1B6fJWrTwF9/T9BG8hSlqLsqlW54T442rrDexZdluJxLIQyCPLJ9otC8EgAbhRwOSEln8BIR
IiFCXyhh7OsXg+oukg1yq+NPE4+/5vuEr5If7hkk593jdMJ6HnkLLdIp7AttfmIxcYq3KkAS1qAP
WNE+v+BqXtlOZThQi9mJ7OwbN7ZUFbaKA67RKnmCQn4oCrTc978rSl6OtmrR6uR2DKoQ/ziQTVcV
vLwDAd4GsEYGeZHmk3ipvB+pTpmbEPQSOcMnF65moo35+WE5JSXEs/lVhk9/Gqmdz0JQe0DNESYj
aooFMaIyOGDiCjRtFxd4spLgjfkR2NiM57rQJPwEio1aSBEjdMv129B1sKeKDn7SlDk90foJUBND
d9NVpgWjvUaGMi5BQ9ShnTC1ivJIBfkOEyqXnn9eIQtouDlgC3NnJ/uvRcEbumVeS9FEDGclUs8b
RMDc6G3GA9+m+Z9po7VGSN/GaM4YaJnY75mK2GMmMJUpHPZr7hHYP1UwDa+YUPm8W/gcH1lL8jNq
exDkdH1K02I4q9MfHF9JIl2osr4OueVFhWzRxq3xdRLnIyxgCnM708WDT0LaZmOsW0BmPGfCLn1H
Pt6uv9ZLXZeZTwi4058NvyOBCmJOFr5wwHnp/O33DtaOtgtk80CWp6+vAWQ1xhVJbNYrN9eb8wue
ojnJK8/pSdMRYSkcww7sVX5IzuTYVJ+a2L9CD36+fn9Jbd2F/sTlSkS1rlqYx12uzZiQQEDkVU74
uL2gmK8tSIz2w0rkaW9euxBoMeOjxmyPF4zl6O8eG5p05ilLD3dTM3ubb3d7xE6qKg8blDk2VwXu
bGwzAtXndKWW+uUGR2M/XokguuEKVvIzmUJ7xnYXeMqCVe0wfS7+Yw1/rgK7zBBCTgtBMQOPhUO4
+h6slLeIKxcscTjhfbwB4n2NlBEF1NkV6di+QlAL/asRGyypkF0ZFG71caufnoxckDjgb3fbVZL5
hcR8QeWh8yRf0sN6fvcedhnfUmxpl31d9L4+bo4DB3ta+PMxgPgAd+H6tjEOHTasO3qwU+3L7mud
TL06pojoI1k5zldpTnpAA4aCEcAoMz5RNq7SAETgYOd03TkqXPx9GJ3khQ0RZdnBawfl9bQhfSQu
TJxFKHsMZqcL+jp2GTxJvi3BMlgNOsFlQ6HUyMCSmewG0aHOWk+6nDUhzqt5aVrGblTAqumNHzjb
0RpaNgZRnxqsyPBGZNu3UNhWkvY5UV77KTtzu8HqrXg7/3MWKoTip81JACENGlhJSEyiVU0pcVl4
gZgG1PyWs09BlmwRak7QZpoBE08y1cJsZ022iZvoKenUChL8AHgHd3G0N3oQ5gC8BiisR90fd9qi
kJoIMDE7VBICy4PZkxHS4RVHuGiQeyuGFyD1z8E3KVUKCoKwHDTIL97DKht+yoZLTVeQgF16pLSM
UOzv0AfJTFNAuzR6dok+aIS1ey1wa4xitBiSeMcrZuePeYxXedwy3g8SCc4Jn+CZa0IsJXIe3spx
pDylLbnHzCFeauHUcOpX9vSL+wytFbQx/4menNSUDHcBn6GO1b/UgaJYj0YvUdpXtWpkyABw4jCX
Hp24ARcXzAIeSl+ExV29SGvUtbEfE1FR0LWUheMey7P0/1XhdcWAO5uFAYC/qldFBw93mOJs6KCN
wz3n7yPzPKwo0QtPYFlUj6oB6yGc6hvt+I9X+mQsWVcB84hsS5+7tTzdzmhH94rtnpQpxTNxcSy5
HCMDKcTdFgo+VkKSxp+iyhYTn3LDSQW3OUGRmYbqAjvozG3zfMxY878Sem0qdpzlVeRw/jZgNara
qxPfBDmRdJbSliuBD+4AXUn9RaMA6+cQSM2LXl18NML9YuQ70AzuVd+SBVqjxX3z5j9wBBl0KMYn
eaH1Ty0EZGtifK/dFDxZGXhHSGqtCLQyZQhIbzaijpWNIkDuCk9y1r1uObAr68RLg2awf/j8/OEw
pqmkOChzAdi3QrZUQl9pjs+SIBF8zBGEX5k8XOzvqcl1NVqZoBv/e6DXjv2/FE2fWG21Cc1V112M
7CQaV7lFY5C4+Ao26NxkkZcybB3dv7YnAQuOuz3gcnWCbf3If7bORJl1Ee/gyImW9jrhKVqdp3bA
G2dr+cHSX/rVmqLbN5t9uNy8xWDNGlXctKbdggCqhtfY/AV/w1xchcxh9aXZzEnbWCsBbZdkrcWT
LbXlOGAdcmZc9ZbbBV+I9g4DS2yxHSqB7M/SxB+fKK1GHhRBcUNecH02VWn5v6VJ7VnxNzC3DtcV
JAlEYlBfhMFzg8E2Gt5Xq2UIZkwz8ha/ghbi+XCglYCIBNmByepHG3TyZ5vOKWKot41BEgvgD2qV
M38MJcmelWL7NZMex+aQ9QuBSC9g8fUCfErou9n1xJMIZX7kyw7l7DF3iwHHiQO2PiFP6XroY3zX
H7TOlYo+3BdVzGeDaq+rMmoVMKhmjj1FYgewDH4ps2k+pHYb9DBw7vr77zJFiS2+RELUzHHD+hfp
deip4DMDstrA+A8FIBbbl/FU9rnTt/wy1GZyabpBAJqhoBHnPSxcrOvmqiZQehT2ZIbgIE92huE1
9FDe0omqzSW3jBS4pPvIe3zmFnt0xmKydOPJ+OS4rN4vF8sgzZaKqcOHJa3l3DfoYQWBsOoIgyXJ
YxWG0Y7sY5PzUP4twMazWy7G3DpAweel7uKhfDgR5+OI7AjU5dgWSGUOIx8T92gJ224GnU6L7Ndd
rbLCtVC6kBBF4n/jFGQPPZ1eTVQ3z1HIcm0AKSkMDn+3c9g8ZVClGvBo+KXKxtcaotZRklyH+W5g
CQTMhvve4ckqHr8bzJ2AUx8iJulV84hukrFL1lKu60iwhQqG/tcdXcCke5l8N80ADJndSxg0H52o
jbH3ap+YnD04KifHH865cGypuIeF7UN6AaqySyT8fN+4eBE4FWO3GTesx2UWfASs+TSgtFcO3h/z
j0DFnocMzBGaCXU7oreGiEV7n6L5TC5cwSSTqK9lxt+kSOwLl+qp4yNOMcdNSACnKRnX/cC0wyPo
nAHV0t+Wq6qgohBBRv9NiARVDy1WjBA9moLuwr1HrW8hGh+BpAPxTAB8PqRPk/BN+MxYmUrFXveH
9fxDOtwWYg/7jsjvP+2LLDrLeuEJQZ8PdM69B0iEC7kdzL5HLyM3uuEZ1agDeKiyrrlUoid0ZArO
LlJnz/ZaqY7jX31rWh0DsPIA3LIZKfny7RI5FD8roN9dkS8dnlJrGdtraCMalhkDrgjPCNIxCRqp
X3KR11bDuEbyYcQTV/FzPuqOK/569DwWseeq/1R3jBTW2yYPxdjlbrS+RdCJHm00fHcEiod4Mspy
OZJjBXI9oFfZ+2HVsYMv/8Df7AA2+VyYAKNT7rUKA6AeH7PMZX2oihlJJKaUF1hMErB4P6JMueQI
tSEU2cIPofzqkOINykr47kEpKce2/Vntrh09/cRHxI9qIUffPl4PLyJnWgwNt3CibNLoxJEk8gX6
WvkGsMXvLCrwZ8yhjEuxC2cvj3mEHSQFaMU7LFQCE0VpQuB6veegqZf03AXxE6ag68yxq4UycT8n
TWJZn5MqAA9ZjhqBb89/PR93VbGWgL78h4ukpt3GmttWMYsfJK1QXxkQrR/BGXTzS5/e1IMsRuiT
dPt+FxaiZ9cAFMea79s3GL5WlCy7X1d91AVMFI5OkyXpmHhOn3WP/ZaI+RHwN3Yp+DvFw1OqiRI4
+3uj17B1PGXe9BhuzdgjYC3+pzcyw7jeWmPY1gylf7/tlzuIfoJIZMBlnTWhPltUq3CpWw4/W8bl
cBvuDHgRJ6NAQ0vIueKjyEOqHF+6CZBeRRS6l4if0ifS/LNqG5orvnjp75+8RvmqMzbnSXenMCTz
fHvbq4qK63YA4dxRxW70QapXpR5vOyf0tktug4Jr0OmwZrbw9AjUKGsHNstNjoDJq6m0w3LK4379
JVBTYMC8OqrDnjJh+1pVC1B2/1C+X4Es3ZGalqFIMIWeDQFNiOSDq5jBBp9LlPoD6ZI3AJHG66h+
eNs0OeY1WxrlAivTcgxTRPPoZ8KCp+XvnfyHXZEpA2WF/90nreUbRvqydZeI0Hhx8QUl7mGavVMt
ja1uJRKjhh1qhthLb1IjW6mCNz6dRl9vjKjHTDIp8Gcm/v6FneW8TEndXm+WDOgJLGK8/Zw+GicM
YO6R/hcezMXqXHlvkhnA1bz2f0u5oDNxrkLP91vKk1mzPWr9R6cbhcS6SGC+5uYw4jzY3NbqoNwe
hXu/H9Qf7nIlmOs6hzkyUZBuS0eGSmssrt/FR2XyQKaRxgrxLAIrRQ3Qu5yTmiFWwD+DPh0j/w/2
vp6nW9d2K0iPB5CebY/nStGDN9PAQ20hMhe/6H3DPdQmo1rZgqUJeVZdgpjphgWQfVv/Ko98YazV
HTbKh9IQgxNeezGod/XKK7exPoSAbrVCjV71dBG9sy4mAah179RzbTaNFAdKEgyDEdrNqUERk9C9
NRa0hUqdwvJGjyDCIi3VS01DPruY4K9pesjSk66sTvMDa8gk/xmLh1rKzl6LKmcihfT2U6LaqUZw
hFxW9bTxGm3WAc5Hr19NB5ltPtoVI7438JJC4008n6fH3eWaUAP9HYgkIobSXRr9HGuhM9F6bCBr
g0n4DKJfksvXN5HA5bJh2L6ZKoaJcXZG+1yFGkAsuWXXctshfMoOsecYW2wgDKDrAc5yC77evV82
2K/UhrTuLaEVEqNtmwgGzLO2ZYYJBo1n7HGZ7vthm6wuQpKYtKa9oGYUnFb4wdueACbYLOa16THI
X7DKeVVxQyot/+puhenF1E0JEipk5BlWchshAxxz1Mkar3OlzzN3wvBBdD2pch58/Pq1f9WBauWH
oIm2uRr9JPxWKcmUkV+bBPkMgLKkdmq9w7YubXsT+4b/5yYhhs2uSekN8GFRH9Noz+hEY2S1/wua
BS94oaTxbbgp2qQAYWQKmUBw9JsfpndW6MNkEYc33X3U8KuJsILzit9ZMJU3mcHTjj3nuGNqcCU8
NN//AsF21PxZyD7OFYFbLucVqf3ra6IGNj0nLyF+KPdiXO2f7ACm5Qcg51RjnZeIRjj2Ge+xOSED
cPzq1NH19wkSN6ktr1i2VFEbUnm/XrG1xd7EMSkn5R8YDlhWvdnLi5R/zFsTnWrszKngX7ZvzYWe
hhEQSb2yqetiXMJDiXna0csL46PW7GIZ1lxaJeKynXf7J9eXfJs8enETGOlq2cXrOId6eVD+RPUp
WnqWOlZ8iXRN6JIfPLC1Uze5K2LGMAFgGdbXGosS8PzNDxqNHHHBf4yVEIdNYs8XE63jwmR0i0vx
DFB4fpExwnfTb3nLWHHU1L3YTaqpE/lrQYEKkdiTlvTL5TRbnNcijFr5RLL7fmsm5Wl8bTg8MKw/
fqC0h7LsHNW822zWbrymFJMxOgOsZjcSsvQQjwEZg5lHeQH1wtRIDW+fW1vs/XERiNjvDdD8wP7Z
n1EN/Xy2FN4iRznQt9H5Z/S42Z89mtsgaL1R1JXzm5jTnwYD+RxjWc4c18yCy+m20KYXXpow4NsH
RUNItNb4oyISzkesPl3lKNxhPckGdS69iPicU6u01sXK3I/Rn28zYjm3b50nW+cEF4LgWVzvPluX
75kywnd1AGGuYzz63CBn+VPQyw0DP8Ul+3TZJD/s3kNMYZZsPx8ZFxHL4dA7/aZJm9yuDqS5iegZ
7cXhh9wbdQyqukJWpEUsDFJeRSYdlOOE71BvsZQyVU6BYNj+Wnc6bqAra6ZmXxFivgKYMXt/4V4w
K7weRj34rwkLJrN0fDQhdtPJmVAQx8olO8r/5/PNWW/bvN4XkucXFMrxcj9aQKKBfGMmuXXmUYL8
pvfpQ570KsawO/eHbMaFfrtnrCBS4hrRSS2Iu4DWjM9D4sKui/qFpbG+k/IAWXw1w8eH36/ktoy/
njMhLFwKgvsgYUfyRazH3hiRsstBv0XCRG8ALAGxaSHRkCjvSAv2r38/EyMcaSafEZU2HjX69IPg
EQf3wOdJYncUJ0D4IAJNkrJ0ZVBTUDueloq8Zslb72Jgi/PpTVqP7jNxEiwY27ztSOFPzTQLVCfv
kvUaR97XnDplQGDm8kn76pkdyCDpZNMPHTTcV3gPieJ6zU0zJdWDAARElIZSkau/QNm1eTmsDn+e
/KsLWP+r7MZBLX28HahQyr0NW4rUvjt+B8eWuDg8uOuAAogGEFv7ADnaytQMmORLgfMfsH4yn9PE
SWdt0m9exsemyPxIwNbdsglTFZhzZ4dFVmitknD7TcPaw0PtPYnRoVsf3kYJufrqQ8bdsb1RLdNf
GKepCbISg4ADt4YtUoqjSFBddjGwUDC9kYd1tcFkUHy13ghABT4vcXDBA/B0WBN+wr2G9fAn0eTE
CsaX8UPeJgKPGh7GH68jCMzZw9YZgDHOA+deaKpRdmwePIT4Mvjs7M6Bqv6v416fvgLj0hzDxs4v
TPheaklBL/zUhfzuxGjWxPXG9EZBwLJcNd0TDllRb9x5JbKAEebj/4CDhZWf5VT9IhgL7c+i5/YQ
mdwm/CHIZnkkw6gleeKC/2dYtvAubY3m8F5nLPtMTU3/XARNv80FBWdHCEcoj6HHBS8Co3HHc2Ux
FXlIFO/zG9JpzEw7z9iQYwTEd2KKNKZp/L/TSchBUkMJZEb63qOY0TYXRXvQ7+AgCccfOYRv1iar
A13h63erYAEUt4vCtfnJXMuTRsA95mboZSebYtpzkMp2IyZHia50RpKts7spefBZgz97+uXDtGaA
Tig+pj5pqoHogp7ROPPke2M7NyEJrgVxEEFmAnZxkSAO2YpESHKYWdcOFBbfuyGcdnfWk/AtG2dW
zHAjaojdATyyUc24nluirRD3BOkWG4rVOhb9sUi2DnqR8wXVDx4QfMgUv71Xu3unv2ADXoXnjTvW
AX9DsEDTDn8iDVS0tzS0X4OIgE60XVlBMstaDj95XNmSJp5CPjdSJrriRAASliaWbvEkASLMn4cE
wDTI/FG0eh4gRnpxudMxdNUP3Q0uxC6zju34hyubGLXGra9RvNBC8g8hds++zxWzYAnugDusXxkm
s7mnVelLYtmggDM04O+nMh/If/UCNQWO0AmU0Idqdf+aQr7vqdod53W7i3UmoZZN1lAghvsrsxuy
F7+RQcYTbAqqmnEYZHmbcwe++xqYJNsguiWcKw5kCg0X/2Xz72U+++hUVWCTsVtF3Lr0wI3qHvpa
/3CFsBQH6CsbO+Z/5sVF0SA4sqKwkCim4o0uq6LlKRsLLWpo/mPtKVJZNf7QiqagcPJHo6+qwjoY
xS6ZNXQ+t3Kkp2rdGWhC2c4IBo9Iy1RGnW0+WxNoxPcVxzcs4cUDOVQQ+dirkTIZakbocnipbfwg
65Hcx/KmdLss2NfWVuDDsBOjOOrAmsVtUzgSB0dspc2+F5439KEOT3sVM6CvbtANwCLqWV4Cx9xd
DkQd4OaVYnW564hYAOdGioeLri5BCDL6cIEaMuzNWJdFgH+bYM/LaqZdf5BARJoymNhoqQyqRW5j
VUs2I4oJPObbniAs55dVJuVkDTogrVjtAwpMCr7ZXWfvfd9dDDB2o5JP+4p6SnX9xwiB/vfcaCym
AyZ4UbEGr7tsZWMEwUC9qJssNFOL6KqGVbqOzYYWpU72vlIp9gwhwp4dR5SpsUR3pz33LR3Ea7PL
+EJ6xV7wz3PcxE6Ow9NaotHxQUm39fU0jB2JTwYH1wyoizBU18LnsvYu+ZrHrR4qjeCGaFKEKiKW
2WZDoATueBjhIMaSo9AVG9t4FKUnLAYZosdBNbzCr+KcvGUUGYv40OMpUrarBmuRH45wuy5ZUzyg
dMikytmOZkf6zcukDGTCPKkpeavGzs61gNQvqKtgErcl5iZal6JTazyLsrAEdI+LpbehOF8b7gQl
eQI6eGxlK2PsBh0LEAM1qo5aG1/LGJell/XzgT4pJizTqHSyv9QCIYQRJVUgSTbar8Haz9epvgHk
0kFhF+yWOWG50bEigPu4P6aRj0yYF+mMywcGVJuBfDx1uaJ7E2bFnKwI5j6cIvV1/Tb8JShDI4+Y
JpDlWFh+bPEGf38rG29P+CzhtBKbDhR+MkIPNKtBdg59f9NGUmjM8Lx7GmRursIaM3pms7jgnK9Y
0g/ttamBVTSxt05d/WZxI/4JJ5TSjaZqo2zwsnLyC6w+4dwD9ZIQm7Fd4XLPoz+PL3c1XcdpWgnB
/JdioVTLRV8ehDy49f/ljmPEEzuowRJDbJulD2LUO3pvMgPMrbIsb8ZdfDr8SbskBXqMBlB/SZXO
MvqvvV9xtbJw7Hp2b/8uEJOayF9FUoCyKd3MgBJVr6nvX4VbMo4JfPWDR/BddWzBCkpn374m4oEN
7aNK7jKKPC/NDspu1Ku4/a9EpZpAorJo+kAbA2YojtbLs1IYay0rpgka7ZraBxV7pxve1vX5DiKy
brJ1eEeX7hAwkTa4SP6MLwti+wfcYFx0HNhtqCNNuv5UVwZ1Ro0q7NkiQnuicP85Cr3USM9hncsB
CnfgBwsHSkwk5ymo7ViU+X/hJ1Tm4sB1f2q8UP3LmbRkSDMxqrP/FQg1ZWmqpeSyCUzj6UDe7OVW
xswPb4AnHuCw3pIcr0X3Gjekab2X2IhBSu7/9ZagqsN066gsCb66ZwKr7WKsQBna7jHUadPu1r7C
nx2859fdDyK3+pywx9vBXU31UKNhwTEPgQDFZDmnrSVo5+qb4nlyMEkDmLCxHx2ys0gBgbHUMOv0
W1bvSVAjCChpTjIGItjbGTYTOsypl5ltxfymXmrOhGf4O334ebicKAM+vU7vjySo8QaweA/v5oC7
F6Wn19l4uFF7kDhoccg3NvlQcVDGlV2hkvClpgAk9q//Yib79pNr0+jlsx0xVQqCBOgGaoVCJ6pM
JsggpCASvYJW+mN5xhBlSnFMPof1spt4CzeLaNVbUs4pwUrUjCkNY7aGbC/0v4ULVN7XPolWQ7W2
uHO+O/i1JdbDl/yfEwMaf9xzSg7T21nwg4YO5Lv6YnrGtnCggK0vbRIb0jvL0hRuqxaT3s33MKY0
r1xTi4m5rrG0+ygKzyV/F379ZNDfHreEwuHdgUkTQL2vngENvhM+1eAjSk8AH/PeEq3a/JFHZUS/
tPR7g9/O8LnX++mTl2H1iQCu8clbrnvq9DJpxoo3mc9PFS6n8sh3QL8PJbujgyaeUVcZ1n7Uien/
dTGXD9wnJVxXk+e/RDzs2LZEFREx/cLhVUfM6lD2y/iq4SVH53nxaUr9kWyjIR34e1a7p8bMlAJN
oN/5qSma17KjDuC/IiUPd+yQbNi8K1Edhh8wAHvloi9cYobjrpHLOhhG7fS1L4P/9b6M66LOUNwc
uKt5wKXbhtsp3yDaNvxGWXH4IZgVqRypEF+ewDQTLzSkexoRMeTE0QMjH3QSdPAGUgKu/AcSiFOi
5IvjECO8eBOi0j7ZEZcKK5Obfq5k9J0xInyoqhEXEe66YP2DBJRWWQccJrQNdzkjGssnXIuEAt0p
Wv2ovWXP5yKBexa031NLOcscp8Ui70/Eimq1s5EX28QuPF6v49WjkYcF7n/dPK6SWUW/gD7PiOWt
bG1mYVB0jYKw9IKsoAjgbaWO80YX1vd7HLlnGvL50odRggUmf3FRJTjAD+vye079Z3+7xdSK5MkO
Bd5+dwBS5hIuERDkD8wwIorfYLJ61Csdn+2D1ygzprhqOsM7dAhnwfexOxuOZ7oNF6ctBTwohcNu
iKRxoBq68Wy6HYkz5l5pdtCfUzjQ5HKwHutOxnqzTtpu64OOmjmVxjysdjt6ETCINy+VejTNFy0l
nY4N6YaJI2vbiPIMNIF1y0zOLvQpx1KOreVgbe0v2tPCM+MNxieJQ39bQTsUurer5OqFOvMt7O18
r6MszvPD6myd8SzI2t7TqBpNmfeC++ThhnEhSsFD6Nkozct96t+SXZXJUdtiZXxbpFp6q9IDGZgz
5EIK6cMh49I2i54UrcBY79YhhsF0KhXFeFzKjaQf6/mMSC+3w8mvKVoodY6Y9xJE4HVu4TZSIUQy
U97rAkyw7lpg3Ynd9BxsU6D2hIoSNtL6r3LHwUw+3WEd9tyjwraqUexr5zkANSuP4jzbTtBBb3/P
p+qXytshbVg1XY1riW3wxAIxvoR7Khk8KQ6fuoKny6ceZkSFn8gSNkOtwV0IJ0F4fw4q+tDWXCZ8
Mm47Ko3e9eGEatqgdJCsmGNn3+tNCfjZ3CkQF8A0JEapMCf8rSYGLbE/0jOXLCMBYwIYyRO/3ajI
CmSUE+EmHNoTs8+IsAdrnxpvEF6K7nqJUpTHZubVLb2+rk6HJe7JVevJNbyMs5sRMZJpvVmqsIt8
QtFw9OyR80x7QZvU3dnjleeo6RpW/RqsNjZC5SZEOeufTUjc6FVqE3z1YA030EOisNZgMl3wJ9iZ
0l27mxCioIncb9dH0iEYufXAKedJMuzZHSPQNr7K6vi3nkJ4iwKcyt6VYPlR5SzmDVc7H4lkJsvF
ra8/o91raKGitlPsNqseFyH6YTDFpF7YcJ9WfkqEuSjf5bFiZirhGFLluZ4dloqhC7i6mZWC+LNW
D7pbDTdBelKEdvMlut3GoDMTwZ7dbBfLctJ3nLk7pslEBcfxcLc3e7iQxfwvNMDr7x44MiYI33JO
8HEEBrLcqzOD7Cbd4U5JewhBP5p23MWaSABgNXHMs2D7KEadpiEQPF/mz27Zot+bwIm20GZe4O1x
7mPCPv+s/Rg8cEuaR7Nu/t3cq3Xn5ve6ZWwwa/tagzW5BpVFbihHrExfVtTPOTZOtBdF40aspkPG
ONHcf6lB25zgqHc/tuaq+43timaAGgJ8NYeKZxn+tajY6QSiyfRAQnrwGrWaCmAKfhRP/IW1wTC7
XWrtnlzj+kIxOUhBvj7co8x+BVRKYzN7yJCUR9LkKJ/1HX1kFGm9BOoO/wHbb0aLBr+1RzQUBzwZ
zaQBsfLG4b/t5a9gnXqZ3bBrI+1Zs12oL/pqjYligaNtcGoxUM7CJw4gYMtnzxAWxs36S+wYp8Cs
zAFaNx1XCWCAOofOibAQNqxbhFENM26k6iWXwngbqjDOMRRx9mjElBtNz8NtDYw8RkjXfApQtMDU
DSsLXVM2VlKaSyPpLXDYLjf4t08WFszaoTCNryI3G2zRFihDI0naT3F8SB2PBJUgAjFcc7fipJVE
kp6e97JELXdOIzmZmrEhfbVOZLuHci+Y1Y6ImJhxKTwIB74ymcvz55LReAmd13cWAWcRm5vqNazQ
u72cO5XDmztyermnYUjkPGRhMJ0hcXGtBkFNqhqjeEWCGPcnj6tqFrehftM+BuEfPzZk4oYXrDRr
Wm5WGsuMAHgewsJwMuovcXC/boeX9xAhUpx12kYwMr7PCO8bLxrkjKpQDtq6MsuUZelE6FoTALcm
N4I+dhF1/g32x4gqR2xe7ASOjCLAYYAGvMzFozswK7NCubi99GtMwk17aw5+AAvFiC/qcoD7EVOO
vEnYuk4vYyi9UhwlDbLMh3yC+YHD6q/9qGP8Gx3QcHsbLo3psbYXhXduiw1s4mKZ6RlunxvYSeqh
R9rVRtp3zDeK13u6KejY0iGP5kIweULJJp2p7QS51s0Tw5pzGLbqaulyZP2sAAxJbojefDumowNK
BXdvW58XyevqwfvF2S9cC5WjS6yhxq+VFnKITQWLpAr3GWE7U0KPsqEMVWyytOCHfs+nMfLSt5+U
53uXIIa39VWQelMarnQPIhGFbGyO7XtrBTwuT97EKh3eXdsdffS+oQyBIAUTBORpGGGhYNB3Zhqr
JfgOyXWq3EAo9G/iO6+WTO5BP7wy0z1GvOHYWBJjpcwJ3jVS4tUM90ngkiMYKme+GGJ8T3BdXP/b
yoHX3SXoH7tmbmW1Ovo/MEj6lSe0I22hBfTWX6IUF9tMaSlxvlbQgZ5DkX/ALWTk50lZeYd3paj0
MYMVFuSGz7rVGmKoZpiYZ5E0CMwaNTBCCiHF5YIcCClMc1uI6hvWQjEKAo1iapEjWuh7BAbAgN/K
GnCg3XEb7V5OOn6+Tz3DgFHT8EpS+jeW/4XvfX/pNuhn8Pc//gb3kR8qUngC/UuyTMhd55xQhugq
WuW48Y+4bZmqLynzlBeMmm0fn11BPRzd8xQf0SfNH8293pVA227U3gzB3FZoeFpIPRVcmUFVHbRR
5KhBnLE5vR68Jd7+2nsQT5u/bkW/qbXZqtD+yoyy6tYuX4N+0k15TssqEDCecVEDv4GoqGY9bpTX
XL6c7+e/RdCY1r90cRPAb5zsZ/pmMp+R7OxsrC155U0hHr9wE+jqnGII9715bgVJ4RA8Z9TsuaZ1
lzWmxuesk/WXd9SYFNu8JXHUrFaTpLjhxgqtU+YxEo3b5zl4cOwby3xpwCV0r03CcJHtiI1JRKEg
/QwIngd1csuuQNdPeiVSUeydE6K+ODRfZfjCJHWIK3vQ7YgNNdJkblNdV+cMDQ8MHc5LX4YGs60W
6XgJi3k0aQAxLU1axb/cl+/RZFHIPwPPz/RbDsT4u527HJjKzRA9ImEFHx4D0rV/mHUgsSMI0SeV
zG+TXhCyMPVmcXhAQvh6BT3nKReHkfJ/9X2+spdVXSOsG27fRS70vZNzMiNl0C6hMUu9Hcq4DBBI
9YzWaiBmHAxWtTQRucPYsbbkMXnDmtUblp7qkaCHgV+tM9vXvTz3EFFJddOlBpk0L/4gL8AeezF4
ZLMSV9XUVsC0iSZBB878nnEG5Uao7IUkyeXLNzAI5Og6ufvImYNeXJOmmQz3aHwaRDmrRTonxOeN
fdToD0ZPoPVbAJk4hQxoNLoyrXN4fo1JrLe1iE39LQ51ShaGYbEWfKHmDxU4DTGDlFAm0CBAkG1g
6sVKpOBwVy6LUOFUYiNXwfHfumqv/jjY9h6DXhvblIjTJ3S7bYhjVE8+puDPPFlS2okInjwAgEL5
/RI2HUY3l2ctUbROSv/OXtHRTXKhtR5BzLVLzISf2edtAma4dp4FKg/yGkzBi7ijshMqX8spScdo
6ipRanStfx6gs3HleOKn/3idj4iy+s/YIkXZQCpI/0/k3G37ZMPHyMjMdLkpCaxUY9rhSehi+Ep3
VEJvACHS6ZOsplj3JD47V5cPZkmP3zhZzqrSd8SrU33/XnPjdm11G/jpm9xJURVqXJ7eOnOxUv8T
S38P8ILJwvqmMtm/UrVn9DTsH8xRksU7BvupDMu3JJ9NH6wLlPIDXO2FQvXvoAxLJi3fQ2M6Pz+s
33tJDWkAfZYDkEBtg0okPjj2fuDuGCZ4MrxriMbQh3DMLs4dY8DvhsewHY3C6Sy3ALWdGtjOvA+N
EYUKn8pm6H8VPWwM6OAR68S8VEdPbSQ9Ppj2rI1XBPmc6eLG1IbfGKS7aKxAT3j7+ODNxDVbdzbk
R4V081AX+wOq7rWavSyOQsEgBOjCHncTBZhnMgiOm3pqIPAshgaAThVSWUCm9FAoKCnK/0mneA1n
YMbSeTXq6vvlBppSqtmPsvXpf2+qsMQSN0aw0CjpbAo98syY3wNcjEc0m1G+O2f6M1c32c8dpMfR
bq6hxaxvsMQGCwm7xDon6lDpkGpcMIuYdWPaWfVZLXPPfATwdp+QXKi+IoIQFgyS/FB6nv7zwmZu
mNHnqHOGU0uL5oPokc27AzAHWp0HuKNjhS85tEsxKQnxqsw2NHmgEyS3lnzL53JyUzUeerKWDjT0
w1B+JFzuuPFrZCunGicI/ChPlcl2PYxFGiTO/+4SlPfhtyXZZNBqgCMV46r1ekbnfF6luDGJEVjM
vwiaatq/8xnXXJlJcPX9Ba/ZHV0PVlEIZ3Bng7yJV0Y63NhF5GUgK2m2FfkP1f7LAHtSPsheLQKN
6THiy3hX+wHyRu5UlQ2aDjSZEb6XbbcWwVLoSEyy1aoX0bt9Gl/8arKSIdZiOUeL8cGaIlKOPYKN
dBkjinThV5yHeCh8oPPCaqL5rtG1qzbn65trPStqAfX3fHyIKPbi7VPlcElhP0VeJZwDxj3z5GTz
Dz5yRBbx8PR1xBk4cwMtHPmwMQ3q7Fj+j1gkwKddq0SpARavIKSdbuY6iT2exFiv1uH92XpyDdY3
INpW7hww5lKVpE780ETTTQSq5RTFyJxXna/oS0NYtEuiLJ1vcl+cbGskGq4/6DkBTbWRipNxvl5A
s5T2awNN3AWnbBKmb+OcWn+Uv+5d3pArJRoGl1wHcT5P1Pa4cW3Ql+aCMhFh61+ebSFFFHzf8w18
hLyY8gtF3DOxJrxA6QInOmOd4t5ozRSj6KLHtLqP6nbi1s0aPYRiQcNlf3kW2f5zizKuYL+frhp0
19qJwXrw2WjGrLfdkJhJzOedqH71bBT4oj2KnqM2y7scYKpm7poBv60wUgRZMpErsvKaeKayKYtx
FSuqUpHOgnOXbP8QMuTbd15M/Xt5KZ0IL9zKDjWV9MFehYWOS/QR+vuZG9MJ7OVMbCVqFttV4VtR
WpgSd/WcJXbCLHIWeN+BCibpuE5ChvOneognEnRtddw00ImqNZCqLlJqQJNA2N3vlZkQf4GMgyqp
1Am9lb/N3YKDMs0ukmHY6TYUOtNeVKW4Nb4/4xGNo7vGu85q0ttVa1ljGNKh+iPY6hUjTFRrVwhR
hKKUhjqFbOXYNMDkelvpICYYm1dHb6sg9rZSjLHZR87lQXj4gO8XllrmkeKOfVHyZv7AfJnu30ci
YhYgSdjV6V1rEryrshLdrreGeTZedNqUHZhB9GGwjHtCtnWEvIu45ggoOkF/B/MWx4iItWVlbWZg
euDsT1c/CeTbY15LYYPn5a9lDnDblKEu2t5n/vdq+RAvObeS3j40LGg05nBDRLAMP0DsgEPCp/Nt
aI8HLgn7v0qA4k8MgU/bGvKP4Al9Tg8kXhLXvqqjIc8+26JdEJnd6bsfS/E7kiAbpcIL6rOTTCGA
m36myhO4DLWYyqakGcxBwZUCcWJY6E3kkTcQkZHoOrMIuvGVFrFYShWu0FkE9quYVRj+GYHUWxmc
9KRmzS6AzcYI8sioj3IV4om/MXXlbIUKAcmBppKaFGO7mMTeCMVMtqfmJoh26oixqP1y+v0bh+Ji
h11vDzixJcBQbDePwlqsZHEkrJUIs+t6HrC+Cto3zE5BTzAJOQCr3HolKBV1awkQSPHNqxph1IkF
kUC/cnbEWKVTQVZ9LhPbiCb+PlLyLirWBO8rrvDJzK6oK3y/iqA8OdQDEB1+g9A/Pry69uDxM7qe
l+yLxmXNgs5/FrcaWzfD+YkbeI0IXsw2WnQhBTxctZyHVI6KDZVNcFK2GTogIOTogpemF9BGddFF
IhzAOwfwa3iQfHGkyW593nwPJPd0Er/lqfO0HcY8A4N9MMSUQdrQhsw9EkfTyp/x/L/TmBjQhc9J
rXZ0znVQIt+LLmCFeMi3oJO/bP/b/tzb901Z22MaAxon0hOBH5EtOTMckeywZUk4G0LUK3Cbx0i4
xUQUNi9/FAx5EkGCe4g1CyPAAT9q8PX1o2opxaF+T/9AgpcpnjIa2knlKz7yAIGW9tjhI8rWe1Ie
aQfWom5/lQ0YVgo5Ay0TEYg0wiylEG/FKy3G5MHzgtjeOYnvTesuao1ER3i+7yrERd2qQ3vh6vlC
UA4e2Wl63NraMdgA7IznySKXU/sJGE2sf3uqDjhOO1LWx0jUaFB1W1caLvvwclbuwhI0jWojvSWQ
GY/GZCqD12OmXl001mU5YX/eUvvCggJpFtTC2rCKkmvd/VCB5fvTfSOO5Itb+wiwIpCO2Xp1wydO
/ptjULLY0UMFpvlrdtZ1iSA8EsHmnvGY2QZOlPI8MhCpzG4kUgESL4r3NHy6K/lQZrViXiv3fiLI
3CQiSBacWPJGq1m+PhTS4lPM29gG4COsRgf0ZXGifOVpKDN3G/QNjbuj/+L3E9Mt+D9OD43RxvvM
00m19cJUlrbCbgnPmY2PtRtVFBD3aMxbQ1lvhA2O5R05s1nTN3ltOTGR9z++kTa/5WC4Iwp2+gYV
jw3A7auaD9vE85GlX2G1haB/Z7DIdi6f1VkzVeMds8M5FFEQyVU3kjc/PwLNhFW9/1SVN2WNjSfb
/yo9qXevo4MFFdqGa0wV6zBdDyaSSKtlrxw8HIGxN0NKsASZH0erRpLa3UJTJUnrG9vXd6skhukX
lB4PZq65OasaCxRri1tcn54+N4tMGSIoOw+XqlAKrO189auV0DeQhXobr++6+Iu8p00RlsbTX0/9
sra5mNpC0u3PVrLDCFnba1/rI++7JmynOhabyo0jsYZqThcW8Jtr9FKpySXGRmE3vcQMeTd1/Bj3
EEXhPEADo/qBQjqEeJt310HKOfg4TYFbMWdODvbwzrpmOkmvRM6lhycwHPvwuZVm2ERbd2Ln+v32
MtoSYsr462/qK0jbEocWWOt61HD65GV7S1lmmCzmLT2k+mtBI6DfoFw2dQEv0b/MCFq9Wuc1m+L/
QkWQJJmusoFwTIhtAmXPdG/LIn2MqUpUXmi52g0kjUF4B+H+uCvoefeqj9AYd7o2zjLr85NcLOv9
wKDtQQ0KtQ8k6ZALKLj9uxxzsqvqOynKBkLAOfLGMnrwwUUR2YVW6dgNPvw3va+yIjRkIIMsTqll
iJFadhU+VRvdFu/TOZ7ZTK1Wt0yohz+gf3tIQdrZ/tZuP2X+rHV5SfseuzCqvcOvQ05CLonT7ZCH
tUkX++BigiFS/fcTlwKLN0lVDbHVaUQVLF3yLR2Zzds6snZCCUJDtZScL9gOtZNTk3YUkEio4mEt
6lB0tGOYrpLqQewOLne7zAvPIOi8/2g0w+dN2NsD2pSNzbcuGeBbl2aeWwiJgP6uMnuTXmyQs+0M
b5xPGRigzNk6fXwbcLFhBy/PUFfGzAJOAYAb+FbY+NaRurkgjCiKMVej93KZMndw2lHBiieJ2bbg
6QtDeNsQJ0TRrJfIfs0CrrGsJZEoebOwIP40y/p6vnMQpLQPLd8hgvc0qup4gu6AVJfsOpuw3IG0
slLeRHraBOirCe4RK8Y7GDEoMmqBXR4390VsgTlKZGfh2zD9Z2G1ZK6IQedntfHJ+WULwS0AHQWA
/ENmCDpmTRQhUxysx15Xgdam8r+2cr3U0+QqLAL9pFse8hEnJINWceIOwbQwpX1fYkcN/f8QeXoh
+r1FVUzoYyzc1r1m9BLO3puphXGIBAfs1jZxmB7d7nChzZc+KCAifdGphz1FZ/kRT9CO43k/RxPC
ZCv3peMSNnyy1z54stvm78ISl2c9VfInEjMmIF6fx0uSCrCsEgBpRQBKFa5e2SXxggEBG33g97gz
ohr9RrRCH4j3sGOa5fvlK0yYhAEt4pFWHhosr3OTI1DqNLTmAf7F8/6MYdFD5catELUkwDEaOLyp
6R0dmAhmEeuzYKxh/asELep4vno2BvgynYJwMewG6MPNxrKDNpDVsjTTshCSEM9woheywJMjN/lS
YFCByfHeb1P/VyntXvPWC0hAwCutq1z05nnIpKKxJrVjNGdiSGrKNgbBi9hDyfh/k2XrAPr8sLX+
F60stc18R3FNBTNIwqhbY0tStuhBJ1rh/+It9QLltW2zM9MY5FkIL5g6bFsP45GjsQyQbeilwCoY
Mq3T2JOVESvVhY4PTw+UMcBpXCtiLm085RbVYw57rEsuQ7Okiw5v0ZTjwgDSMQ9FYawK0YITQkcs
QiMBXv95UCjXPuMMToBPQEsLZmS5YcT4SUDLjZS4A3+LR3Lv9a4EGrLNZKKyojIzwbbFh6jMZssd
FA/XvGA6j/pfRz1D4tBcCIu81fZrmBxCoNbaIbsZb1I4/AyrJNeBaS4eCYjyYvkqIpN6rVVS1fl1
pV+Deqi+r82vBah67vF9VoCkDuRnP2BSfVF+R6TIp/AOsQ0B56/BzQO4X40470uX5nELitW5/0kB
p7W2CeAdpxxQFn/LNaVyK0bjaxUMGGR3Cv6jhu2n9L028cGc1c84P6tw3Oet7GxaJHaMhI2xHufQ
NCrKgtMvz7FxquLSj0qkkKHBgPxlRQ0H23B5jDslsFDyO9hj7kzcZRcyO5qIrUYUJgO4lVhRH8Y+
nrE3+wAl4YTxIkzqEfinykKZuLXBlSZzi6a/Sq685FZoipm/3lgj76LuIGKCE6Fd9tHdp9lHu1YZ
FVqXUuD/WfP16LbL2Dg9TIlkNsKRQcHoNLIKWI4L4JPRl+/2grGvhYHRkGdCgodEGV23v97PqwrN
c9mpjIF3XIExxwmBBOsHGTVkhQ7enRxM9g41EaEOgrxh6IkXsKQeEu2VS4ZcFukSRGo0jp6s0n5C
34f1nztOSS8mkgO9LPOiPYo78xox1FeUY0xeOjjDZkK/C8rtHk2LOVcuxiVhgSemK1/uJsb3mxW3
P8UDGVOA59SssDtTAgSnSt5maKNrqLVzuWjXw3E18OimSEd+WmAf9s4wxmS8NNHikpVh7BSppwEd
CQmO2LWsj9GhbhGV3wuYJEn/7j0bS/njp3iHg9qgo3Pmm5RFDH/7WG8+wOZ0UqtjgqUuDNxnOErT
+IRZlWm9WezeQ/iMYo91p0IjZWlh5fPw6nXvAsHTbqHypPw8vXVRAqTpGRx2xI13XR3iUi41UfE1
BKFpIgisMhpa1dlfmO1MWvMGGvpvmnOX6Dx1SitF0KUw+cTjU/wuzy12DNxbwqrcQMwbwkedeW4c
Mr0I7JAFJHUC3vpbQbjoqj72Ry5IXbz9i4HLIIvFgeNbcaVCdW6pRPRNDd/oVSPlau15vtjDbAAW
989RcUqggJIJ/bVgGnX+6cnrbnnkfwoysHq9fYnC5hQK3hG4z6tIC9akaFTzRmsj47YbVc0dQ26P
I7BJ9I4euTZtyGpPmau7bpPZ6YILxS9YXjd3K3fiDCRhZGqwL0fTEdNiHpYL5evm8Zid5EeGOAUM
3z/yTB5D0CRBaYv9bAFDYbqM6gdCQCm373keLtJRNIPsBMhZ56U+WZmWqNUn342AhlpOtW5Lqfnm
pAPszw75JeUdm1TXanNA+jktvpTM/UTVaWNyIgkR8PDUahxnDPgp3qwkOy3/01HMLMyXbYbRCiY3
kD64xMrX7W0nUaX+ZUIb/XRTctS6ycVg2Gwkk4iq0lKbKmrn3fvdS3+LXN2HE11yaY/fBbKNTiv/
brTQu1J2Iwj1hSRLxhj8vruQy+Q1mBH+7/DzdngMsm29f7laT26jF9IPYXwb7WWtZq9OWZHQJ6U3
pGrlBshzNKPakNKuCgApGhEBJRy6Ki43qGsU4jOmrULZTGQ7USSgpBI7ZrYXsSjEvsprIP6Z0ASr
FWJ416wFAfoUXuBVTsEXOsQB9l1reXNgCcWDeBtKoaF3WJyZypWduX9dVdeG/EvB8FvBHRI70z2U
3d7vTqA0iAGX4Zz0uDEcq1wvdds9th66a8JeV/HBzR1j4/yL2WkAJSy48yNbT1Efuqivm0z87U+J
mGTZKjw4kLuGFGLdiDyywIj1n/30NQn1eV++GOcyNjlqnteEc6L92tXia9hngxfhGKDh7ka+Xrk3
eCHciWpH3C1qKH1Nbi9oVpXmkrIirW7QZoadsy6CUURtAmcgLgJCuoeJwbJA8ZlKu4Jqj0jDpT3D
9CKepE2QN6dlYsvadS4RqkO/cx2h+OoONzEbmk6Sj41ismQ68M3R5oWk/q5JLUTEKOZEr/zcDPgh
TzTSyYFzaKtUAePleGS7ISsZocuE3GMp6FgNIB2SI+JhI2ySq1tEMlRg7NOTadZzDkPwXF2ak59K
fr8053dWmaHEM2EdE/qJ7DzFe6oBXV/n/C3sHOcb+JbRgP4yVO6HwN+L8uQI+ZoM9SfmYnU9YRBk
BKeHopkee0ttrkfZJ7ct3UnbShCBzgjzm9oZHzebm58pRbaiBYODr4j/9/A9V6lzyzTjKnNObsak
o7hCYnnXskWq84VdyPS5z2zALyJeaRMeZbrJwEDZL7d61gYb8cFiDRSh9mXAKv4zdSZb6DamShQi
Me9FD/emqw9Egiv0lailoKkfLkE8RCH1fsVMmdke1OFD415dwiSde+rrZ2P4unQsOYtLcrCIuLNm
tAk8izWMyowGODukqT0wFni74F+dZqLJBj9TbjNPm8pUgvXSpTt6cyfNAXDrXQKbd5rTowQn2iQY
pZpRB30A/ec+gVhYHtw9pW2FjCLkzC0OKee56qkrYw5fj38eeQ4hTu4Hk6AFsmU7+KYUBwGsQjZg
R4zpT2jR4AJJxUfStdHcA7R/tSLfHOpr3bKwjSt7R6ydtO6+fX8X6EXj+sLTV/BxglDOuq+HS+xg
Xpe66oBiPmWklohRn46vp9ey71LO7gdjpY96NYzH0zhrkRWQmHOq9RXPM1m4fG4EMozr21vn0/D9
eCyxjJYGe5oQ0RCyKTDmgpHQq1fw0nxcySyxBtWrlQA42tbqEZhMXQDXAYO8kodKmfrD2r3fO2wB
IN16dKdciV/viPpLK+J1EJdqxl4h3QHCrpT+IjfEoRvByJC1RC9/VHYUazEXR1/0K6FHFyCmZ9N3
HxJbl30nhrJ7vhp4vypwGwrMXDV5QtpIIpVWXnPvVzuQLhOaS8jgVfZp3fl2RcPJo+u2uRKUQwCQ
B8Z805Cgt1aOya+y8pBrq/BXJx9JeZFF6bfOq276o2c4NHLW29tGiu5k1aEhksTr8nJnD812HNb9
jGDDcYspFMqnOaOu9kYuMq3wtg3XAuaayikXO4x1P6rTuvlr0ow52qruS0gsfZKN4q3m5UHrPgjn
9vYbRlVEVJIu9rNiFpGri9uJiEBqki1eH+Q30fJy0UAq5xs6ZlGeHUGq2Q+ucX6oI0x0EZwN8FyT
UnZxClKIvjo/EUI9pccCgRYhkP1mLIICFOVv2OByv+/DBF55+LNI+VlW2ssZQhG+X+jaVJxF4hLG
3UvkRoZsA8swg0VzPVNxMIK1SOXJh7i8MRVkmCRZDkUAlAXbYSmj8oEBPGvYIG+P3vJhiP4cn8sH
qGUuAC7d5vu1dL8A61/Uvn36gGKdpPIkNzrYdKWNcN9oOdn98zbelavezDo97sHhYZ21kzUh+sUi
60IVj3kaQ5JXEGKJpO/SJdCrFAlMXtnktcsh0Thm1c26Vt+6E4sMfbndkm2Qzs9LTh7NF09h7WjB
msRt6CDIdE5+NPaHXsvzMo0tVmzsaQeBXoVSpyxb3RE5OzbRTwefPVaq33n1nAXfFhrisJzCBu5L
uJO/yV+EBDuHwgRZa0LxNE5wS30tj3bRlPka9dvoW2nLdIAz78PqOaRXt5Sj8nZKBOdFs4bf0WId
3nioE5Ok2TF+qX+eyuxPRTI9xgeEVsXocx1xZ6Pt37XFccuDYXtULRuVGY/seLRQNQOEPMf5PvyV
KeoWbmKCW8Xdo6cqfXgF6BOyv9gs9/2ajdVtvoSJhIj2q7kFNEPfsmCZF7N9EOTAcG9WRYPhF1/q
IUZlgL3sbZJIMEyFXQAF4FeWzWG6b7uTlEEnOFLULCv6VbrD5Bb1ZQIjDzkDyd1corn622dcBmHy
13YtgCHunWGlGfjMmZzLFb8VR26VUl1Jj40oKyt4kYYPa+mCIbkSovRg2/TNVe6mzxhMg8O2nLPV
GK0H6GvtP9c2sz23a1zxDqZQK9fZR8Wtc3oeo2hzU6Qo3SkQoXBjDeRHeA85jI6apfHeWqRiOPFk
i7pfdnHNkKgZ1+DJQzV4tCJK97346KrXOWhFeUkKEn0Ep6DyLRtH8c0hFL36J/CbAm89iycz8j0n
rAskDmVHkTHEem/FKrs7w30PNTZbJiRZobH1cd/h0WoH/xaxEre0tobKlDI3IO5jIP2xdOijbFzb
fKxgLGIMhesjrAzlZfj6mwDKWvkHm7JQ1Cr+CXm+j9NUUWPIank3v+Xezq9TLYtnwOoAg7vRBRjj
0QjhZ3A8hrVTwPDaSTJf+BGcwwoQIGGGBZ2PaEpCEg3qoSucqthoa2vilkohRLbYN3MzfrM6JvbS
bkhNvQK3+Eo5mD3uvtCXO432fV3akvGDC3qchkuaVBDRhUppv9su0SybFYmgBzy4xCiK7jpeLI8r
DZPi+C03YbpbXEESKNo0z63zCdfu/s3W56YrooOKo1k3sOBE2HrQhJVL29gRwwOYd8HJQqjO2JX3
6TeDNKXjPVznPFsMXkEjdNGiEgbCxmgo4RAzCpXE95mMPiJZJVaBeo0+vKNfa+rAC1PJG5jXmsil
T/6EejyCcCdrKLZHMMtJsEkBPqBH/HVCOi7AQR/nP2tevwrtjDSHvzMl7fsAvYDVZ1KjjKAbPnJO
5ero8+2uLif61lUz7JRRsfYpnO3boKXHWAiT00SXAGQFaTJ1f6UI2m7M6DExYEvshU+T1tuWq+ep
RDou8rBp59Z8BJFaXHuTBwrBR50LBvERJABSkGo56i1cGOvwx7MylFd9y0LUP1iY3A35qdu8LN/y
puArVeZEz7LMlkULjL+wNjkspTQu/ymFaJVQIEWzjdauLmduoprFOsSuumqGqcgqKW6lXDY6i7aF
dx93AX5mzbNMQKSuj+jb+c+9dG/Puu5tzKiXcJHouTWY61SU4sf24taR7uZG2c1+EIqErHurT/XK
QCsJLaUVc/rTLgYdApwhrP4yePU/5nln6kSt+LwkPWoUH2R9qeeJ66Dh1LOUnFjSOMprWaKPStDo
iIXg1XzGU3qiPVxYxDOBX+aTeVAIN6UpMwx+V5fhwthNCjSFj8NoiP4JKVHQxY16pNY/vKC0U/Es
JE2k/ABhsOYMBjyob43UULC9p0zueiIZwgKBAVtudv008Wn7w0o/G54vlW9W/VOoDj8Y/Augmduz
opXzb5mfxBJ0vAqhGpkIzSCEZgNWsdymnY8jrI6hLrdgT9ER04kSUtEhVKASwAmt6/MKgenkT0AW
IeV0ts7gE7h9xMcx1Inxqde9FBW/y5EjECroUnMRaHDABkqWhZJeVmt54yHzTdfj87LfD/6/ZKv3
01eecVVeCWex93zVCxaMukH+EFzTJUC0pAt+0KNV51gx3w+53AeaZk2ARieJ/n2eJuPf5DPx37ua
Q8P1i/JsrWu1jZympSz0XGr19ElRKgsRaJDbWjXpRtCppA9CC/cMtYjauotOMqtm467AiIslAMxh
WFBZzDnKajP17cRz8zcekJUELyMnITKTjeyDh2xYMo4XVEoFmsYF2aU0pgt41nRbeL/Pvs4uITWv
lLhF2hGUEck04oW0kidrRq55ycXb1p4s8kVAIUcAykplSilzPfJQ5aq3b3Z3KGdt1pOKWeMFypdU
Y+RubPSwnyrIIQgrEV0ZOPvKpmOlEPDf+ZG2K/JUQvThqfEJilFQtoch/AljO6ynMCbVK5YN6d2p
pC8PeM8Lgh0Wt/fdih7NH2ULZhIayHC97VqD4MX/gd9l2Q7btrrmRhu72hizGWZe+xNS/BbrgYw2
7mZoXADYavZsMHdNLme8UIg9UPTyUMSwb2t1qNwdib/2Doyuyaq+mFYPusMNjXGczpIXHLoNVpEx
UIqg5wA1ItSZJNkieti+CBHT9DPetMuRYuwcoTE3Lha39Yoi6nX0TD3rB7OoHC61SNlduJHLrJ/+
m7c35xIycO7DELT7sbqumb3ZgaPaY0WWuE7S6NualZ3GE4YwgPw4ojOcv3r6iuMSow8W+CSzCYZs
xWrAZtpVmxvQNPsFqDD8IFJyjNg2q2rbVy2LZx+Oe2TUMCBKQslDTepXk4dqJzixChinUyFjNh5a
xHdvWXJtEAj3VooGqOAIhCGP2dQ13dB3ZxOr6FEhV3eR3OpGtdTH3yG/LUdoOD41aHk6oo+kvOMv
sKnT7QaUiqsnApopwV88X2Mift+tj7X+NMXRdhuAmgJUNidGb9FutSKacojWeLEw6Z1Bsa9q88CX
0O0IePlMziB76LvNVng6HlwQlg3KjjEF47F91cY2UCTMWNapY//oEbin31kkYT38sOnjKGZi9VW7
L+VO5/m/Z/PuG3MCbUlTxnQeF+hvnvvp9ko5rCXo8eX/HCFOPSGkO5F2mFBtsjlk+eakeZIkX3V1
aQ/lVPnq0n7+i/xiLpiPFSa5HxHl2H1XAlVtXuKjWmjLsHqyJNKUutQjD+fxVRLQfAusXwX6gw3n
yCUcmEJoA0D0u1x5+oQZa53Xo58M+Esn+jybYoAs398fqksPbV0dG+GG+OdPpr/I4E22kwVpFWRR
jYZukainBj6ogoWRKMqrOp1ORwlSP47lQwsRxAv3dzL5DHbiQx9D1wHOr2+yxdiml7tbx2yDsG5m
6DR2pBxXLXm+LFrNjjMa+vzHyPhjyjnwS7STIkLtkG208yKPx0OQwtux5zpH7L4mPgmMDEw7b1Uz
TX5Tb2GvwChNkWCvRtlpSMDm7X30WYR+VUECStHrKiBcdiFmpxQDG+RJ4H8OJ6i1iy9+0VF1xUSy
u8u8G1uQMVpzRmlZXDjw+6C1d/swPBmYvSLk9nQuN9BcfFWrx3YKFjivb1u4PyF7FbCiSgdZF1Ip
2n4G/PgkXEfdsp7FmhhSogi6CE7+btYopsHq69qzW68W9/j+K70L/xev2AjA4i7lVEVwBpW7EA0e
zCjBE6nES+p5c/tL65mTpVec7SS7Qc8qJS7oOlsuDUzjLFmLRN1xLUpZFD3tI96wSpG6szxX8pwD
/618W/AZ7yQe8Si/ipc1FnNfGLU+r/Z/7h+x9ignHBOKuB1NVmXgctR5OjvghBcPKdxneiDZioKl
L7THvJEqeYhp/9YFhbevUQH3YCPofmXWAr73CWkEDqW+Jo5P/f0pkfDpAC3KHVcZ6nfraeB9lGev
W2OCRIda66/AhqT1SG+3ChMq+vB/IWKSkClbHrvaD88HDv3/cY+PZ3lBXbRdHMJe1f+EHROnSkTn
07tsJ4zOMVU8R9dzaIJ7/ktluE9s/3hWuRCwY/OGDAocESpLV7M/jbTqkKxFWRcFJP+FBqcXWlrE
G72AV4UWkqkwv6HVnmHx13Nn60dnv4FLGW5n6yayc7S+RZmT1VclCEXAFmISwyBpa9cqeMHwY9aQ
vV9pAgfZle1X/wBf+kwa36umRpvq02HUc8R/KobbnvBvMV73LOz/QU1+uVTxXHFICOL4lvMZlcU6
A3Wz3LnLBF4sT+qf4u0XdQLgBmRqAi6GjihHwwlUE6PZl1fRMlrJKf4U5uNfALgNNB8djR0FC6mS
vHZpf7W1lKKYShRYAiXUbdqL6RpFgATLt0/nILvtXqAEbBMRZKMyDkIHqSfirN+htuCzjx6JpoEe
ql/gxxhwtKJM1PGW76B9LCh2lanz2l5WvQc4+bdoVeTKzfqNypCNhu+03unmuH0DrqJtisBGDzel
3HG0DJFOL/zXPgCYod6Lnte/3JcGSe7VX0/xRLpOSWj/o71X8fZ2RTS/0PtpF69LP8usyKOxllzI
oMigWXaYIaqxBglioOdfwofYDaiZRR9IMAlzpgtuIp6tZZgTYQpZAQ8dDBUqwEg7ia4/h01tIXCz
eRmiPEQOepvdOLphPyCDli6LGGBaTUQDpP2SQlRIC2kgY5elmA4zUKAcgEIVzp8qIbSKZoa02Xqz
lqSPkPnMZbTN0O8MwzUmkmyM+njGf2gyxZD+j7fsLFMuJ2EDdMjtRQ9roOOxdsXs4vZTpSI6aEhA
iYuhh6KD1siF8zpgB49xTytRra/03tzg5C3Krbb3NADhwn57Wy0k6FVry9dv9nvbYbSvIjf8/DA/
YnouxaWyAl610rTbal4CkkHwTP5dknUuy6hhDEQO1Ug/++6FtMXjWQ3whHavwG1efEcWntYTTikL
Ybob2seZD8o1tJ5uKM93erstZhdtxSOpYPGXkeiDsLyBPEUr+Ii9ex3NZcBjGiJWYMFOoTledJe/
+lgPli25pwm/0ukBFhN5ra+94Xp4ymFEACvzzU1GHffdbdrqKH/kfHIPNaprXPvSgKJWoTJ9gCY4
XddMAwzQPnTNjTfXxxj79IFbXzV47KpljNIF+B+ZYPTC0icwbjhyUMRgbLT2f/HuTAAOQ9ElmNAB
9YMUK08jQ+LHHFIOxqrYaVR3HYxC5mt0IVGmr6FdRiOAKC03YszkMakIIfzLg9tAPHF5mU1FxERV
Izfj8fJGzFWAg9t/KdFgM7TGF9fxcZVZgcyReC1OJeedx5/qCRVZ5obmBI2xQyYOVqTOkgiaQBqq
4c1yWUc/CXUk5V1xqkJ5HTvrjbGapUhZb7YFuAoqMBJTay0BWWjr0Nhxt4Rvapme3SQtnaO5b9UO
4jXPQx2/yW0h7bUV9s0jX4wyBjk+0xKEF6B0mBSbCvpJxvVa/scvAPkhhanIb4A0qC0M5L0zdMK1
uOmq2vancTCupTx29dSzf0fmimYxyZ9NQuNVNFPLLJkgd2D/dkY+h6T9fGtwCaYrOpZ+NEuFrwNJ
A9+yAbhqDy8jFknR94IjqPS/pkjJPIi7qE+5aqq+jFG0AyW7AFhSEmrIXNkiQoirVX5WM3rKQbSP
SuNIvjF2KFveYTbk/jmQDGnNUt2cTaUTZ7aUnFG0Np46KP0jJgkWVw7BZFfKmnl6luIlQ//KlKn1
GYFROkaqiJLx/O1rF0Fp/piDyzLl854YWrOFIYtdm7rrRtcPFhctm5/4bRLPnGkblsm3i7kpe3iX
jqQvUdU0UU3jw9rMG5p2LkBh6EoHxL5V8Zd98W1DR5kzZ6n6qa3w0GHfGDqncVUSu/APOmRN3XZN
avwRBZxvQ0pBC61Cw/cbezRU8SnWqCr2W9q0UXwQEBeziWWVUoCvowt7eit84YI01l4HoWtLEmC0
RKlyAzzaahezzD6GUzemkeIYpTjJWJkGoMLAR3NiYnFyPj4tWYn7AuufTc5Jp2sUM7qkvHSeFcx1
Xb3eQhDBW5O3du1EGvt8kgQgEsewhtYBGpcd3kmKJOT2L501oZQGeUPSC9JESAE2ITOf2WJH8Cq1
pqO9gCwH+mUXJeM+W92AghhUexy/MHi4W0nD80St835ZqajX3bAoz3p2t2zodD+qKdEZopa+PZXC
cdhE7IpQGUhqX+5OZ10q84pgUR/IqTuKPk1TVTlwkRmaqzQi9ncp+SkbjxPeU3As/tCwzS2Ayc01
RuYhDJ+NxBYTR4ltRyEODe/u3W22R5zSBWLW6HYIQcZR1PnIMetgU1g/sKclQOWDvKK1sSS4py4W
l7wFDdcui5L03/mukwlbDJfPPEcTkOk6kICzHSfsNp4AionzDV292goUYfmG35kauVcwL70XIzN0
Fp6l8vBVv6mOnrl+qTcUJ/ffA2yxbTRY/CEkC6sM+BgMnbA/TaAziJKEg6wBwfV+ovTbVtVvXxSr
mFiyMpDAqrP7dD7oivzhKWt4mnqnCGbg8jQDyutRnOsDIhwHklvknigWReGI4mvpH+kHhL8gLJd5
3sBrEWthYBYoUN8PP3UeySjABZ6dgpg44aRcUYFlgp/dQ0VoacjBjfIGwgYBewJcmPDmpQFhTbky
RBzQvZS8q6p2fhssEeCymTUbcMkmNRJlGTmn4z1rKO4vEXtVZLIr6fskde6ojdvU62FQrLsXgJcL
ZtcneiH/3EyOKCZVPFMgTj7BVyigQrPlVKv84OUuHs1owsWNgLft1DV5yb5tYSFBrq1nvouajHB3
c3FRZDFFVu+YKrMmE+wmZ0FoDqf2/16O95+1Dbywy7eNO9xJf9mAD2K83B8WheWdnC1uj/IhX11J
jI1D3Aw/7ZZ/Qx0GcUaXuq+y/4odnViTXJ+sFQjRRt0pdZgKqc1TnJQ4FwECvioljIgM0qSaKfIf
kX/KIJkMvz8IbZsJ7z9YijYOb6txVSYl62AVuF+M2MymRPS4f1oHXmpwdv3tPrVEQ1dNhCXwDqta
hsVfcF+9a+krB0pHhmN7TEDVStEqLfMdKlzlBzNCS6rW+5z0ppT6J3U48uJ5U2Sood/NwzPEqtiC
4VotchuedjiKp8omhi7Tu+vA6iTR1sZTWWxvZKMy9/mDk8KkYTYeLUWyxd3DFwCKlzTnqpXX8J/C
YhD/AM99xNjs7RKw9gf8AZANGxrOzGEydpSxhAbzveLa00t7NRrX1ybfBYW2SSqb7Dfym6lQYESO
RJ4LRlgm4M7gX9hsN+IwEIOGe6UBPKBzWiXvSuXwBZ/m96hRk1qqsMeYsj/dvtldohra6F8uCo47
S8LhVymG9/8vZoCn14MJf6KGf5T4Qe6cGSb7Y9wNJuvn9NT1bFa2U5RbYyb8SAME4JS756D2fViR
Z0s904zlfOEMK2TcqhJP1wObcCULXixNSeMVEqmhvMXTdi6AO+Cb2lDQ7D2koMOxcZbyUjCEVfbu
jFpBEouy/V6n7Sa/X4sVluhVFYkkA2z5mVSG3yWYeTOMPytoHIsPAEj8cJrVIlN8gTi3l4LU0baB
4Xzlyxmp8qv4ruCy4lX0KFCPBCJ+W4UdqK9dO/2aKu1Nb6qNZKLQb41n7njI4yr6rV9ov5U1UW1v
KngzVHxEv5Uxx8Vk6G+kzwN8Z6NiFpGT3Ebfw/v4w8KMwM9qKQIxDDJU4z+XVPGQpAxoLh5sjWC+
tnyYy1mc9ajw8vQPjXVM5Kq23r+q/9I/W1mTnOPiWOJBFz10a8CH3EC7C2YqqXH8xSOuLYcrxaA1
plPtglFQ9MXWAlYNASqeigrs75ri4Lzmnz3FwINGgvoG+h+N0mxqQFV2JxsWgG4InZSfppXlhEP2
OhcrBF904qp0Usi3iLRC+hMQuxuJehTJSQg3MrCDWpITtQ9oj+EXPlRJHneHzTJo1AIzoGwD9gmo
YKJJP5F0unIFCVbhSLTkzXSy/GOgVzVItUEquB/MaJnCkARZcDaIkCQDuDgdTvHBVHdYN62Mfm6M
fM/Rdo9BCZLzLj8Q+3H2Bbqo4hUc5on39Rv76GYcJSaWSMpmiGeua7xWqsipYw4g3aFYBUkXxIvh
KYuyWlEY2EGmRODwD9t/ZbwrhrLY+vYOtv05UDroXS3CJy6Mz3GgmgNMbwR2Io9UElr30FvIg0LG
ELkPPsZvAWaJKIK4pgbb306UcxRif6oeE6pVEmlwfzr1fgYhFO2zrzkiJlD0GDyZF/QC7/4cGJkL
C1+JWF6WhGydk/A9cFkrTVT+9NkXW8mndCXKj02H1nn7jEfEtpDtQJQeELFkuEK+vISaBjrTPFzh
xfYM3qkwMmj9x0kgBqPeHDtlsCtd9tstTDQ2XNVaY5V+LGp8VlkT69LhkVMxzt/UvrP7QiKGgBwi
uWIWa8qX+EMB4PWCAUFfS8lJCHlA8VetUySSVWOjAPG3hWLv6bAZCUoIwLBvmoz4ohrPxqlFX9oE
Pe3D0TcOk0l0XEk2BINPnXpu7z8SbTC1wFo4+zw9pJ/2Xs8Ywe5kcUApdgrvtP95aXzGtg+PukRj
Pe4N7dut1WRsEyZrGmhjeDOqygsKVCCM4VX2jsX23h7obDeUZlgt4/HOXwmcAyRmGmgpFboZMzjc
aHsNoMVwEXgq0ae+LgTzFs8lybM9m9EgiGMy5TSqDJPyesoY+VcnZV4CnGbLI1kpjh/fCUdOOWrc
sj3WtoFejb/4+am2e0qmICno7kH3N0PCcRWaDaQWIi7EwZIzqU1QRu6NuvwQrCs77HRC8+PvDHlM
2b4fpViqHi5V3LU8A2Mk+Np8NiZLfedY/+SsqvjBCaLJNpRwVBbxVnSGwpJ6P+5Fc9ojjFdGUX8o
t6LHqACpsA20eIvtUjpftiqGjT3oe2hy1d7M10lb7tgVcXCnIFGyoKDLL3hm8OX65jJQQGLPgALN
+AkK1oENkKY/5e68edavVfYafOq9OBFFwyg1fs47/2m2Y9RVeupRd25HRuT0n4Hk5k7C54kz9FzE
TC/O4jfoQsWnjVQRwMjat2MHtu22DchE3v8pzmVhdIkWZKGx9yzFNpnTntdIpBF4a4VABXGsbXqw
4VSxrf1QGomC0UVXu0KQklslbZkwKBEN1HA8nABvsRMBLoDLDy7/lyjJwHBHXN9YkmB39+IuVlwp
szPaWFHttJ9FX2UlazSQrBYLJKFhEirPV/Sr6n8mDUPsJ4995Yxv1/k4JgBv6sNQrtrTYAm4lyv1
aOSLMLmDZhFni4jOoHMKWb90QTt1QJzzGRA2MbsxyAgRZwFj6VNwToSwy3vfmluujhO642gQzSS3
IjkMC7EkC81/JBGzj7Bzu9n7aIlrZ9usqBjlvxFRE6iqSEZkowkgZXLdWAj7QkqosbSq6OLl0uuV
1mgUe4vojGYeglPz4lUw2R6Cd+ASP2fsCNQAA1aQfFDZa4EpImcqeO5jhEOtIqGyNZutNokvi6bU
47U/0cmfGeccfDm+v2tbqomjUIeYVnhZkKM75ADEq5UzsU9z7MravTAa50gGjQF/42FdtQaKx8fm
Alv0uBg1zehoGlrb5MDXxsRuHtE91sGtE3VqfFpomLvkhaICmzAhN1EAALNfz88eeBUfIbXAGqyr
d7JK0RsmnL+2ibsDt3hxPlbw9bMnFBBnwgNY7+nIH/Tqo3QeTJcrbMfzjPMto+NrC6j+LJlS2HLT
VMxEjAV6ueOLe8ncyHwvX7JHbmAZ3xB+gZH3XmawgUwqFTMSMa8sIPuLC0Zk/AZvNuePtgIP9E/A
Orkw49/GeH8qLEOhXI3/ga/tkRe54HVf5MiJNkIBPCyDVq3F2DwXgMs3KOrxGFXX/NOkCqrJf/zd
UXaDyX4gC/F94KAZK+RUi4xFvUPpDzthW6iw1+f+ejSRkV5gdIVRDl3Tis9itdqdlXI7nZLVvnpQ
KwG+u6+M1yBBNnrljUsZchrzALEYEj50ecib72r+n64Upl7MYpXMweYE79v3D20bQ6YEvSICy6HC
C4IY3enUcSH5kUYEj7OOSTCie+IyVZSxpzqhJH7QB6AAwvj9EYP+omLiwXgIi4VHok7SdCNllL8L
p18SzZqyC8Cr1Wtufh3WYpUDDf6q/AD/MkCsBqESTcN+LsFja2f78SWi02swFyUdCfMct52EkGF6
PgwG4c08sjIeK8VbD3K01N3Ux2/yHiyRF9MTlMV3kCyo3uasITQ0CuTQFnpu8UpSTf37poRNmnQM
J1Pu7nuLoKV8133mzToCvtUeKomOMVJUB0w2PprEkUGi0FZmfWCWwc4Z0j+SJz2au0IKV/FwlbuK
V+kW0S4xv09SzLcMDztOWza5j/J2kRhQ+3G+tnaRj45GM9mgFObvt2IO2dpoNXLEqNlsa3YeWgp1
P7qtRQSy75We/NxVCYQVj53r0fVIeX7NlncV3MaGcHIgNN9OFYGLgo88w8DCSvEFe/U35Pqps3UU
GwRy7QqHeVlVPok3E+8jlDXxfG8XcPhq5OWXCWAFP/ygq4peCryqDAypUipbaPm/Ui/c1xeGv4Vf
iVnqXsW7Ibco3ErztlFfvS/jVhOvY7b5DH0Fq7eJB29av8pMr0RsrONUqDi5zSh3XcsDyPJcfW12
ShgQN6elBvKjFnpgX/2rKzb+aX60xTz3MJLQMKov7HIAd79Qbfg5RfySmdiswlu4Ip0GOFJRO5+X
2vzcDHa/uT1vX8dBq8jEX5n1X9fZYFPjdueCuNy18vAiZmlqUhr7K9xdohAzgjXqpa5l5ncE+Dxb
+EarMrkiSCPuyxu2hcr/QXqZSmQ/J4O8F+vFQOzPwnwR9To2mRtXx0/1hRiBJ3pZjk18uDaiMs1A
Zo6H5rkl5rRXoqZrph9aroI5VMpaerthneXqZsS8ManHcYB6bj6CldcEojBbbsIUetM7NSz/r5p1
YYjhjH66Epqk1RpPGdJW5WkeT7+8CLY5KlArEpcfq+11nnMeroHzKVXgUk86vIqzFsXQnKVuHs/X
25ryDbuwNFH1z/tM+mmzXtRrs/R05WbKncp3d5rU2CLez8meLI2MrlRolbCRPo12lge3Db8aH4MP
OUp1uXGsJEb2GZSWL6mFNSsfZ0OXy9ephQQn4tWBlZAhqGur3UwZhzSTZJfnz5dQMA6sXxiwXwYY
pWxDxGZcE9dtKk0P+bm49dWwj/zjMY/uGPqi7H5q5F8OjyAv4V21PhdE6AdguFCldQ6HhnW3EbYh
xSl17Nsl6YRz/VhnnnmwEcN33Ha1edCz9uAeDMukWfaZzq2aN9GUEca9KkW6a7HA0ipbo0nTvys/
rym2kxwpZlSNS5cB9RO1EEL4prgPYvwDwBn57hnSiDvEPF/me0kWO7iXz0AwjlsPrzdDxOldynjX
K+m79FHqnqF7JCnFHYodRDT0cmOreUyyq+glYdxrszR6Q21u6omqe9kZ/U0hqUAE22EGk3tZL94X
mOlDC9gVnkJv0I6AMrwr1sCdxTJw2VKJBD/pPLVtLz8NjdxsJGOp+PCK361eZx6/48fB4eCw0l64
+to+YW2cd5PGm8M4IDXWVstCTFttxWiybK7jZE95SMju/5fEU2tS4t+aSWFlyjiiG4Yqv3Bx2x/c
Ng5fGBtlCTZuNmAsG3x/jmmHZkHSuwGmNgpnTGa3pZzSHhW0OmaGlUYNtEjp/pbp3ky7nXGiIA3T
Tc54oYGQjd+2aPOUiHWQwkNCKLakwEmHyoGHV/ZeRc79HmV8c5lb0hPwzzlWIzMpWfk7A9IC2+0a
m/747e15AV0VJga382j9FPWH6kpXWNWI5MtlLWdoI4Fsvft8xVKYTmuQIp1ro7b6u8d+rR285D6d
pZ62KE6LMumhdgggWzSSAWTcSFnCfUbuVZ+JpF9+MkHNc95Eb2LALb4IQsPUco9H2Rlvjsb87tVy
mO0hwFZ2iQidzKqmCEBSvuSiaQ4u5JaJt8L62csOnvZ/wFA8SzJr0yI3cHzet+8/x7SlZ2ltd9c0
A8b1f56X0Gd8jQDTdAZdTURs3NNs94nGckqvz7aO+9NuQtg6WHpbBiaMgWqi1vqEwH2pEXdYRO37
gaxph4bdzB4tUBFmfH4gv7beDdBLav1qvKAoXsJR0fG7vf1FpffIZAig87nE93GLOdG0oltMuA6D
PEOmLhl7fJZmnJp0IEenpwIpH+IlMKzYQZjvOqhibWobchJFb5HoYfgt7LIvHmyNA8SLLrutUmd2
MxqlUEcfHQF1jxMdk6EAYp1474OTXY6y05fAfiD/PDZssGCr+Pg2Ggcuwq6tJMgTKfikKtybehVM
TBulko7fPHk3IXhpjJ8N8xXlrwBfVmgmQOl0MEHwnb7lue/3eDgc7JXXmZA9RA9NSfG4VSAPyefc
483oQyYdTGNtycDgAbs6RSH5ZYXFyZ//qoftXhLtME1kdCfubMtl4WzqGE0Y5/cWTfstgUXBRXxG
f4XbG3ZnTKtNaMMazkSZTZXv7cUubPSNh7YKNSWyJXyYBM+rl0zP2N0U9NWsfUxZtXZYVQGk3a5V
r43hfDMUc/L7t/dYDoQxDpdOL4EkcGomEQIKLzn4/XXIk7/phQya15rr4q7d8FHqUFnn2y85/gSo
jppd1dKE2eWnJhQi/EH+kes6RaQRJe/EIUoTgRJBKwY4tgfccL8DRpg2tpALG9EvscpNaUGtUUxl
ewLWnFFfurIPdjfkKuS4sMvYAlp7AnZRRAOEkSRr9c6NiEKUtLhImC30FvfrsXyN1JqNrXPr5WDV
uNt53URjJXLQyR/zCrLTlh0cSH6i8N7ec47IaWF26MpZ1Z3Qngyci/jKiQMdoy4ztgpImN3NdQf7
06Zd1Exc/1eEg8h+FtWfQKl9crJ8Wy4MIGXhtXsbU+5gcodjSoM/USXWn/i64CJkJ5s2Cawjrv6z
r4eAl1NZn+memHTfLxKMK1HTS8RsxWhkeeNnV4dzhPVose5O50iaL3Gi+4pmab/k2XJcrH5LiQDT
sHjFiJ/BpZw2lJtNETPZCUuhoLcq9kwK8NpfNxhwYdLtufBkjaMwKu1yeYly113XAj2psDYBOL4I
N8Kqyqev+cOX0SlqtRolb8QsHzinbMruC4ZzcxBlTfpC4z1yK7iXaYG2XBPGJ1DZ6/7ur4NvA/H9
73mZA6INRd41Siz9b5f4sUawnPdslJne2Yr1caBNU0/VzlVxPd+sXFL3WC5/S+x3cEbw7rrFTrNd
F5vRdEniuU4mAkA05QFHd4nz55nsOLZV7Jm5Qe3OuPyRnPXKX99DRX0QBmpfkKbVKuK4A70HHk86
AL1Vh3nQXFgRNC4wF2Tu3TS0+JBWtWskELJlKAkl7tpv0GSWkYwxkPgmZTOsSeefcM0GGH81U93o
A4aogjn/n7vBDmY/YFniwajdFofSWtTjO6iWQ+UBq/SV8qG7c6Yp0OS+vkCbJyzQt2LrN27S0/OL
ohqfxuw8gfnc6dWxlndpGZYVgLdOQCkxc4/jlzT7RN9+V22kgtXiGX6pKuAwfcWNjNXrkHKFT6mk
F/SUmywHIEugsiJ5KUIuW4ZempKOFK6DbhghlCRNEpc4fCv9+LurN7yRRrxnvfDiETKKJ5ebIwFd
n7bUOKjveM0Z7CS3OJeLO7Hd8EvP6lYuOOuySkll2aBD6teCaWHe/hmcyCwo3V8Wg1YIKQpw8f/s
bUQ4JH7Yn/w3tEckKS8dHXtVXhDRWKzGJZA5QBvM8ucRu0sX2uYUD/zFKXgovaOYiO4lDJlzqGUa
wqjkaZTrs+Ojsje4JMKcXvyQm+96Cl/weYr5FQTcYUU0sacgfAScBhURagq5Yt6vwKm4IbwYO7Zo
Jw4Ns3QV1btVdVr5DApwsjhNKMf4prgWODr8jIILnoqDrbn5mh8MWRCDWchVhrKEHz4/R+eeL/Ge
tXL5NrysNbfi88g+Oump9CdPO72p+WSOVo6WSrubbsheWD4v18WJtEToyuDAtW9li+wHiI6OC3oN
amm4MWvjK75RWKraJHGZmlRnH7I3phyEAt+S1kwLVkO4mkq3dnX/oNW/wGgDqvOyB8Nd6w+mR7D9
urHIzOsLfaMpa5u6k4ThGZlqzjY8nf6WEsiW85ZrvnvKATrTe5VUk33aGT8Nd/4Ct7qtrsykCWFa
sMjLkRC0XZBqONqx92Q/mI13MrghWSmrJwQwOe+b4Dnw7WuE34cMA0ZF1QZ173D5Um1CdeIsNo1D
SecdlHNAce+M4F4muzSwGPwNbykGgveABhAJQCcb+pWVf05wub9U1zszMsx/6lckVjDim85oG8fg
XR5IM3YVcCxuSBPnCOgZ3Dc9NWSaWsKMv2D5nm4Lw/WJQCvrfqvk6Xpz99CZfBxGz35Hir/6qDAe
psNb29GQF3kgf2T7crbj8uBS/TcpRTlvRJ7r/WBy7dB0ygQhs8uYIqo01NV3Kxs8MtSpObm8TbgS
48rxJXctNkfDDhb0vqkzr02josddR6KsYYVE3Rb73IH5iE90xdQ5Y4eNBNv3uVH/W/AZnVtegCTs
3WlogBclkdz1EoU1XR6OmNbtvjGNRqIUH6ybTGTGXpk3YyR+4bqicNkF0umWbod8t0HYBJLVWtok
Ahi1iO9qkkikntEXf9ocebr1SIcaJCeK8bPKdl5ytNkbGJHzvb3VlOfIbrvZfvWEojGb/CNAHr0x
UTdYAjogiMdhFSlbwc/E0cIcDxtRsCP4SEuuqbGSNnrPimloEt9WgCR7bpNXKrNZffGPTk1lc4U/
BWuUeplXhVRnSYn5vKFLs2yHIl8H9renHYlD/VuTY/scnF7MYYKPLg/3btSG4r2+OmFjRcGnINM2
iN8UyB8s/hVqN1IGBkT5CGQjtd6tfs5Tv7i6IpCJRuWfBvG2Ce4VAGAshTIHQaT548wn2KtXtWOU
H9MpbOlApCSkQskrTGQGBNNNxAMeF9o+rIwhQM/i1UCKjgW8B3CgRxLPrzMJ3SUBPsd7MTEGAnTZ
x5tH1+CgGersQfrlE17BzocRab6+MGGBHhUVs/XJloIb1CKdIuyD2r9uZY78fdWvhD2M3OI4prVX
ZCrhoI3uCr4hWgijxSJMTL1SKlcU5/kYWXrC4uUP10S0/t6FbcSagvcKJzMeroOp1+3xnq8d/ARA
0z3ahkitf10DkntOyRfTPHKLHC6cf6JfxfntSs0FryFYydS8K+9bOYHccbXtCZrPjkJAmj2kB6c/
lYZh4tCynXJZD6VL3OzHMKHK8IhigsHGOgczf4ZgDU83IwjXNBb0LoXvPlxi+u/0NSfDnkHd/3ML
iKz9wneCy4YW+pCUwfISdHCx8uozhgPjbMDiIRi06mbhsMHW9prDpXHmpl9j4ibJcuw2QNPhlZj6
12cjFap4LEl3eY5wFkrtB7I7pXjly4hvoMxF919nErN8fc81jkLknswKwxmCTi36OcV0j+RZlmCq
K3kzNDpJhkhUlr9UpRWBKZS0AoKY1nXzIH8uznmF2Yobfj6FHCHqyJsTeiNn6QGGXWhXI4je0Gnd
IHKchrsPznn7F1YEdOv+tpYhDtnfYiwCE5OjpCXj7HYjmlj7ULQrk77wwpLgPypoCtkGDiyqTXuv
zLqD6iHyMDHbDQht6yX1f7ltO3bD7gm1h9NfAUn7d0dLnpnxCd/tg3fIn9GzBq2dyF7QbFSQO2EQ
KAuM1afmHwDgPgDln0J6KRE/auTuNKuGUitO7ERSAVIfVbn4VbSTksimYkYTlHQaftP5vW48Rdp7
kKCQzvjbyippXRv9S7bacAG9r9p3B4jT4WBLzKboNm6wdQbMcSwzl6isrcanqm2Itiqco3FhDwqh
jtXA4VJmsNiyq1hZ6+IAE9cn7/G6jdV7yWRh5ixmuRIRPl8QrYjANf8TgfmxEApU+oUG2o7Jj8mK
fzpEDThzWIKqfTdEFFiqfNNg2bPz6GRzY4dltdAKhfaXLYze0tn0GZfnfw4MIzevuy8tf7/5sSD5
d37w089IGj1AJrujdbH7csNqpxdc8VmIOTB7ud91XjN9PtemDa3tmfnLAekHP20oetdrZIr/EoKt
C4XWvGY7w6l9mDndVzazyWoaRZB0DL9HZzvEbRb83wRPlcfDp77JVBdwO09dpuHYYJdoi5xwQV2J
0hwk8ooK+jke+jrTzcE3F0eu7SoVdx8IBTm2uMJ+e9dxhf++CMHhPAlCpQB2uFSN38G1dS/5+GcN
ZCPXI8AT/DVz6IPwl1Qg5pBifMHU0UvsIiZgWy7/v3iYuaBAm2e939c36UE1CzA8tMhqJ5cYD0aZ
eWwLX908rfCCYkPu23WBcOAd0tOKYuX4nazFazhVaqI7YgI9C89IvwSkZkWF+yuXTGv5xA13l6Gs
1CvCkReHJXJ+L5R2f1BPBZVH1HgXd8K9cGnEJFt+hhgpdDGPA5HziiqcszuEOYHPOZUig8DSVOdU
47iapiUQDIpQsAWIl24TWucOOTMqJjv5iUdVHVQ+FqnN90alsGa2DeHI5n0LIDWUOMT1C64OiTBk
awJVuPXn8jnwpFKNKpj359iOdEJp+LQX/UoPN4ame/TwXEHTsrcFC8OwGJ3DHFA4qrwoYz9O/KzX
XPxYtJFdluThxnBXw2d42hm9y5uA0LCR4jlG5UozYosa4HOTlTOvfqKk80iPTc31cJcwTtmb4Wtl
dD5kaozPRQ6GZLjW/CmTzNb5Fv4gH4s3UHahFEdo2Dn9NuqmWOxRV5aSyhhXr8n0X2dvWJRkX683
Owu0DZryf6kSnFGdBf7puAfIXm+MRS+e4MOVE9xsV579B8y2wNdmHX1tcKhoZmr31XGuqUS5vKSU
d3OKwSSRUnQkUhgALUfGRTwfZfHPsl55dNdr36/kMp9/qa+zJr4hnptbohbP/nw/kx1vj1fI4gvD
8VLr0g1jSVoygShXMe50v3EtsD1ve/9jUtltzIK39OvdWTq1yFd0U11E5WGCHGfRGysVsjfiUCEF
t2SxQZPCj9/GmGNGlj47i0KSzwKHAEZhavFMJ6wxb5D8w8PeNCoxzH4a7ZlwjsGBOqfydWfkw4pv
Wok5jNorLo5mCqqkZhRj+dNXZwrHCxVhLyhof4dJiK6VrUfeROHkw3jJz05p4QSSSv1ywKfM+Alt
6yMikFsDMlwgJyE6HVpvMWzErQ8EWdWsHoSEd8grAeZFqlRF+Lr155IYuQuj4KC88ex69d+/dzjE
WVn9CDAqUaWW+Frv0uF8oagzfKSTAevHDpFxvrjzkFgoPcis0xN6SUEYWVh1QWCcFSUXkwPJEg2V
SUERLpa8dxq/jQdB4cpplkn//i06iOXdqOFWxW4YvpNeSgNmYNdYiSan5m7tOIqQMbr2YsrS9zEs
WBkt4LfFIsbrfd0yq1JxVewgOGJWmoSOqC/IhtxqD7R1XhGS/5n2xLUTdGUMRyYvwnCPF2VWMPcN
B+NhZDQOgCXk6L60RLHEBe4WbIqosImX02E0vKPpCg31pjsnTH9uanmvm89fTqxcOcuiEw7vYnbb
jqib0XYw5lBdR/bI5AkNqOYS4emx8nH7MV/XK65OKF10XJIALcEmY37jVJ0tK8+kUIVZIA4YAvJ5
eStYd6UNgUlJOzglDX9kcpNvZr+0BTwb1d8cy1WhLVNa1yS45XXO5sbA3TKvHhEBqxDUKCikh0mB
czLGOKtYRDMaRxHdI53VZ3uFz3oyb+OxSsTPv676qMTA+F8LtB8xI1itiZ1BwncnQbrDjMZ6ez5e
FTlqPW34KBmVn2k5jvlvojTVzgEvaaxAIiALMGjN4ZpHMtz3PZ1PyWQRE432a37VQfcuWZT6floc
guBo9zDsVgsxWdI0KXyVy5Zo43nw+B3UBr1KA3t0QgtlNFLoimGOivBgFf1KwtyZeXMa7MHPc6dF
x5ia1Q27/lE9kYyPbhaLM+kjVEPt1+E2r/S6WW0T6Ppe4K4uDxTJFwij8aTdFLrjsAgMEzD8Zgvc
psTXqZEKj4owUoCcx+PkwBsB6QlmSP5M6PWA3enAdHs8us16AXyS8Y+RM06ptykiokxhZTlNAegu
gML4EeVFPTfCRvVG3G6VkHLMY6HXduW6+TYrQQGQUtYXv6jzWA7PfE7gmbwdZMq2n0IwJuznSad1
Oj91wFZDnkUK1QXpV4Qckcb9S9mx6lDATHACABZyt0QOuHJakfTXnDhlXqyaFT00kezSM6uuomDU
7f8fip8qJs0hPs66RlVlRKpwKk9+EqtCr76J98n2rOSYaSZKOpe006v63PBBT6GX8McZT++gqFQ3
NV6yYA4VyBLPY+C/LVnkn2l1Isw4rsdF34hMWDsShDXlLWMOaKs6iXHylL7AswxCNA3DqyZqoqHQ
ymnuGGnNxVpQbGhnBBQ3TFhWESrR2asJQiBJQsYY4/lXoQKh/u9qNOUPy5qqN1xGw3hlg3CI1bRb
veE/MfXD0mGuBwDF+KrW/woCh0agjXiUgvFe254oqfLNglJsv5WwIqq7/NisrBdlzizAbnTwBHMD
u+OhQT8QHBIb601MEhYg9DJk9k2uhuHjEEyr4/IpShjdP/JtzZEY2s6poL7yJ6c6uAr4R9Hu6Bmb
ifYZYFvXsf93+tBqEfjoG74fUm0XW5UghAMJQrCoQOYdsmHJhv3nOQt3QJwpoSeS93yyKtGsYWBR
yOKYGvia89cLakNvMiT/wI3qDAQ7WY7woJdroNfe1S9BwEIySVcrfE5xQxDWa2tAhIPpJlt2mtiM
L/HXUBn8bdD5VlpVre99tCSqgIjo95EuAEovnNpeeYj8h3+I1gN8erTunLuMYRnSY/QWo6zpZbjZ
M9NhdqwVUNEd8KLyZg0fKZWQ9C9hZccoKwLTxV8UqRogpJQENJJNahqTxvC7mSNGrGA3tuEqPrSD
+CjtOKPd64OTYY8wbWhns7kbw2Si1LGfY86gUqjoJ9vQUsb9ExXD5ziDvgJgTrLunzapz8KrnfGh
9n0IPiAhICp5Z0f6sATzQoPA6cBcbdqj1suWIrFreMNqwkAPyL2k7fVs3ektnljr9XcwTZJvzS+4
njbN5iv9Ks0TPQXgU2voe3wZm6hhAjlvV8rzSYaOlkOXj9Mw9RTwWMTnsTohhPzads5UcqMJyVuN
nn61dU+Xuc88dOjQZ88WZHEfMRhBjayyKVhzRVIdf+answWcuenUm5uNXrkMPpVCHj/wndI5JOJY
yPGIvGTvT9ieqtYbAVBnjBUwqThIE8+vB0Etgz0kwnitcoyMZ77Rd5KrHroKX+9xuX/Gio9aqJlJ
5UA1CcdQ6l+zX2khK2ghnRO85n7dWYvWKQsuBOigRjP2PYREHCdkG5xjMoi9Ho9MMjwVJNQqeAT4
Z5trHjMHeHGqWebsyRTfVlfbZODYkyf0hR58CZaBLZJPJcAh3d5JnlaxfGUXAHHaQ23CBT9h0d2V
OT6Je4lIwNPQv6NXD72/xXz1xY8HG5nhy07LhRQFK/BFM6Lu9+fcTjf7Ybpi4hN9Q3eG3IxKGItK
ms/1t+19tAufwMRAr5Twae+sC32gQGla+Zpc9nPp/ZUjHMak26MvhnYVytBkExRjSXSkGgGkgzma
8cEKdrvH27gVhFUG5tSqkINLMzYrnM5WLGavMpIuT+LZQpCp12di0ot+ZVgxYoxZSKxLqcA2Lie2
TUD4OcL83vyFmjVAAp11W36k0yIXOrpabGcVOSu4rkV5TVkVK0I4z0HB6raBw4BLvs95pP9jJbrS
9L3NMa0zsfy4005v+/sh7nqrby/Xes6/QppyauAoGHK2ne44G/J8Oq0WFGSsgoUmi7NoRkMeN/VR
osCdBFEHAGvyNYoYEMGyzhUWh36dM14gEPDF+48Z5uo1ubXj1SAtuqTJv6l/0UHyYimEi7Ju5Mue
hXlryZCQ2sMtCEUnPppW7PKRFAMyFHyCS4pj9IoWveGaJ3Nb54izr1ddo34M51/r11GhR9MUrQ1V
xW7jlF2hQl3V3gKQ+2Kh2gLWfhTKclnCAjkf3QP12XlZ4qRXx+nh2dXb+CtkDPpD5wtiiqwXe0eX
HYNzY2OmJoHytaBgFsU0crxUX4UIzQYNlq+TYWkAnZL15ebDKe3LCk6Rvi24+R3H+aqtUVqkTnH7
zqiYwL9CjNS4vHXeD6nNky0iTbE9Hr+D9ihALkyNG7GRkgGgnYToDezG3FH03iAKAwaqE02zSN8H
Iox2BUIpiQP4V8ELtY2zxT2Nnefhd7S2FsR1N9CALXry71ySGKGqfOdOMWIlkUH795ct5rO95cJm
Iyg1XKvivknGukyypfwvcNpgljhASahoUibz6u30alKTLVmF8sO7DF1UDjIAi4SNEK9vHpj6F/EM
tJWvdAI4hltU6tcRqiRXyJEGkHsloaertoF7xwI9eP/+fPfiuJznFr/KY70X/aazaw4HQmGGssrl
HNkGIA2mvhLsuBo4iR0Z146jQb/IKnkrSzU6gNrfhCp/+qB99CLZ1AIKVePaN91FrXg5wiwIVd2e
5CWH70MC9cool1Sz0t9OynrxspTvwrVzV5oLoDBlN7TKPsNv0Do/zASpShIGVDnPP6MvMSAnp/lq
dFjWpvuHsS9XmSEgpKCko6RBp943r2+DDnzQUgqhSBm7kVtUgAuL3g4PD5344L51uJYlLf8KUmST
truMy6Dtf+Lu4CwyGIEB1WzJZsXtvw4j5i0SpColRNMUQThH83Bkflz0fb9b/eoy2szsSKYz0HHX
8FodRuM/Zn6mhK9QL+BZXzdhiVl8V4r2CX+5v2Tdqm773CS06vAu/27m2ixYYVpl7HSUGYi5WA3K
mLoUnlQGe5AJV9ZeuRNq4y//xlU9QsR98E2sZ+xdYVFtIgGYiAldGWP6qHEoLTlcudabtjAq+6Xd
gPOo4yHQrX/v4p4iXZ8Fi6TJQwwNK29jjhXNn2V5Lj3Ta5bV29ncrneX2BwMdQXPWJtdRHBFi606
Iwn5SYOPA8zCAN9P/a729yEIDLvOVbD7VNSWUn2aSZwMpcCJ/nb6hskhtnNeypVzeAbx+yqc/XKX
FJPNGELmVtsuSYqfk8CcAGgCw7GYp+swK4oAAQjcD8Cfj/TAIWPUu63iBViScoYsAVbG/bHi4z76
lWWdb1M2T9H6jf4O4bZPeHTYO2SEru+newQStdCX6qHu5dyePu9mf+t3BmzwQz+DcZHB60WlO2Tc
BsO2rj1+CGlo99aFzse4JZg453Jr+SU9cUdkAvCop68yq1Z9TYYz1Ogd/z3kFpjJcA7D8C3aJYjQ
N8QVOEcjKfaksocSTzN/+/evzpMcygXHyInPn65+UfcY8qsXq8kN/bOD7OWAkqRjJ5MErpKg0416
DMX1A0FXpMqurbFf2OcAZ0iUKHlbCDzpRCXDkfG7s56CW6daysDscO/LTjyjxNUuhb4xxNDNjixW
CnUXIe2udpbDd1A6gybPGA/XKwHNpkvsuCgoJ8qZkU97QtEENCsnQJEBMWR0jJbse7664/2flupG
fxnTY2tD4PkOUULmBySrQlebrJwHZW1chQ20YnKvAMTtPAWq6clJeaThHADC2arshC+AZOsrrWN/
eKy2rN6DYRVrKxQHXdijCYAat8g9IXd9s85EzSBUP1eH4Lz7vll6sZ/tEppfOH+QWpql+HPxJrx6
mzLZteXvsKa7h1IphLuBBAK9J6yJtxYlFw9LA+USaWZTbpIzj++G4kjroUqtdwvetiz4rhQidbZT
I7VEEvcpPx5xYcJFBw2bdcUMEOkE2H3vKsBKRF7f7KMh5/CED2T0JfOCKdpDWHhFgz9+bqokovV/
HXQIsy4eyYpt3hA1zqZ1st4C4eHONUeTv5Y6+hWS+fgquc/cy6H+sdBgbfvXcEUazDPKyHrbrGb/
xFa8QqWxKjA7adeuxNJ3yes38aXmFejgYgS4tUSdi+Hk3liMfqZs7KNNzB4007vDZI+jID1C8dQ+
o+j+0PXTlFW4tYH3PC4/dbmS1h7H+Br3Odx0p0QQRlrszc6a5MfGcpvO+gUrspnmNOz4LSipkOw/
gudmuMlpWp6ZhncvqlKkvGZ3I2CU3IgKDwWbKie6FvS8qiLfeKthHCFhavR9DlG2hDZSqd4d1RLR
csWLJCL3mzMQYpcicfvjs2Vw5FMTDLpm31tiKa2AMNOnKvL8gYoYRaI/vlirFZ+7Pxqvwl+ptcQX
oGQxjwoqJoqryrsHoSJeW20VM4f59cSe/GUaygvz8ER88ZIBw32EVdZxdYh+7804ZZmOkXR03+1t
dgS/I1rMQgcjN7sGcOLplztyPiXpmrfHh9TittDXPIZ74yi7o/v4gVPqGj1iLwg/DqHcvYt28A1w
igGyeS7i/7SljJrPJAIE7OIEA3JCO0pkuAoebNE8rPkGZMIbXu0uOYOjC+8yZ7PAFMM29exF+Htn
TNRbvJ1P/bQ1WXQeST6zHQ72rncuWAiEn9CgZrAgTktM88mY0a+MVxcGmX6gs9jp6X2SobespfNd
I/Zkd1cip9PjrIfoRHkOYBHzKS03OCkdppezQVZiG7eT0T4WoZ/bKEzPo6SWdYs7vPE7rjO4qCWB
CMySGeRYetA6eKFxwkQFH2awhwe4PjBrYBjc/ZaEw9ufetgm5dEavddY7FVfFMCugHxYF5jDQ3gY
2CJMJWiU1tJZ7aFEnvz22208JIXVh5ZCWldYWjT4jmyt/zDZLL3homgjpadVMPhm7i+VtN1LYn2R
/yLh2+JgiStidR2sP9ioSyWxZy9Rfv8BgW3zuVwVrQFsUcb/9vOMFKn0xdPYUOhL0o2mXLthrQY0
VgI+8M0AP15iK/LcFNsZO4rg9RIDznz6E372PMM2B+ch9X42N4FKNBz+KEO/vFOXXHPUwe0twB+l
QOQxJMe9fwWeCs+qLZO1nsQ16Vm5omzTgi8XZnxewDmXDdwCkMC69KsUgvMA7+XCmlg1ia3IgSII
8SF6GEl1kaMg8xtunBQNwPVIdQPWuPOT1YqgJda3+QB5c0KitPoGxz5H9xjueasuAatVdY06iEWM
o72hvBWOzJWqJ+YSdcqZWHXZetE8axwEo+MwBgtNiFeKjGH9BbvQpHw9tNZoQU0Zd+T76I1kCtIJ
/xuZY/Q3t9HFAcU0DLRHcTZ3olTZ5PkWCWU1azwCJ7S1SPFcp9lYlg5yYe2hwXl8rEZK+Fi+g0fx
qYvXzgm/l2iUrYoghqpp22NOl+un4P3OD4zccRDF7LNyMkqm27bNkrMUUx3bFUhJkok8GAoFDXNp
IyR4FFzNhtD62CgATNYl+kTnwKzsYJxVp8/CzhemcajIJ5Ni4QC8jgGM9Agnjj1J3oAapRzYNLYN
HWI13CMS6Aim59VfH/YZhDwBDoE+uaycHMMwyr3zG7XshMdC8vRnQVA2JhfhTlEf74Jv5QaOV8wM
Yw8W/uCHAbudmfRjH85UAdE3cCbk6qRWT8pihMFsSrT2V7XEAJDJdxa6GWVOyCqsNxDZCD1QYSkW
Pj/WUR/cFkpwFAqen1km9Wl2UDRiNp9CrYt27vQN1e6Ok7L28ICCm//ZujAlJnmHQ9HhoJXuBxZu
mJr73/8hTTziFOTGpQ50YI/4sRrxyFvHOlo+ED1FLmNnyVbPuHeM94DiFIu7pIMOcVM2NETrv/ZS
qYHgC/NXmqeor4MAHWyJGAYqNr3BazTJgOczt/mFNtQgw6VxLdOmA105ifcOvlOS51hQyy5/BCK3
XfH3LkoSoUweN5vCUkMmV1lfRG3/NbhFJxNiZTLSqCaRFDq1UJ/KnMYIlyiMJ6KhLRf+TzdClPbQ
ITf9sNU6XoDpKOzuY66BgigNvQe+zJ24qbMHb3APED8pS8lpgVcKfCipEh5GKBNU5RdkATJR517y
47Bns0crvm5HjMsz7DhvI9yAgHgsNPk9XwkxgXlNJT5J2n5IexdK0AQ61ToeAztuECa7mOT0q4pB
DyvpFxszMRjIwkdvKevUmo7DAYLhOJC9xDx4b3cw6nUqln6N+UTerfsWz5fhQre3pezH/jqEP63y
faDY8zZwRv4zPNkhrwyQhu1rZdt3aI9sbBkdu0ohuD5GdSWTxJ91tohIzWE728+s6RkE3aKSinF5
idXz6trlu+J9FSegQyxEjxMss2Acp7vv3AqPP+jl8xNJELKJrkJSjA3VAIfCGTQffux0Q1BzVvML
cYLeHMcvnXNKH6J9oJNcjawqhyRRaE4zfvgXhrDXwflXWg4LWwzbGDrpC5pcbsAdBT6S0+qPIgt3
uDEBBh7UtbL1eRg3i5XOOQKsVV6tp+JFK+ATRFS+qwSSxql5uLMWUSfekcAUaC03eFeHUw7l/uld
DTWSWDLeToiF6GvNKQekLAcuV+sflpIxZZueMObWCKZYraYqhBE1wIUU1i4QHXKdVx4dyVP2pErf
lpPSiwqKa2dgBnZTMbppWvKIZihKpWJ7NmsgFcQGdhrNAc/ov5i8OstTno34ZD2JRDxKUJNOQLLi
pgODPfiQNABuhFYZ8cKZdf6AV3q/OHzPZbelISDdS78T81pNk9cR0f9Yq9eDEK7USb3O0C5oXwCn
7G8Vceob5zJSYcJwx8ZA50pJ915Vqc5jU0+qXkB7FBmdkoibFQavdW5EDa3q2uf/8P9IHGmLDXYo
IykbE88nqJwL7oA4f/EBNCwYHOFX9H9RHCGGPObkYqFb99e6ab1XWyZHkQz7VUY23vCIcR7C7qXI
BD8LCa2qRPtxdvi7wzchzkn+TMRuTxqlng1YoRDFsQOvkTKwB4xVCFQ1VVMlhutW5yjzMOecO/SU
an8MckJR/bWhAS5SMUwGqICyiFs/5BuLIP2l/3LOe/tBg/ST9xtqkiVwPaiN1oa4BK4aqg8/shcE
emHo7n+bE+e19zmNRtoSMUMfdfTgvuqD8iy6WIoGzWARri+QwJzgmGYLRujXsktEcFVsmbRI0DDT
eoeLmD6FJD3PE8+/8L1Yev8OyuBgDOYZPb1cxEOQUu+L2knhbMvDxfDomwDSM4nZh1/7iAckxxPm
7xhJPPDf4plt4MF6KyQoapOx9I4Qw7ZUyqoN1kQEHR4gtSfRvhyXaipzos8HQ7j3q4X4Aa2c8WRY
W6onfstmDeKDF8HitPsRSfQhtCL/xVaWndfK5VrsJ0GJcB/y6TDMiErv6D2Woj8+S61wCokNBeZh
q2jbg24mJtQZP14UMFtJf5ltwUqUzPKufLns5vWvS67eL3vDgw7B+SA0bF7ziq1g/zBi1fWd5tYd
zgXv8LCDznf2p4RoFdNLwoXxemcbzUPcugOv5ATljQWy28Jtsgq5IhOFSXQRni491AT4aD5XbLsa
lir+A8cvQGjRhZVaifpG6bkXZAhxBW9hxSjPmrWpgv8heqpx/1PkLagYPNVBFxgkndN55Cs9EPd8
YEcNhAfkIndcdEa6HKvnuhmLnoOziKgM71TOAT6W92IknPV1H/ML91g5+OCtezGsnp/B6CiZgwTr
0fio+qh/xN46R9LcuqSXuZr7CA3a7vvbpJbxRYhdXcVB2/j81lJcoFErnM8qci/4FivnyF/v9hNy
0MeR6+esJEqnQS+U+o436n0WjkU6LPyldknWkH3WOWPt/oeH+PLD7lxZvh+ygksLkgGIWsISj+9k
Y8fO4qO99BY/z8zC8gKIN0y8pQmGvAmDTWsAcGZ5GKKvMtkl4SjxToZ346hvGS3DUEQWfLc9uquL
PsWcwXRTgJjbDo3qo4G+Li0M7cDIfsQOq5jstCjaDUjk+WTXlsZ8oW7hKMuBbl/zG3bcMnnIyb3D
eR8e5JLtHRiR2/RP8pnTcToqS/mdLEp6HsURwTRyxfH/nE4vffwPxpTxG+k1oV9uR/0FKiNU3+9X
EzhP1puqAdBqkm3u9J1hxxKDt7jCi2PgEWB4cl0fBqcdfs0RBBeZ78XU1eiPcvtdNLwyY58Fkf6r
Ztg2P1mJrAy2VNW/pTE/Gieor97D66tttWgncdHpnHwVPCThgaEk3efuMX2WywwqGdZG/hPFskUB
4gjo9dz8Br6q4t2AcA9jKy/Qc3nrZq+4Xy0OPPSBsQhQ/Kz4YLo/v5ATIS/rFTuNmadQbDWUZYJA
9oGXuk0/nkqWLlTBVIfzeUgaXUAjXCZEzpT8+yKD7ILfYWGKmkvl7no85zbJS2AOE7Q2whHQW9c5
zcsufkyy7IXBUOjIPy3sqJLY5eSBNr1qGuRdVIWrx9kjJQEzFh6IrcSICngbmCxpPqO7//ghv4Zt
O+A1rKQY1qSsq4Tn2s1s73uF2ydowomPHNcemaiARSB/uyT0MwByXYcQfnOAiRZI7/bBJdtX7NMw
e0PUZVXfVccPlEzu+QnrqSKRoDYhIjnq7kxXPsOH4nTDV6M3W4+Ei7XAlO37aZGTdESe7knnQYFV
3uRQePv8b4V3dD7Qs9TIcBrJiAIhPfFjDIcYmML5A+FE7McopVrgPF6rsi1jPc8I0jhK9RTR/cgr
0z+wlTm5BApEhVCt34jWeamrm7Z0um3JrAh+2QCKvvxcEfI31C7MZT4vQO7BaMVCclksf8uiVeg7
XZpnUPqwFNLK37++TyTM4744ZX/WE/TouGGhw8SDgDB0HRW1ZfgolK4jDGtgqiVodSg264ORvBPy
bnZCjpgVtXsBjzqosCKn23oGID6Aku2Gf33EDridf5b+47wQmJoDgXusMFiZQZhX7k+TTwBQH8B2
KpO/FANNFMp0MaGVMh3raYdmF3dhSDma2spNFrtIj/vyH6mj+sKWMlU7q9N2C8XVTVxYQbjvsnNN
4x/u48bMll9L/BurDGgDeBULkQPLZZNPN6N6d2TC+M1m6yMvK3GesTW+kFfIQ35xwgJtxsYiDdjS
XMi6bEkUQZAU3Nbz6zgJFWtb3ROeDxPZG5ap0lu+cjq2bWEZhaLBg7z0lSYaNzm5gPKxkZ9KzLDR
y8twedPDQ2cS4qvPR9oNq2lE15moW0wFszmfQS/pORPmKmn3yblKyjBDB9Ea+o1GfjQExsZiUUNe
UtZaOUlaEwAtIS58xxFPgqDwwkpR7RhMpIOLcjUc4SL7g9eMLF/EeLDwRhGRfCZhtjgsSgKUPhbi
nuZMKYec6JhHj0ZQy4zsVSiQ/18peDfT3keUmwlrtB+9FWGmVJheXA712OnK8Cxs6zrWQjt1Gwdt
lPyoDgDtRY22VaAuGLwoFFnHHanGWHW/hUulyOjLT622qttQMSXiExJr1iQ7GRxMiiOjtSOApTKa
BCJSDaefAeNgUzf9FPxdCjf19040yuqN/NdYCN01qvcFjcfxKFHY5OTTjpVqiaT+ZbpIGTv6LeSy
ukXJhbnFZ15JxXx7PY05dpDL/ruYH3lybYPy9fI0CkejUUmKfmhxV15QLsiisuQCAuRil33Uhq8Z
HfX/qgt7tJOq/+pnLG+sj1PYbPOWkYQXFzkRoicHrwswzvKN2MrUyv63qEjHiU1WaSLBJwmi7P8+
Dp447Ub/F49H/fv96f7O0UG1munC262AtWmtcA4o3gB1MrLTe5dOB3XK2BB2B59ky5EIm22mFU8N
iEIKVckiTpu2yQhhgupzyOCOhnMKym3ZcFpPMxCEl6rbtEVch8PIUNqajKyAj41XPnn/Cgq8IOXn
dbwoydKfscF2BYZO3vx9vftQWPoUsq185IK97orcy3VoPQprNQ1PT0hWlkaIoKLEHSgjOwYexMay
9c4syO8KDZh7xo5oQHpK1kzj99RqshD8oX+K5KqaJDgB1nGHZjCodX1k2OWtUHjFjZgFTlHOW42N
s8lUHcy5uSA4/dBTvF1t2k0Hc8VxhplRoSG2P7o4ysKUwEc5/m7t2K/aNKIjsb8b+AcblQrRTs5W
9YupveFxszpE0YWnod44KYjCKRxhut4Z9M+07/IvbmIV/3bOU4BfattUCopwhTXFs521hyIturwQ
nd5WJyy3Bae+QulvVCR9MuQtISjcTaAu4cSmPfxR3ezrRZI0/HoIx1afWTbtSnr8hXQoWqcRSHNP
/n5hoBEMXNOwuQlSHo2RJdEEf9VAQPrTrUIaUZNctu+oCjtg3hnRZ9THJWqhzL9k02MZ1ly4AO74
qOBMd5ayuug+a5bgpLsoeeI+SOZBU08pYJteoOfyyeadv+5WYz7PXdVXpKvirFpzaww1QaPHxTsV
B8X+HoaIHtkUWlCSwHh4HEgSwuRkd6W3d/JTmzs2Ac5la1Biv61wM/Nf1md68qrFEKncWVmNXJhk
K4XUp5ZQsplWhmQNkFnLH3K+9+cbhXX+rPk0H/TuJERAArV6NtwgbDbHNkWvMEohyC3ZsOUgxxNj
hgGcO8DOOrsdc5mFoSKGjT8cm6Y79awq8dVdTOsdmsBweSkmcITOLzYVJsDlB+NTvsDD8Nb6hPCf
AuDreTgfXhrv1gUTcf7K5xA0DRvK3gBNBnniBqf3nvcz9mHY/abHVYfz/usKbdSHn7laBTzw3vfH
zyYt51ZJEqiDiJnyXdX4YC+ukLak/meAIbX0OhVwyCcgWZUuz7yxU3VskkSiA3LEAdx+OdZMrBnO
rInO82ly5gOpr2E3T6obbceob5v0YtmFhP9mDdQppyPK3jXRNeO1yrLz6WFvMMheC0Bc8+kHs55s
/uVLTGBPdyFbDaeltXi+Tx/5E5SJGdOrJRYtrVuJjFCLg6O6VFRXaZLmcnsDtkZbazX0ySj1llO2
V9BgztsepN+qyidpacCCMdwGCtzgCKPycuJdY+cm/T3CFI99W5BZC+VyqARsYNKmbblc5roOc+/f
Z9valc5qIWpfSEFq4o7/aOr2EV24sqhRJEsk+hdo9sbQNCKt3LDETZrRmPfi+F9fGBflGHE2zS0/
Ac/4B2+U6Qu8Ic6/0JMyqdmtHHOdHpNArx32ADkOjsxX+LLpPB8jKoldxIWxXKCCc14vQvcQUTPQ
OOe87tfsEaPGqAfEL04MCKWD5La4f4UVI60QTrD62+mdtYpl6fVbbVmZLLXo/yRnbobfgM82S34c
lzknum+6FGdwKIf51MRYdBug/mN71Da42Paky0TBCumVl+/df307mCtIN1GVBCySxrNOvoVP6NTq
YbX7QPbR7y9LDo9uWtGStXPj5n+0aN/MZ2UDs/ZeNAwkiEqkg1z1fZOl92a1Tg3vIy8cNOQyM8FM
HMPxF2dmnTLnVsZb86C2/TdUyFOnlL47MzUTVWITS3t9t89xQSOyhZa6euIdDm7ThIaPWoj5VODU
6AA3tzas/k5DjaDlYYbBg5O/i0WKml1CkCekgqy6CrSbqEjDFg6w6c+XxEATOS9bbPKuUyD6dtuw
7RaNTxpYdBhLs2WQwQs0OyzhmQ9535jA2OBa5aNZSNJINtY8zinggjAExJ2otcylFFmn+iGbHHI3
DM1M1SwyZQRlIQIxLp5IiZC4fa8P0THB1JaG5lBmwco40GAO7k+jfCKkmPYv0NMLRIbpQdzujDKB
AZLw7Vg1xirm2qqgIQoIN5kCj9xxYYlwST46PKPntkAkPv8FuheMT/7oxpotyVT9rnB6tsBjkakM
PZJwwSeyaEGHoARimTBpHpPAaqG2PbsV8bbMVkN8bLKTNqXRZeDiUlPJ6Ce80vq3XWgBA89sUt6R
YCuU9wHLS9O95sNxBWAY+s0ipGsiqEA1wXS5k9X8f/uW9q+kRvNUO3/wvMcoCawoAso0GxtWJ9ST
ay8qUaRLAS89WJ7eZ8+RDwSV3v6cLUzYRvD8ljlapJftrrfZ3RaWtLxOnJgBWuTyGBRHVx+wRv2z
pvySmmm3AAEtDOhAYnZoo68EZ/zNVovRv+W2TBE62vHPJ72bj8KNdK4H1V2m9QuDq+qsd0i/scpl
tOa5pM8GJPF6djtmceRsj0iqFC9CvGMriv99tjyby+S2J5rY6cr0HVvq4IbaxSnH7CkGA9FCM/ge
7tjMU2b1NX3l2A9q+yQes4K0WdB3dQgtRdtCKkQba1IrARAYB6UBHH1Y4JJ9wJNPoe5kB9fB7TKR
l3Xe29AF4eXi3msRolkbDKxwGfIr6RlPLYOWANw5Cjfblqm0Bs6VAGgMST1EiVMpXe4WVVx1tptk
ggX7DXDaiqLPCBbS8pBuJQeJCJ5PUo9F4s0p8h4qNTfjXOnOzljbxtMDKOAUyCmfFK09YsnbSQmf
XfUPlZDSCTtfdd+wr1jgnt8woNQR5TouOBgd4TI72d9auJhgC3B+RVz4T2doHvR93UQNHpLKCi1P
xkp5Pz2kmq286MnFWC4V40qgZ4a2gdDb5/J+WW69SeauJ9f/K6srxGJFS/nTEU16uB8bjnzHlw5M
IDkJrc1wc16rYESuqz6r/1mRUxDJdQdhDHfoL+PCP8pRclL3c6wHTttiCc1wEaGXlVtvRRfhlK6K
+zPnPx9A4rS7FQVrefOOgf7kP7nIHp6YpHXUYMYlkQ9YaTDfUCsTwW6GnkpLOHrEXGfnELN5FFD+
iDVycbrm+9Xi/qrj7TjsyKqnFCZRxdu7jrKUq3VQIOUXH+Y/mp9dSyqlLpYHqtBs8n6U3IexLnSy
nzCOSzOSfS7hiDY8nVVTYim3RUGTub4aCWq1Ca6Ida9mtaN/gFXh32dOD2ZrpXojsYKcJv1clZzH
tjy+7sF6rGx/oQm70H/teXIqsw1kikkmn7nyHLR62ex/v6Ka5nhNbKd2B+fjmNV9iMApdSOVxH8Z
13b/SaTRjNJSG3ymdhzgj6xtp+JoRrCvqUTVrfswRASVGbqfCY/BbLRPRUKrmXVgNr41ldFLvVwW
hRh+mVtsb0HdwbF/dHFKb06RlIN4DG01kVZ72/0ROROghwJ91h0uoS/mfE6jqCISMOG5p28DhzRU
okWM47fb42Zy7WT962LB0UAijDuGeY2L7Tl9snAhOVy2za0SxRviDyVvRsB/6hrrj12yXZMl1GOY
AivZg3b0F7nCZomvPk9ofV1rnVlqH0GwCwDq0eYKUm2OvAeN5QKS+CH/q7S4iTEoSGR09XapX5Rn
+NXAtvmKmffin6FLcBFz539Fz+3rEG8oEeMKX1AYqF60tM7eqBTeOy0rxIo6lRd+HG3cnvWh4x2F
jHBbelJhcdGDKKmgWVB+OBE8Lveswhf7+LcAdzed92f9IByXnB8VvJunipuG15ectUjorMqqqKKL
NpP+leJJm5G53gEi2q+D8xdkYbTwPV8EuovAh4dkLz5W8Fc7N/4o3GvGWnQItzSZ4cHbVAstCz4T
CkmmHdcmCsTEAF8GYnrdjVgr5+kZpjq7RbI7zmgQu9C91ZboFjuR/PovUTGmWiTjQvH8Z20jc5oS
xnHBRmZ2SYj8wm/Z8zAAmG2xAvIoxPTL/vXe/YCnf/1PzHFdlUv/dNcKQfV2ghJL8Uo/7/Pya3Og
RS7DLiPTxHbjCsMYAflbbq95CRREVzAE4yXRfppKx0NzIYv7WjYO7dOdaZTehOQL/74aLx43tmfe
MMygQSxXM2RdZT2SHOpBNMyOKD9jPDE9gBfMATYn9YAyoPuvJWUWNGMba+JHkwZDAzhrkVxadvbL
YaMLPo3/6opboSyO8AFwmIkWy7b005dYdOEY/lBtwgt7B6amURPmKDc8d64xfRjwobibAur1HHfD
C86AOL1yuuigwoKqT7tdSOIIF6tssZzxcKSi1Vc1pgNnZGh588ZGKrPZJgTgOdSvo52LAeCijqfK
1a1lCO4hOfIgdTN4ZZca2BBoBHo7OsWU22vmCDN4Qbo1pwYswYaUDIsmVXP581I3WjAEFJyVupZc
GucM9wtMNsai4vBQ/efs2jZe8/U9uUxusTvCsBr+rN8fR+eswT0v+VMqWwtGzbgr0dMmRJ/MVwOb
bl/N4Pu4ZPQY3g6ttDdXB6wv4KvSTclN7RgeNjQG2sJbMmmO5WcNU1ovmtE+PhzS4OxSrEts/gYl
y4kENmMfxJJWHzEdI8jj2JMjg6MWcYGE8ZQNrTXg7BrBHKo+3MusMqbsCqjoG+vy0h9qZaPNudMg
Ps+UVPsRv+CBj2PGp1lAu4dB9Axd/N87PCcY9kKjJHMZKywpnVR7R39TK1oZ4lMwjOJ4HM1LTRXC
PooZ4KcPJQ5IkbYayxufzWETlIvEVhvrIAC8+2rMBB82AqazS/y4Ip9dYSQnHet5Fpa4Oo20Sl1N
J8Bbgz6PnH8fSGSrOVRYbltUWiqtDdZeLNveOA5KzyNRzOFy4JFQkVlwSrdWSIeJOr7wzT2L4KEI
7TYUV1odjpd+Ik91cBWWx7SukxX7DITRIcnP21UKCDHgWbvnCuJen/SFhGazMzf8d/7lEG01PBOI
EJXHQFADFggKqLvdmS8AYyDePG9kWLCWHfJnqknaJS1jP4/AJH3qW2KrP8flDpasXh5Yz95Hi6E5
RpE0XBc4FSWmbu+81l2lNsgNuVe/ZvLV6mGWofmAggQA8tLCP/Ndl2VkPkEqLO1hykc65Q/zvimg
nvMp8QzqZl+uLoHVOoIb1YLcnbBGYk60ey44zW3gFVw1Uvqr4fngWk7x0JNIF8vG76Phn9URTbXd
6+VvrU3w0P8ZIRkdA91ZDq/UVJnzEmN357GlCI8uyqNjTuh/v6z/uZ7uTcmKx1ByL77ByxGJqQJn
ycYtZuTNZwg8muUHWVZv3BqSVAzr4dfmq4rrjaCchx1LJg0tvF8ZTbwCjohXFr47UcT/E3CHaLcG
jo+mB44XGX1Qk0VY35EpambppsWKOzZAvf6KBdOXWnHfN8F40M/zu+DzoEEfhNuuznIKsefBW+j/
1j/wPQ7Cs9A70jwR05usPr0Xj4NfsQRxbwJebyd7ryYcTq9DkOkXFXLjBSV8eud2E9VpHTSARMdW
fa878KV9kDZPgIjMVa7I0C6zqeYDKIkmw3taN7VRpiyS3Akqo8AIRXCcClhFiCB+fAYtkVo/bUyr
JP4dofrh4T+P1HcEou/Kq79zxmpiQN+9oZq82XGMoulAqI1WWu5kZI70jbrRPuTqhO0OKV4m2tk9
ynoAXtzS+u9aT0AxXxCDMFydPPqeSnO4n0ntwCatOy7RvNU5ZcbeHZmYhjOlB6hjO95eIh/v+RkK
rb4OFkaJ9a6uHPJb0tus76hSIrtwQvh3MLadctjI9cX6aMNWOxLKubSBaXIoESwPEOKm+UyXBGYt
XsfrgkSHG2yhrjyPxIxC/t14QwanCNCgNmRsU1ef78wk4LIVvMJCxqlpjQuUsV0jlISgfsEEzzdj
/pQOkaQEXft8QJAXgexA6NKGws8i8dtt6tbe2qgkhPxQf/riQBly8E76MoOaCDaC8yd7r6msviJ4
qGfBdxL3PddVrr261g/jlBlz05R6dPARRyLdnKmFU+mreke3GRys7ROknsnvNsgfnT98aP+bdaWM
Md176qIbdpj2Xp5SnDnHPszC6WFehfYYoLKkZUrZMoW6VI7JWsi3a5EIS1HZ07ymm9wVwV3cVKfh
ETlg2Blh/0B6qRlrzFOJMDZqVYQx8kNXibEpGQfQsDKbeczSDVOoD6JkAf666BZ8a9EHW42cbSCj
EQlvqkxCB3D2FpyaSnZQ0zU0CctboJGher5bLI2muF9l+t8Mgz7q/034I1zgWyuEgXw808pL07mk
IGXp8P+z669Irof/d2256ZIOHYnT7PtcHzEtnfwBwbWDKuCzEl9fDB4Txu4rzZTbmi9dwnDhues1
0EIxVGX5llrIBD2CoYwtUBpPD2N9JQKYpTTkzCEWNr4wmGr0aqEgWVbgrDilNX6a+rwDSZYFrrdx
o+NL6SwM5ofi2XVzQ4lEOLvZxAlLeMlkDEO4b2jYmCSDfNkiWHP1qgNL329XlurSt2jiTge1XHem
IHrT47C/7LjMcVjV+lbeOx66dakqrDb3RQ4wRuZAkJyIrknrc9uxcemtNynIWW+6j8VaB+03WLbe
oVAAOemnE5IwA7Kw1++nAbvfhriljeTHcRz4gS8GnpuqT1do+aIsIzVF3OOzkBQXxcuwHM1SJuwF
NhK4Ioj7Xcql6HctnZkRw537jf/lxvb+xz2IYSEyBd9KaO7/J7KRnDfDrpb8LW2VpbpAUJOCLmjk
8QGtLt7TITJF4PZMwzxr8GdxNfXhFr0ggCFd7Rm8aQjzfe7+xLIoJdmzkAt1Wc1xT8nGkx7zwz2a
S/urPrMcwvYTy4/4vqyC2+TbjpAB88+gw/WO54oPh0tNngDbBrr7XS3QlFrVXLOiADi0OXdVvs2M
VkQzdswH2mtL9RQ4eVTzKcgXJeoU1JNreXUtoCAYcNiAxY8pSPS8Ds8DRuNs6Avdlne8kJHjD453
JOB1tWpsEaVNyawQjiXzDPisJaLE+/7Z1aYwHSl1kMqvajARVRzXBBR1TT6w0oxsytyKL2x4czZN
fOAmKPm4iSAZyZOOMlJkIcp5DyTlW1HyNlXrllh5mm2UQcmIlS9f3qZZ/gplqmjo0oLfvx6O/dL0
5KdzMe96q76/37nHy41G9tY4ihffgdZudlKDIElqIfs1ERNmL2P+MHdgP7dKWnOsoLOVfg8FRa+x
ECujcyufrq/5lPdZVpmCgq9O24Eti0xRx5qOwDYEEDq7PdNDKDo7IE2JhnXQfqv4SPfFsg3HglWw
hjeyQlr7+M7wxZx6ZA8Fvyy3SygoqXQ/s6W+sBcRyDnXzVJ6jZ8cGtslZ+ofgCIrZwPGmJPkOiW9
KFFKnff6avzWyD7W6JomXvyHzNkm0FNByME0bqq3HdHYG8uNSnz8bwPzzg7rTrsKpuGQ7Zq4dK/A
CpVnyCejDlb/xNqF3/TFFt919Wfc9juesDCYk3qqziMapMLZUOIjhV337b60GevLBSRFCVd1sQCb
O8HTwMPP3AUxmqDsC5El7q7RHEt/u+STk+fddzgoAIV9I8rnk9G8Hu70uTxPC3sZgFduyqYg0EgR
jXiDhobnRmEfJEpOMvvVFrHbdyeSjuc2P818khbG7sP3WM/wMHCE4oIVjz1soEugOAqhlqzDdC+W
RND8xrrZ6A+8SHk0XHMFO+YD3bb8gUdNfray7XFtUwJXQxIhARrv8xFlUbs0OYrzRr7ASi9GCTVq
7P5hpYBq4xjE5HhH90Nu7hnIRrEvXX6VFSHrgyXN5GnxdOr1Zzwn/KxYo+I1EncGDoj3mVe05Abm
+Dkj9a7FgzpeypMBi4os8pMLXh9NDjn2Dr6kukJsvtcfIZk+gLvXSkjpZ4Hkxzck1jJ0mfJ2s3gn
Npy2OKTpGcg1Dyy734ujSiA25d1Sw+nGh4YbYhYoQTphtgB65R0sB3V07WdLOqA+Qn/VHu8heY9j
ifCcrBTcTMOZIowIZH0SF0JTZV118uYkRbAZE0mSRjgNNaLrjRNsmzC3BHLdGAHgAKBeoVGKLwPH
gMoKbAzEyYLX/371LfDW5KqpOvnCJ8ng4/I8+UaLGEziHyTOIeYlwDTViQhi4ZRxvAG6tYZYhpdW
cta1mf4zV5EDvFctiRFkjiF6U/FJykXrUtzeqzrSqZpqEUyV+LXG6PCVsN/JKcwN6eniyNwUQN2X
7ZqElO0VuX6j+z9obVHIaM90JLM0YwHkXAuyljW5FaQjaySGkIa9uQs/70iaNpxvaWj/xfLdnS6b
qNhvQl2jf2oetToRlaEnmBjId5870RMSthDFAkg4jkTpnWw23aPyWieQUTXmwyNIB4V8lEl92XuC
aU/Ngu3iBq6kkLitGKH2NrE6no29uwwN6+9gsqLOKsQwJH6QHgXQh932vynSu/iuzMkyKRFQkXP6
nF82qonASruMJJoz7dvM8RXmGvLUPFkKkhSnKhoO+ivegDZxpFsaWA1QMFus+VX8giXXFlCjrz/q
03lsu9gs4jT9/77pvvvhLEZrBfhyP2GfXpYJ/WqmwZyqyChr0LP4+zh29AUqJEFIYMWRXGeNLwTz
i6JLXS/jbFTZ5CSfIUV/gstae/J52KNrku8LjahjN8F9gAteJB0RWiQMq91eKVzQ2yGxXbbj3kvF
Jh3QnP6x8WU7LDWBgNpPmUPcY1K2F6SBOf3Lefv8/9ZtZcxypa30gU8Nfa2NS8Ik/Nvutwtj9LhY
U1xTQ51cCPZ8kb2U1uru7FiOzbpSzNG8PaVy5ZTTlYdb2/kJIWJOA/lqgnKMNAWxDKoGLks5ON3Q
g30mbe/YF9lxo86HD6z50u7SLC679lEmuFwkfimNY6BPp0a6pfuZnp5FwviG14+mtCNasc8uGCiq
hVstlO7orXT5/t7jX5laVd99G0opMyVQq/e55trqM5ZoGvVchyBbACxReOOeSfZt6Po4x8tgz3Zo
zUkRE0cz3gJQB383I1puKGA2L10vW7MmZr2UT5mL7aIu6fAoLs8hPglklWQtCF0rjVs7rGuE9K2Y
FfIZG06HEpS4WrdeKjIStnhgO2SJjEf6e98z0LObj3Mfsnjft1AK5F6vleWgMQsoCiyvoBdf7hwa
1qd5deBHms/wCAUH2C1Tz8l70x8hGfvhof4a0CwDeL+2XW9KK9eny90OnpJxWrX8pO3Eo2ZBrWCn
DP8QO6XYJYRqE0+Bs4n5t8btZOTsaf0vaK8t1w4a47FPmriWz6cLnm9ISSZNtKYaPULqIthVy3bJ
5NlZfk0dcsFzzxc1BlgIojSk+V1Az+5UW3+u4fGQOZnBZg1wL5e3XYF13sDyNrf1uOTVvaU6FisA
IILSpNzm4QfWrLdevmO7GNfjmdYkrn9TZ9Iq6lyiUl7/ih0kZsyPJAUnouYvG+4dsYj/XZUFAb3J
OvtS90yvXPeGIYUIpKNrlgbj/dNv28STSp29+ouzB6JWa9UvgDjYTj3//jByzQft5ALNTFWCgAZ7
ykBzPexMoIEVZ9ZTW30Q3ikHFYEV82FqLNyvu365mQ0oYQw8wwxVVq3VTL079TkDw0TVBF5WF+LL
SBWP9EpMc5k5LUs5Wu3gbUqf3DcCngiEdAz8r4U5adrZPSBsLKDHGtJCQKUV/x1JHB7ZsAHQh+TD
DonqLOIY/Pbd17ew4uOlDk0ZT2FKBjHjoxMb37w9bpGl2LgDhA/hDDzRDiQoKpJQXvyYGuFRQNUW
syXfOZPH+swmROOK9Wj0ZO2YztdY7PQuiTMJo9bbxj9JqZSn8pGbeFNCWYEc0cOMhEpcsy6r8ni4
IUUoyg+fjZ3576CeO449aE4LgOrv3MVfzgDKXlGT4Lvas1CfqEKD9xh8/ihL/8bw1nW3vlJijj+G
G1roO9gjsGrlCenzrKM7eiwJZNZZ8xofHLj8e5ORM+TL6rbR4VhKO4Z6gJqjbOijfNlKF1PTIrqq
gmamp9f5XcopvGNUBNQNNfoPACYujgAJniBN/rX1qHdBXHmbNYzqVx1ppS+pn26GuJLrHMLs1put
8SoDDjqtAE7lqV1FCXM8PpEyDB1sQ76y7ZQL+KJ4goc69okN5Uz6v7LX5wmQct+UABBXKJNuEHkm
Lypxu+GICxeTbqWEomJT776DrgxLtxmHJ/id5EZl8YtfvLFn5qIxzRuNmOwhrZEAl3sMhU/62EAD
x3iDpsv6+Il3HobLnGvN+S//cuqF11ygOxAwd6Nq3Fo4nUuzYiF4jvg3JNJHT7DQD/OSzElEpnFI
I/RzYZ+GAGM79Z7GfonITrVDOu2wdN8ig/2SXojUQ+vcyvYywgtEOBGnSKO8702e4nfkMC9Z8KBe
GrblyLLvDlTFDm+KoZDiehTYR6rg+zNjUaqXf6SegDzQskThitAEy0LpkOH1m0CrLNXfC+45K61y
b6H49ygokxrK016qICl/SmZKf74p6jKM+WjN2fUTBqKvCzX9zDnMkcxkA5iWmkXphbkdkJXCTNHP
A5dmoesKn6Tp63LlxxNm4Bz0HoEt5WVut/AuDXW6Ldb0w5Pzv448w2LqW/ldBuAwc56tDBNKct2J
9n0aCoUe5Cryk9n5nWteovIHwnt7kG8c/usU4oU4tGfFVLdEPN3pag/gpwc0obSPEP9OaozMbojI
FHtc2KipbFEajQMWKx3HhPM0j6NFLrWVfTcYD7MIRV7XQ8JUFLobGrJy/+cknBJMO1TyJo76RDpS
G6iBqbICeX0dCUN9NBNXnhBA79eFKYYjSg9HKfiYNFEwPkXnkX8wIR1aOyYaM8mJWk+yN2QQi5e+
O5I6Gs2KDpVv83oWGwkf4vlXNapt05DRK6Hcc/0vV+gLu1yndi3nZGwTX65GO4MmauCHaKr0u8B0
i8tME9vRaNc9giJysaZIC6vgV+ouoKIIYRLsd1HXPaq2PWMob6wrtDxUYQqv7SVUpRIdCHzt7pkC
V7qyPxr+OApb9kmoGD8vgc0jST5LRPBK7Q3zyOKL+LQhmp9wJy8PpG9DKPWIBwioWtLsG0Dr+84G
zvyLTabgquCPvM2PhEyOYp4/6LlL1f2gkR+7NK6nIh9p67FUvO4ybt2k0hau3PkX1qhDHwHrfduG
UOOGFEqfOPFt7zJMx3bAmEpEjDKEKT0lBDvxg82gI5+wIdBdiEd3SraDPKASPutus3gCE4/a4keJ
PE0fNwLr/62Vtzfrs2XxKVNgvUT38MEPsA6PR1GOUw30sDpRjb0ZRRTe956WbdnCkS0Djwr/SfPT
s4C/yd3u8k3h9u+Pt4dIQOsA4kL5W+S4pGYhjKG7RbmvZ2XH+K35Q4uwz1wMIhmjc8HarDA2cJ2R
jD3Nvibk7Ry++KyXzVe213I1+nEp3KEcrObydnm2bjvKHU+ftwZrwoZ7z9x094MwxM/pMY4+rkdG
shyiZYlVux/Mtsng/oHb/zQ2+HKeqKL5PUxLx9WsfPdL/Z0BjFsLWeXeWiDMLQQmPpHVl3BBF9LJ
A/dnnEz1/CIQvbDLIrKNmqljFC0M+Lju5EtbMyAd5cyW4NKUGy6rtxvjKFhYPvrDNx/xVfjREfuX
Mfr21wUoUIpng5JQ5y8FcUxnTmNZVeu8zxvPEn82TxB/vKiFN4IHg5Chu/XtmEsjE0QLtC+JVW8C
CMnq4ZLmq9uhNTIcASGw2fOsQcWYnBAzFqBJ2FZKogNmPSTrRD+1JmtooouzfDcjmz+oDgFBnBHd
zut5MSCqEIFdKEL/nQxZNco9nEwMFjco9Aiz0rv98pXMDIPLsfIF+b4LpdDKYJ9yjwIZt1FwlTGY
hEsvy2mn+0Urgg2hXy13fxAbhHw2305/OHVFXsObluyybu6DSlIXYBIqVr3c+me/wd18jg2euqBI
FrEq0UHdws0ILuTw129gJlfaXMflSJDJG5108MgS+75PnnPigKy3jfaCZXXXSLUCgU82HGy8viz+
B2IOglIeTy49yOSR7/EQanaQU9xtSbVsIk5Fs3oVs/JuZNII+W2TZYfAXH+mliPNVl/XJg0DQq2s
tRTZ5+ysvib1aCq1bFGfxQJc1e3LgokqCUllPz0UhZZ70JIeC64KGx8AGbGeBHdgHyuJKaInNRjw
UYAZHUuKRXjfJRDTHhBrT+912DFbLU3sh8n4XC2svjKOuRZP/4O6OWq/irJsxOh8SAh3E0lDnoKV
51wi+sBhdNJMN9xNfsN9OtuZAUo6NJG3Zn4VgxuSXDxjGj+D4kuS9uYbJxHc6IJD+ztWo6YEhhmz
xOYb3a8shrREgpYzlr8XxdUUlgFAGsIFeNGCi/PZA5TO4NtsC1/EnVSH4yKu71RGoWA/3eYKbSbI
4q8x+2VeuCHzyTlgg9dXjSqTtJUYBtFK7T3/Z4JgjOvsgcYDQ344NRC1JovwgPPI3OrVz0y2MnAi
v8+8PT1n/CF6q1ypCSG48reSELV98QPiriqABSeMTeTHspo2LDrtufJaW/qyrZNKm9KoO7+Ff0mS
/BseKkXqfLXlHYNFbfgevXnJXPmGuC2R9X/RIc/kFxio6Hb9Rp7wi2XmxfK4YgN5erC/b6YVBIIB
A2le4IERkUbDXCA6Er2ReU4a6MZ9mTA/buKtChHGhNRz7zEI3fwcgepaynmApZ+cmlibNnwL2AWj
Snb81Z18+jFEdT48zRhqB9GdG0HZ1N6F49hRoE3L1tVBFrQXN1Nyl4p5P+YQ6Ecnvafhri2DhIdv
mdpYuKD0FC9NQigiOmYZIHUmbRXcHO4BfVOzV8QgLvKE5OT0XsqzEGrN6bz0FvDZDxCbAl70yxVq
6vw6kSt+s8sz4lyXFEafTj5zek9LLlf9wfhyCTUfrUg9IL9ZFc3wNeUlpYx0rNJFRQDOXMV4nrZi
pFcav/v/47+wXobyTCQWavGKxIPTVhk86Jam/ugTb7RUM4fnlmNHO094BQKEg2Di9eD4XjT7BI4y
MiRDMYOegkkKRD73UlJ5UOBDlsQw58Gm90cpRJREsuXw41zPDCvDJX2QNeEpxBpu+hNpud9GpO40
DLKCRMxWwExiJ4cKfM6TpFdWLP9Q4amnyCCtHoL60OvcK1/zGaEOzyNF+Ek0vmtwgVZSLXbgEuHP
a5zbjMSW9u87+Wez4KZh2o/E5asr7G3b49UNQ83pDdWIMwrtRgv/3i4u7QMlb2hmj2JqW2wpNYux
hPuT0o20ZpOAQGcR8E7ZVvXWIjzsYLG1w0Z6sOX4UcYWdkjq5wdRV7Nsimt2o3bOckLkLLRh8J1s
P9avOr5ORNYf7l/UWbO2FAs8EaX2htA1/E+1lLBhvM2R2t8fZvfPx61zd9EApjHz52sFc4L1iDVo
yJxgkU/eWqripXd4e1TMKjT5YaWtp+RMCzheMeJM+X1adgW2r57fALC58MRc2obgTTOKghUW2W/K
TBlNBfH20G5gRniYWWoMp3cOZ7Y8q73HDmTSVF4QgMnmNWQzVFeNPel5rCjjoOwgUxxaC+EYVk6g
7aqZ1qNfyTPUr2xPERwZs4ej8cJwPM5oCXsic0wgtIkxo2pg+p8XE5Iz/iUsluWmBZ4/xBELcltG
9NYmbQ+m0PO5DoBZvd7wY1S4NVa7vMmbYmbBLdbU0qs64a5Vl3pLUPCwYeyTjCo+l/3P9vTCLMEs
RqfSINOIxQas9wc4Tr7LyYRWZvzyyjDYGdPMGopLlDuVwd4preVFQmYcBF7xzE+t+qAXe9k8Jsin
ej0xpWQ7PrY+9CaDKOjc7AQfIOa6R9Lfz9S+ftf1u67VU/N2Ql8WWKk1+zatRZF8J4R1LzJ2hbYz
g11FGEQfZzfLkleMfholkMfztT5z/LhrnrBdPxh6+KlnSy/wN1UR3iuU9f2bPnXG3K1HsAxCtufx
l8fKI9VXqkIJXMPm8TU6+gw62Q1Kysmiff1vqATSkfYnHHURrP6orhBSp2JS8/Z50shLHkrzxX/S
VVxxP2Jz4QGKyYnnQ3RlpYizXuPZb/VgS3fX6g7+iKXOqa7N5aIl+o6JVf0p20yEccHzcyf99rT/
6mkgkmduTYfRgOk6uJ4KchuLEBnOuoESwOztjC88PjbYzUS7WU9/3DK9601xOpKEZJFxT/EgI1g0
dZ3mKBO1yDfP3RSr45OR3cB0IW/lbn88KgqwJ+J6+2shtv8lX40KdU37MO5sLSy4sqbJ2zt4Btaq
0T+98WyRlBXDKQPv3IMU81u02JgUIbfGiijTYuaZ0NrCgkgR20gXZCXIHxLjVvd+toPomN6U5kHh
pzYwwABpNqKwx/csXZBS+wHiMU1XxgurCYrBz7PVv9x4+o7JPgLdo4QSiTIceQYQo5hVXxvMR7z2
PgUjdLCAMHb1meVc5veqKYuO4KErDq/5vdjAgb8xLyZN/LU4jN7tbLLgtX5LRb743ZxwAwb7tAXt
+awE7crnzjEQgClbIQ53UNDlUKGAGhIPnMkSTBHz7jHolvjYDieNx3LTO8U3zF8JebRiakcXUG8o
PtLIYrfq5rfsJhIGyH8c9kDniYqhLtyMDdH/OFuFxn8BjZG8PrE+9Tuk8iIt/87Hsi4ObrMhaZAj
1bhTanOHku59Tx8YCThUmMKFQzqA41EBuYu9/ADpzbUpgzE3gUJKQnbW3qzb7rEgKArt1M2McNhi
86RIRu+4xA5NL5tRDkoOZcVd52b2Ej3zn+bR+1wF7GMNdyu8f/ULGSjuYHyLExvvKk/VgH8ywslr
iT75dgg6KCDP04AYmrBheW+rT539lsFezjmPCW66GjdcmsRelp5fQqMkxONrlJPm4wq+Z/hkqjTm
K/0HlijQinLnPzASTw4re9+Ii6qcniqg4uM7ruLsZPVLLXlku1Y44McbdYtRUxRGioC5DdSyayWx
VoDtmIKjNJpv1cld/GFeg4ZNbWgsXz5QvZhYw42+WJE/XEHEv93vonShAuOL76/poSsxqFV+w+v+
THHYzSs/lK5xXJwpXZfQ7eW5NxIIfddCrFVIRBvYAyHaQv+kqK+SnQVx26mPN7qB/5lA0seECDWp
ov+57NwZtYHZOV0kjc40pnrnSO2U9dLUKgnoJ4ZQr9ylwLOrxvLS/yphgjS5f1lFzTNk3sR7OZVa
Iqeot/+QAYnuWkKEq76TDtbtdEyjDVnWiT1mHcFizTBOGgaUg5dmTDvdiiZ7hdCYtdtFeEdCOGHW
SffRcP4XEzhKhIpWtNXtkdcVH/uhfkV3xG9LNQq9dQ7vDpIwpv7hKOcjr8B1Nk63BEn322lyb9Ks
k5Ul6Z6d2JByXwScjKm3ffNokGqKovcieVsEkJczokw87abzSVHuZIv0ghZCtl5nAatU5xWUbgll
x1YmcwBt78PW3W7CYMe5OqRlAzdV0xFwKUXEYgHVIGT3k/NWUsBl9mUucXWut1ibVwytktSGSZ/W
KNpMHhkj+tbIWaPErC+3kvyoPUv5pmmiqqK4oRDpw0mvtqupzZkV6Tbv91eCw5XPpxyutjmou+uO
aPh+4dKjnxYCrg/yLB2pKJKgyiAdOaTtG0hZd0ve+7QZyfuV083JPJG64W4SOst8fZyWXn89eh7R
utyP04uozvhYUALQKPGtXhzGZjGKxHjTujkL0zBJULvwe+na6VhUOG0iPYr48t+DlkAT13rga5T5
jJy7CZvPyfPfzOBWsU4tE0w4PMSD6VAsuAPzhICew2ME2uwp9j2kcv+mgsKflUWOziv5zZBxOGXD
LkF8So7tSzdtyW9Y8gnq+FZUqkC+gPM+Qai9bOsK9oYcYiu1g5b2NcXmYgwmCtBuY9TA1dZAJlpe
s6CaTveGFm2rW/qV2rd7JW794u9HToc5ExnFmZIyNePwt8fwu9BNlIzCtQQLNi7EKCyHaP4c4Pm2
e8kZbxfN27epW/GnT5cQZk5Wys/ZX15IaopjImqpw7MJxF2tfGd3HcPVZsi3kzVHahLXL/FsJ7eP
LYfQsSQGXaize6QWb+V/757jzB4D8OBS4Yg9Np6UW2eAbsY9xx8xKZ0302sV87+ITO2v5Fjf1TC5
lByN54So1EzlUW146uJqnN5/AJiATAIPZVqcfW+ZYlp/FCD+9M0UL587u8aklD6d0DQRYhkqsPus
ENIrFB/AvZAYHbjWJwk2djVo8jmazaEP9bPUudHFctwLHA/CUa12BwEFDuHZzwxS1DlhiZPcsHau
pOB0BkUVwnN3wvpEUglkzgMB3VhDuTsmM4a+X4+wCVswPbvDaWQUw1FjEznOy8kxvEd5lRoGaLlQ
arey7+NWq2e0GVlmwcLu/gU899Xkgyc0TTGllEEbv/Spenl4wt8OJhlMqME+qgJ+N6iETVwNT0N5
+dYZzvXUT+c0rAFaV9T5TyqQ9WNZ5fd1rQl8e9H4mutDByXw3gcWvBhZmAc6AUGEdfNeitwXtEeL
WbwTD3iKKt2l3r4Od3CUl+HpNJreWFECvXD/fo2pe6wpeE0SoK5gfPf63gk3SIPiSC7XdW13fa7W
E7DR77vdOO6Gd+E0A5xQOG/RU6a+BXkHuGHRSsaI18FP6jxhcQFk9k8btVyy4PxHxLIpzq3ZPUk6
sO7VPAcPM+ThdBapq6/N7Fdrqci1v6nLlORAzDBYpANkdtta/rEjqTc99aQbC5PpDPQUCX3FlaSt
qDlPzR+y/mJgzzf/yKBKaEmaH7QfvXbIz/LgY2yROadWAI6KSumyDcAXtszgkTsYQlXrPW53377E
VAvM9Nh+qkQuSQfwwDI/b+/nLrcbZwaoE4qJMHjC2CXk8USHBP402JmAX+8xU3Tho/TmebAAnJUe
HatPbmaHV0Dqgb4D8VJBRRr0QvObwsEiM3UmC0v8h88kzieTgM18C4/PQEQfH+S1fwhZGn4TLNyQ
WVYNzHQyZ3Uc9bCjb+nvL/uKmhNGZYP8eJz0VjreWCMguqyfRHffU7DYEIc/TEcKTbUqjo2ySYQV
CPhRrMbpVtclzQ07FUvRGqgPJl1ziBd4Tfe5G2B+jbHYsSz5cJxa6K1hlKepPwK9rknsnMbPJ0iA
XfVB8qHMhkGZAHJXK78HjnwKoAd2MRqwRqgDmtD8rD7BGlCzwa+bkrU6U5a/UM7K1fqoSbplzEYQ
QU/DGSjAYfmoDZrVsyJXKVf7JYwzsgl1RZflxxlKhbacNlvUkAKPbG2oLcFyfJQnhRCpg9pG3VoD
gSW0INJ5jJw0UAUpA332uyNBDXwY5iVRNFgTaSk42tDI6gB1b/ez5xwJQoc20AeYBWlgWClnvt9S
d1xUxacjclwJBKD5Z415KDYrVLh2qRY1+NwwAvifbTVMT9QHgeL2QpwxHIZ3RtTscQpRr/GFfasN
+mEsYFPZYD7l5LTcmlPLXo2AnXfJL+/nV92DC+inThRRR+lhIelUS+wG0ixXfEStx0DBNo0rpO74
Xhp6+Q10EoPW9XrueLzkUITMHS4MRGo8LvfMeorip0C6L6VUWsNcyotIzmrVyg9YPa986YZuCW52
r7Bc64FU30JUvAYscxWD0tdRz1a5gZq5OqXJWV1CnQkOvsH37pfL9ffmO/c4PtAx6FzSnj6jnt2Q
4vNM2fXgian82B+0BGroar8IY/3/C016kxIO0FZVcUcCrsPiaqbm0+dbjPJoscWG17M90plLWg3R
ZJuoWeykeGx+xWeEj4sWVv6A5njdwbWqgwRGcSDrQs2IkmEQUlz21Yl6ii5IYQbUHBp99btz5EjQ
F+BXaUhhFqiggYQni+Nan24g3XEPEd1BR5lmxOdoidCbTgbXr/dzcaFofUWp5CED76oilvHd4IoW
wD6Vn09SY8FwmP05jBHB1SHLByNuEv3K0a0T21eYzLt02b3TI8VkR11EmvIDxPURARXBKQHNgN29
PS3hq1vUWBUkQFiM46OCHkFtzKkkEjys8JZ6W2E7DGCUDiaxED02Hi7RVxIFrWkSGJGW0AgNFeIC
pNzJ4OeMAG8/PpTNLt7szAHsSFBOrmBfpaUz8RVMxgDtLl985f/shbZgPeKYxgDBwG5gnMuMwDnT
eXzoCc7DCrYiIsKxPeZA6OGGkW73sjI8r1rYTDdr59ZXraHQBZm8KLBja4v+ynPQ5Uy8Hk5LtzJv
sSBvyzZFdtYzEjSC40cP1pc8FbF1swSLmLpikbFNM7q8vYS60o6EOjF2XdLTU3AH4kAqASYauwQ4
itjVVnKoP/BV/OeHaZcecud0evUl6a0Z+yRKyv/0AEvvea3y1yx1SLaY1nLoAfkEpsCo9a7uuwiu
1Pm2kNQvJVKfjR0zrtlbqOMME51egwaaP1iA03h7wBtVOGxy5XIa+7P21Dhuh2NvNtYwNCvRy9xN
HsYq6lOS7Mo6KDYqmZG1SDzsiKdeTMH7PSbNPDseDtpgbSEGXNmh1lHbjTdIDqF/8tKecsT1wKPt
lyvXpTj5W/wSoPK2ARxC/qB7cbJJDQ1j+hZC1EHb3x+0t7A4axFBzR8S4lG3Fn5lIgYXzT1fucYu
c/aUpfdUg6L6XO1MBInoB2JsEEjZJDrlErFjztrABfaSi3r6OJSyJMLmUYmLvR+hQLal3/Ytr2MQ
HgSZ9fjK526uyfniX70C+4h8obMI2kne9FTbLcyVqatO633VDHbcRdbi/F9FUYLg5hqqDzhHrRri
WUSd6u25LCDa77g4vcyYR+hXoOzxv7q/t95HrHL3OP9HVQlEVgjwiuFR2NL/YShp35+NE8tHjhm+
X3UxZRule+Xrffl9/oYXVF7PD061KAxFIzPhDS6AmYZaLq+vQogknN15JWlGSs12nMdy+LYRTmn4
Sq6rml8yVxlT8UVkJqEtUm6XVaekwl/cjHu7gPemzgIlvt2ClzdvwqwYH17TVAMpxhN3DASfdc9O
mIasOsBfK/8gtuwafPzflWb2aLAusc30KZNiGb3Z1urJ0WMahpJVpi7v+hDMxe3MlEl75EsDf8Fd
U30WgK49EgJeiRN+sXuB0JR1JJ9VzFeAbsoZPQ9KW2nfeMMVmPZHk1jJ31KYzL//+K2kOXR1sSIg
NifkMgt36lncciMfyvb8W1MLsSqS8xPJP4zSpUxsh3mzoDFQwf0vsByWdoRkvxdHABLfjSo02xTx
O/eN5uYEdUjUC4Ajwg+d5OrVjp3k8djEMg9dRT2fJWZb6lkcYHFBXtV85ZZnBN1iYvSXQx/7f6a9
UcCAWqdjGq4WyABy1ffSKyrNPWbONYpvWQh8efGNYkE6gd2Wqpe8lWy5CjBj1Yr5C76KYt0L0rKf
g88xViBvhG7Ba5IPJ4BZiwW/V9WGVZBQt0w9wqL5pIqjjwPElPRfWS+AxfdKW8LIr0bwQ3kQSd7d
NlSuVXQOuVR6KKH5qQoV7JkRTLxqpVERfJ9d3HluxE0UHmX+QA6w/Pv+d74ScLT/S1OIJhnJ+ACk
rku2pdAekTeUTEZNFRubwzPg5KsmwXCXC43HNK6U0Ih+r6uLkQZ0RVdmnv0wC/QkiRLqsjVPXYMo
4fZiWLyY7pcCHt0p+tGjjcK4mWBHxNu9ID8oO/rdxUS0l2kcoRgFtXy9fhXer8BesISgS8OLtmhq
vD7P0pSKg8m0dAEz8sukzRi2VEd5ykad6+q1ZRFzN+P8yYXG/CidrPUlIT2oHyfD5FXW0mBUsYpY
5PC8Qr0C4a6eXZULgfX3T5wB/vihZTz8yL+tX5llthR09ZiHOGoh0gObnQQexsvJn4SMk/SV2VRZ
ihepsHnke2+Ecwt5l6DcbaYcWtM6RBBEYZr3v43Jye6ketxmW1qsHasWjUFmA6d9CiUGqDGgVz+W
KD3NNRD6085YXPa9s15Hnous2oDX1WfOVb8i4cXDPs8ub9YBPj0f+1dh7ykOdjmw8Do5RU5GR6lz
UgIwbiVwvlI7xYg+ZlVdEhgOxw7VrKfEscjwjJHO7H4gyKtor0wn6PBd5pD7zJxJLLamHtLSCOxg
9Klbaj3nFe1FVw2wFxIdDML+Jm1mLd99NYVvo+dTBwnTuAtET3prG3Sm9j5NZA8x7WOBeyPGC5e4
q2vKnOJxgmSx1rCKz/JOv2sNFOPamlJS3bZya+B/M/adOBMvEnJ91zYISWviMwojGO7WDqUJecD/
KgCZQqQzvV208KTLxbbygONMgyel77UyDPhO0Gfeumd0JAUiO0apTirdQ+WFi/1OeS130Tp1brs5
TARyVJzKfSHf4M3iMwxx4nMWf0EWnjjBzBXnnb+EqrPH+7OWecyQ8h9Rp1lyQCdfQWrLu7ww9q8I
b9ZJ2zLaaSpc17av+z5/q1Cytuh2th3NoF5FvQrvHsiVB2GCez7WGdGarUDHIMgmdr/Q47fbnDOD
+94N5JF5TghqXHZQOODZ5CECPcjWX1pzGmFlyumKPv5lT67WvMjc2etnfgRZ9lQOpp3F4WtVAoB/
L6n2eVeEkzFNl33c1F0puGBuB6Vx+jYAWU9skBOLYhHyfzGeq63yzlHE3LYsJHtaVP4SHJBbOFk9
Va0BaJZHwGT8FTuiduL0AEIrRj8f2nMzoM6z2T4jwoI4s4C0X43SvivDfcW0Or6mboX0vvBvr6Kj
Lvm/X5N5aq0J/3vv+n4Fmr1Z/SjZHWzpjjmfUHtvudwZDyEq4d6N45TAZ/0K/iOFUlhSnOVJrMdg
HQ/Mf9LwMrzsnapc/Z8e9fB23F7k2+Ns31ekKL0LUYds/PNov9umDkr67kIdgy3fY3/iqJUqfeT7
xVLE1tnqi8OrNDsZkLdHUuKIvmNxlev4NCMMYJkfaRD8TtVdTDBWAWeFAnGg6yyCqHnC/cDwPj5v
KbDCIFMrpNQTAG8S40ve8cnu+eRU7cbmRUbRS14qPKMV7PiyyfdmnTm88EkH54+5fo0NK6ZgSeK/
3crCWNGHks22vSnMrD4HHsHjZdJ2x1Bx6NxWAlIS4DINwwjusmv92nr2rOn4QJKJc82ikeASFaHP
qET3Ujc1PqXT2O31Pd6s1lt+2lasFNBG3GhEPjEc7nXzOK39s4DTvC3WNoaGq184doVob5n31DJ1
x2qNxvTv4jY61lxjKE/gHb137U+ZcO61GGGjAgfeVbfUtEZufAA5WD4DUQ4BoeMX93lXH7IBokrB
j31NV0+ZGgN7hODFm7wmWKIOHzs2MLycsn7uG3qM//FQVKTSen7GZ4VqxFMVwOlZgiY5Hwmc2P3K
yCSUB/AIPfWdIW/kHyrwvuGQzsXXoE7Xh0AemOXx25lo8D8wxzSPM2oP7XF4oyIfX631nc0gPwcV
tovJ/AA4u7EwNYnStYJ4TAtv7r6VsUlGRSnBA9UNC7517IqRmcnosFhXSOFY+KtrYP9R3zDonb7w
Sk1UzKeha8xEU+QvQiPXyJxJl63bw/hnb429McAoV3mvrcdYVJX8gisAAfJtlnkCGx0SorxvIoXF
5SLBgH6MxrZqnF6O3Q5OYtaPeULA8ghgwkzqI4wZvIWJd9pBufo2aXh0RgCunpA1cBlgUOTsnb+f
suyfkJ7zzgpGo/ukEn3qB/BA6tmWwlFaL97zChvmD0QzemOQZYjrzdIGlAEbhyw/Ixhbh4Vq2Kaj
Eca0zFYX/4JdyPvZXWjNBWN/1fWo8xQrGTRxLzx/9oh6gD3qbWXGyxZ9AjZDme6rmFLWRgaJjcet
t3z79C6utUQdsbEQkWVYBpAFSunF0hBCMChoyh7Eg9Th0RDauIFt+px/69kHa3X3Bk8g3ywb6QD+
PpxCsRQbUIYQnn3SjWYWLt2BIOU/2DwZLnKivSBBuK9Pna51rmyIJYylJNbr83iYnhWe1F85IsCq
tDsWey205l//v7pVGNePAVx0f0EfrfbRmpmDMO7wPJWcRfxBhNYIsA+U23qs2eveKJHjfOkN9jra
ydv/pcuk221Z7rigqbH96xPmmPWjujK/ysOG9prUKmmCiEX67UR+WlM5a82XKvfZI5B+X6uqB0/L
NJti20p4oaDsvAp6nqEjp7T5RDrOu2YpbbaSHljXQNntcX8WWj4ZpMuroa4HxXAJz+vaHJD1eUZB
N1odJP+SAbXM+ERU/H7XJ6k4Al5UfFcihipywNLOkrDaG49ER2Wn8U4dBkRsBm9DEPDzIoYJitTA
Zzns4Qug2VqQTDfX77BRrl5DeWv+Qf722+d03F1kulxD1Fcfsp77ZZQzpg6yep5bZ/AhjOANOURL
9VKHT44qka+4ceYKcgxD+O42Ki3sqVDzXHm24inpooVnayXP0OEqM9Hk3jupPKOThAdQaBL4jcZ2
QkorcgLhOv5N9/YEPtzLU3OMRVy8FYckXmENgpKKZXcDI48DnoTxIKLylWw6ZkHGaxDfW+jshwl5
UC6grIoMTIwNCTogQY6W191gwX1GmYjb0dWgvEObMNsyS/kvNtHCUounWv73Gz8jd9N9+vscLmMg
VnV/Q2IW2/WdXEZjF7Wq48yGLRNQK6Yj556jcPVmrgjgJmKgh+pCecFxdgLYQZkNNvMgIjOZU2ZY
/0br5c6xTcZGEf2kxHq/kIVTy/vHBEASpkTNXwEcmEQIwUbVCcl3Pj19GK2o/DROFa768ZzjpMz1
fO5jI+DO3IhBGnsq/3Mc68hyQet3Aw5XffEGJ2pD4x2pWOWQUoXmKHXgTp6ypmrbJk3M73ETbO8v
0hV7FDESaOqLwGPDYrnQ9T0uNC7/RpecOvDQIGUUs0YCpiaBzT3xXc0dZiH3ygN7WaSvVAPaHMnq
S5vshTSXbv7hqQSorDJRG/SidN9BOFWBnNL8OgMtqXSP4ECxlYOYglNh5/3seYfNegG2LUMhhA+I
42NNTScvRskEDwqls5C4h6yh7+CyytvsI0N0H8KdSU4K09CGPGVRKRx110vsVJwP2Za+QwjCoexv
/KZnNbAOxCdlFoaOWdiTi0zkeCPBF0mn+I7+nITOmSsw5tZL/U9Q88ZFmtwDfNHb9pUIoRyrD/1H
8+uShN2lAZ+QulpyMPIMpD1FlY5sfneHeejsRdYXBsElYrZ6Zcag0v0C4sDzX/IVIRifIUbCx06Y
1wccZwkg+tJOyi2kkpZPwhzu0LUNpYNXJt8IqtybvCT0eeMJEn8rcDlkUY1XvMIcOBL5xQc+XlCm
fY6w9rDchpldZKT+Z1a2Kxnymg3yEu4PWRdTIXcQtvaD0hhmWZIeQfXLWNHrnaJGF/JoLk6lYpgS
QUUmsSGPSSXSylfjB0rzIA6HsQau+oQ4sEZBbPt5tmwl+7A5h0MQDJzEaE+z1tdV2SVva9hBIZrG
L5Op7Ohvp7pU/jAVGKDy55nHi9Ye5YXc5NLNOE/p0VFEJ4g/BuS2zhWi+QFkSnCP4v1PkNU0TAb3
wzcVV8uaJmRNlLThrMJSPyNsYIPauuGuEEgXgbEFcehwjicYIKWkUlh36ECirrAKHmmJpg1mnFCe
NYh6w9jtOlLbyLaqdpkP3toxKyDvzmT4viYDLQ3fGf2o4EF/gCFXepoKUmims/miqNgGmx+dsiZo
I6K4r2Zel8FIJNiKziYgOplcDmJR4bLxIePa5DL6otVgY+sKcIwRRawgRavHIFmbwxgkAtAlBHWg
+R4teTTktyy4PlBNFJlWS66H53GGYA5NpFz3m5nvA+NuIQj41wqAiixQywCw5v5nLtWj724iybGj
4CF9hgV7cnTmC7u6xjy3wVNOnMztZSMOFpI7fbFvkrLAJ8qzZNGh+3R2RyDsMvrfl3Lsas+asbcw
uhOrkUKyAgH1i1Mu3KjCPepj2uI3iDeF3b5+0LOxmAe2kR+jyZph28RSW0pGU2wJx23zIMuGwQBc
Y02r10cEvJGlXU6qwWOWGVJNsjE0VsOwX+Du1aDXjkda6KFaEF6cBdtPIfwSst/9M20WBEsdyXGr
962OOTOHxSPzE58qcz3kJw8teCPaDX4jc3K/1rKvO4zT2xSWMjelwwwEAUd37ZAL5vYKIIneQpi7
LI5+kb2plXDk/d1SFji3k0VzF5/4bBxDCa6sIglZVol1qdnYAXG7NOomAtqJdUhHC5YV2Kgu9JTC
CEtQG+czKijDc8SeFB5GukXbolf6bIBOld+Y3WevHJPGAXYNMUGVCPSOWH++QLWlPcgaZNUf/fOx
INNJz/SgdhIAOvLcvJ9oE5BsS2Vb8n3wAxbilh57Dwt+7oKUlbOZ9owXVxl5mMrw5FfHNQhbTNTk
Q7WBdkmvCC0YVHxtC51ULlRk3OTmK8rTycFN7iyltzp7Bf3eeAd8sGJi915NS8YtL8w7naIrnnUS
CqymkiTnIsDTRVEUE/zgMc9uygyA/kGGrKeVNSai0RJGCFHUvMCHclfNQMXsQow5hWJWCZgkv4YT
rh0epUpj2UWrl5b6MgR7X26ZgNmVppvQshB3IjG7u1+0MDuh1IdgW4C3YMF3hgvYhrWJTXHsF/4H
zwrx/hNCqsjnTfjm2rH8OTTRoFxPfkmeoEwcuF0a8EZ/CA6q37jPM0vHtFIgKv3E0NQ4sdGkZrfo
rkyjjlEybh1WecPMfhqDjmosilv8YzzVtM7VqPoDBKw/OYuMW2QdWHWnqK6zkeiIhbYQU5ETAou1
SmUPFVs/bqPKa66WidOQa7R3s4YrW7pCts+0GJvRS9esB1j0Mki8pWnf/EtPJ3cs4md+Q/8oy4zq
WM/85MlOzcSPQBjtqGRurIa8J/fKtCNXlrIr1QzfibEHHmxsRbt62C+CkjK1GA69HQnFfUe8wPuT
GEfPTA1+3+11yevah1xvSh8ruWrunWldwqldc4YiSEFCawbmzhr2xr9d4SLM+sYA6fVfeRtmUO6r
koobOtVCII6onJwF7eaZtNfpOJ6Luf6DtLOzMs1xxzooj1GLiCq0nvRFlJx1OTH5Ry5runojfnqM
zq7suCQnKEm0a7Jfc0qCK25cpNBx/h/XvivhBjuWfAlgf6zySF/pgPT91WMXdCYB5fGeaAIQXZdo
A5SYKG0TdMXVtIaYP3P0NuEU3bQ+JGRzauCpGpN2bTDH+laF8NJD2FuQlwACVWjujPI3KqHWXCxG
h9rTZI9ditpVJouRkp/0/F/bv2h+Vgohp8nCAiQ7Xk9aTJ4FiUWcjbx+biwi5+Nlt/6dlzkovtRD
dSDJMvEyOF8b10jdClyfetupwHKVDs0AjblVBqB3Bv09YL4fybEbfwWY7KJHwSkmQTDikCyarPUb
R+z4vHUe/d+KXRLkCIeQpyzJGXKDM2y5vgAM43wYVhCnAav0DCDBZ67bC/oRpkYf5f8qk5+Lzjib
Mm5+kt6cwl01b8HOTG4EA0x4jQKq+pJSuco6qJFGPjrVMht/GzROIEtzCcpkYgsOnvW+suQbCBtl
v2j5FNRxPjU4LnCCOJEeFrQlXToj9NrZQtW5bez4vnCHTtwc+paYTiKl/sTgLyzcZ139y2S0U8bM
1IRbzUvO1jbtxfZ7wXpIBsdTL9eUwUS/SjVuxUhM1x19jErltwKmEmbAXrqrBVhx0kjnCu9TgpvJ
HjS7SDrAt9enutFyXskIWf9DDP4D26AUzRe4umtGLfygFd2E0uACDKf4a2RMbVP0kDOIYIdlEZZO
i6U7ZG/1E1AYXE8mie7SpBBqS0lanRKdfrIgxOFARwHwBOLbI7kpj9wsy880BaAzf375+Hjztnrx
dCMQoDUE1xJBBneBiBAJOlylk2+nPe3qfNxhRfMMx4vgwwtramNlndzj6lz/BLJhVn8NpakTqFla
5+ll+fwZPvPsrlIDmCjZj1s0PrGoMjHPefk4PO2PUrBvNMN6wNOe5tLCyXdgiS/ZZFMoESkxN7ex
JZin04952xfVw0prQjo3HzH+Qarahl/4AKrCekPT6B+eV3xKQ4TGsl63kZiT38X8iLg/CfrTtrgd
tm4zMFC+mjCeVZCKdbz3/hCMXXyvEBdhOkBAVckibbcUu/t65vMMaLcvt2q7HVs1qT2K3D4quxTM
aC4uziUuK+RgOhJfvdAYt6XMiX93LD2utK592DckgCklWOIejpHOficdQi6AIYtYu4iAjWT0FNqx
/PobhqvPKprRnLs8at/VJVL9vQ3FnMJRjoleuBlJ/2iI8o6UGhr2F/IReZWhERaEABdFkmilRW7E
BHspPy/JcvxIzOcZVlUrMiXDCAQ6PBLd3Rz1IiIRSbV4MXcqAOUIwvTrB1HPv/bR2Mt1l/kiB0di
ihNYL1T+w9BM6s3ccLbgYtsqGX1ObDKGMIoezuKlrB+HYcIWGooyMqM/i8XrQnGC9O58RFZJOGdw
z4sPABPBCk48dIPP9F3BdKacRGRLdEgOlsSF4n/jFH2kCCKD4BJuN7Zs7r3aTVWG/AP5wxgeq8t5
m1yhLGNhpsym9v4LQd3MykHMyyzd0/vThMokVElRPiLEBDNTbqg+bUppebmPfrSHNH17UQF5b7s4
ljC+GuOrSN+XBdC+wBlsxBGr7mIyed6FOWeUXl5WFMmxyZ7F+MoMkFzikokUxr2Y2ucpY4i5IGSs
hPY58P+T9dk63LLnMumKvvNJIk2iI35nXMFq75LYsdLqG5HM8KIg3IBTD0Y8+t87Xd/QXTR1FfIt
V1Hy4oIZt/4EuxhI6YUvBIsxEo/rJrwqdoRMnd+XFTe7x0j7VMsNjovwGPFvNFu+LJk1HDiqxRG/
e16bJqvdM309PAoe6FAwPK3gSM5nJXIstOGLXS0LG6cs7ZKCFlqvz0DBzlhzqpDM+VBcGJZ0gKmo
/L7cFGvEA4aZDoIZZamOo75aVOC+dzEBtOyhBnGEzRoxYPBTSHMOOOkSEYYAyo3oaiv2uwgnABCg
AJdLenOGc0/vogKQUuW82LgRvaS6SNgTtArT575jTgqLtTMn0DusY3Ot9uG4Jb2hThJ9kD/MQFbI
0JA6KjdqxNs6M+edgbJrrz6Y7pSY+gzshyZ1GVxLev014YChbG9Pti7YtNdKaqa62fZwC4t/hxOo
qxbxd6+R9dLhKpB0mycBAiTg5svqGatm3GVMUCoM2fHZmPqSIPONarSySptOqnzmRcnujscPL9lH
g2dhyeKmpFoGhIt7wcLMw0087Kc9HCROLi4SUDQtuZzVamy6h5xJQMROlpK5d5YYyvB+6wHejczX
yLVuEliu1CZMA8uSDcDV4IokGSGuJ2PAtMkSlp/hfeBK6s84+Nm3mIlLN8vGx7MpxD+lDvF4MA5Z
T+gCaLOr1Rq81blD5Xmki65dc8ctx6lPL/3oHcHXIbSgMTNsl/n1HKJWdi755YBjOrRYpEeGAZyj
4QgVK8Sm0sKybJDkWrJFKii0bwTwW5mEocwgPmCtiwb0nc/F5FdIMeNymKSXguY3qJ7L10iFxVS1
s1WO01bS1qlbSDMhLFT30LR5pirZiq7StqwgYUjv61398e8MAinIg51JgRjmdO4PX0IhvkTJCXcP
0PQzhkJD/ZWGsScZhtwCNbCYfsnn11UP8VV/9oG+AMSEYvaIuxHHnGs8w+h0jyCxRCd9m7hYpMGL
4aIrRhxzizRN8xCoraZNStr/+smkXav+r6Ymi+qCNrvoJR9ILAigcrRS4wkBUw8k/csg7qW18rfz
YZjWyZVT+m3UcdYHtqwfIoNUnMF3KyDN8GsRuUpoUIJdZPezjzC5hHU22x/m5uR+LBM0BaQuaDrA
tBdZueVrDV6eUqA2giNiiIN11QPg69Ei3p1G8vY2I3iiXvv2xqEoF/k3mExN4sQ7juIxcuG0A3a7
KboCv1PVh/D/l2xcSqPJOcQRRO1IemHG8Bi91ohtIRjQKVvY0/Zm8YFTjzReSYpCWgMT92TQRVIy
xwkDYGlzYoFRy3+bibwbI7DfnETX9dR69m4Yg03RHe+ra0FGbnAedl40SuRNqfaVACc6xvD3qkpy
8b001u8v6Cl5/3L4TZyINfenORgDHYKUwcSSZCVz+qeUboJ1Fk6U70zq1QBRE2wszZzvR6ZCgDnt
druVodq2/iYsiBr5ZrX9hN85my0l8crKTYzhoh6FOIjaZsflvIKSbShA5kMQzHdtNdhzF9d/kEf5
qIW4PILCz9wwVIyyt7K9Yi4a/zewhwakVfn4RIo+5B8EcVvvXu9FEh+fcOJ628CqoLYO82WMT8JB
qmHcWi0RyremJIoDonvKh+uGxaS13UoPXb2n1hrCgBPcABlJ61F0x+kEW31+RIBRfWBdxB49jyV2
7DnYiTrhLaVGKXj8RyWPGkjhedrsvA0jtW0LEHHuGgicbPX6sSGgKGjyylD7ijOhvdF/LxBFXUbi
8oJlvJ4j6ufSnGl9K+oFmcKCJKqCyOxCF7BpRBGG6twjONZtiCXbxX2pdY+ssQSHvOasWYtwQLuF
2ZAVSoDRfLKZCEc9CJlp617AnWMDRSKotN9Fs8dRM158L1ZiA6aByytOucQUxPBnTQ6Uis9MFWfb
Q8Dh9QYnwj20Pm4M+0pjW0UO6fxidr4qo5lQ83ROfFZkVzYXQL7ivzyu66gMg5Nj3K1HdHqW5MHP
vuPjFHaJ7HURuu6xLyOniTD7iKUC3/Anpd2o7I9vJa7ADTdArp5BWL7GyChBPF+5BO3VPbKCMBjK
5I9j37z1ooGTauJuzTu1c0p6IueTOhCV01Yd36QLVAbIrEFPYsTtP1EDY2sXQfw1Q6kO+i1tUnTJ
f9CpurRASAHGrCiSEVX7cqw9LnbLHc68ltOLQYzMl3jOryh/l7WSL/QSXJIxsXpivkfqQj0epvPi
CgvIOAOj9t3Rbd0/LOp+osCn7etz5G68jcqDFQen93ll4qjDinitClCA2SJW28s8o4Nj+SIXGsUe
sA0+cdqjUXzOLPH/QcLmjzU5mf6pr9kW/ncxIuQQDMkDe/Uw05tYWTZ26TV6mGZKhq/FDQBIkLzi
dBo2OdrzEnI/ZlX63okV5ceebRp32Hd9IgIZW3k8VmBeLIUqSyIY6/c/1dH1kQ94frhNT9b7N38J
IRcwdYkEeza6WvsjqnX6Dzl6I7j78LY0CA+I4hAB7Xz/XczW4/hcPqZXnMbyVCYVvCDI58t8u1cM
m0ULySL3e1tL/B32AEg9kcBWrD2J4QwRPKNJNt/Zl8ToRIybuNTgeG1KyXMkruDZWyWN+N2vx64y
9PGY9+1z8r3l+eB8ax/qWaj+E2WNjq5b78tkM5iyavEXDkdKj5hZqcCdFl6J7JCWHzZdKT3Wda5/
YgGO8gqhFmtWM9BcjdE7f8B16IHPyNIF2HWFGJk8VZgBQ0KKcwMiYWEGVXHYMAZDqRCY1ILjnasH
lsZtS1Pz9vWsrQvbSPfk5CcgcykVnV5VR+3p0AllS1sosZHgmRxOiocsxnpayIHrpJrvHb1I/EC/
HMqBbrfWoucHmJWKQ1s8IwJdwz9w+uwUBF333B/qrQnwo0fslptArOMBhpVF9wAhPZOYv53Yf9Zj
LKiObVJl27VUCw/rElcqzGxQcGOBtjoQ6Fw/RaBO4uvjQebLr62wMT3/V9Kw06hpAa6D6Tzc9oYk
lwC1ullwE0ejznbWSJONmMRDLWY/vzXlF71gu3sK52DBng/sW81xwQVPQRQ1kIHL0yqN+s50vGJs
GH4GyQN6ueY+YozwqpsHkCjVtULheuHezDjqjLvnpkwUDZm/7j+S0qprQIuP+qG4oCVe09ZVhwvM
L36Trx+9f+wUDArAIN3v2fYMDjre0uzh1ZLfGbtuBCq1/ys/UUwns7n1gsJ1lCxkWjZPNBekQnnA
Zx2JFRa0zoIiosOMWdx0JX9o6elI7HlKTRkcia38z2Z9olu5R/p4A4b8ZYkL6xKZefjw1Ee8K9Ia
fwXESttkd3/Ocl4/3iL82LizvIvpb7aWSwsLegOjCrqTxM9qImEIjB2uGGfKWnn9wi22cubw0oix
93iQjhxCohoaNwDGsQUzN8rYu37ybzeiR7i4xOmH9REIctLu5SI2GraZc93k/3LEFTx4mw1yviRq
R4bINnMyFw8X/rTySF+Pr+HeTwFGCCHsYF5qOp2jvb+2gmHAFhur+VwtGAFJRhINLtErOhYuYrto
UU6h+UcCIeHj1dHr0kwtw/PwsT7A7DKr6ZJ5nugn+82wQKqfqhoSVLlIMNFjLO832LCzfMfd0MGh
PpMFXJ5sWBRGjPfJf0QlkwSGw0AUwCwxZCBkd0HlzaCmuDzQQR9iaRqvNdMyHCjNhMe/4KULRcrH
6sE20Hpa0pq2b2V1zfcWqESCc1TUuHMshCft7PT61UZ2eS9HjWi07lUrHAP88zc1YWBv6l/qFqP1
+1LZwHsKgsJ2TEmM1QKaakWNkwxPKG7D1w549zTB3/G8zYblGxbs3gV2MXlcUzB489V2I8CrcYAb
uSYXONEEoCiUKKFqe+0TsEx+7gTUXF8/bwQSSWPzUxHG8odFQm9kPELxA6jVu5Phgm4DzP2O2JzI
eAmL78U0G+ZByn8EDrqlMd2IdElZPRqToMuOaAS3KUErei7f1yWCYrNu9XI7HhIuksqhYrmuqHlX
ZK/s9bVVSqdnEVQHV2JYkAIC1ww4DkGHY6Rvhhz8Z7fwV/BSsE4e9OCAp/TkUQ6KSbKnhhv1cplq
j59NXeyn6GYX9LmU+t0ZTDDe6UvCVO2uva+VyMxlnbtyfdHXfSoFowN/h5F88XEzcniMpErgGL7g
ad1cqVNVVLNK9idH+GTs43hb+n3cqrMr6S2xpbHzpRgC/AbvjgBWUMHy0TzPZKxKnTd8wZZEAhJd
wji3Giig7aLF40glQoW2EU2supo/83PTLWrJjy9oL/V3r4MFvZsxKt2HRMHMGMmZPgqr8iJNj760
DU+/c6fOwkVRqUeafqOxCZd6YvSdmWiJ6Tnr4lFHBJtalzhLHfDkbhl45YsZd60rFRzSW8VsS7Vd
BIEhOGomFcZYqx+Q5KbNM0oxQ5jTCakbUIL8TDZTZHxbSOuCT0coSqBsZgGfjxV6s2dihMGTYIMR
GNF1RK2QH0UdOszlt6rHiTvYc/MY8EXzaIp/Ux1PdKmdtbGNcTgmsGghYAU1oHo9dybqgeK1fdzs
OwBnSxVklkOjT9/KwRxJzVU9HINCtUg/oDB7xD7et9cqtJaMknSSyn6vi34Na/uhNzsPX+mFraU+
LhUBVDpr4BNlBn86889T1OuNz79ZlRDLZtC+rAMS/f5OiZXUqzADf31d9HX9pdPLRAzqPsuG1cF7
/einsKySaDB45C7svvCPNSnBw9foJ2nxb264FW81im7mALPPHVrgjcL+q0O7QNhUL6i0Ld8umcuz
mVUvtC6MiLB5Qd5RJKlclO3fQKwEgMSrI58sSjiPh0VKynWDMuRSGGqDyihkaynLl6Hx+T1iyAKc
rVH9IDHo0J3sN4fuVDAAw9dltYFYDd+jyICiG+7XmFH8basNXDr3hDg/mTLiueSdP1Zk6Z8GQiBB
MNN92vbPfTGEAkKJjRSHRAwMRir8AXAI/fg4tKIDW8Gyi4LWi/glCzUZ3DT6jL9KaqFKim9Z2Vvw
7H8zSYhl8f1HqpK534+FPr1F7U3CIQzXUNeczzc/0e+qtXy21xwEc2gg1mVECymeReSM1xeaqdPL
uX7gum8mOkVp+eJ2aSUf6S8qfJFuaNPbchANui9dyZzghK/b4a3/njm+cIUC35KQl3pAcwA9ZoJb
vfqtr55PxxWjLfjxftZYCJLVbIFap9DoHkxCLGZ19HBub75vv7DJfXJg3nuuJ1KQdn6qDj3EAr3A
C+pBlWH0x7ESYQYqdMjbTL9Nrd+SROwWVR2ezlYRCc99bzYp+Cgim6kON07UvebaWm0NUKAaFQbI
ejN2/IYVApew0UXIYBdbaw2w35b0T9D2hDXnezSHwIu3uJxv8IIEpdUJj51x4AkXTL/ojRTW0pNF
pxM3486ju70uyY1/ldjo7K5aSTIK0dcxfWa4ssxIobw5zrWxKlrkYZgub7RcS6/NmGm/1Nnl+mJU
vPmwgqy9D8ki3fPWeTqCGQ8QiZzETsUs1fn0yXq2m6zVEaqlqZgdFIQJ1TFoq248izPDEvtMSpBd
oN2SKCNx3FWrqNcNsfFJBgmCON6BPWB9f34XeZtlvMt46/zigjC7hyIsIiRHVEzmFcpSs5AWR2S8
I8MhIbk4HNZ4qe6AARyOIQNhU8R6q91FTszU6klWrg0TC6ZgVfCG7QG9BPoCZsYWC+1Ip3dc0cyl
31Afuv3+cdhUoOc9ODDTjQ7axlEBqg9pzy8U1z7MUL7G4yXjaifaUOJlZEc07bpV9tCfMr4byFBG
47wtSbgg+R0iDHZvwR53s1Tx34GM+OX8cRiGRh2nhXFNOfEU/FN4qLvtN/735u5vLXIJ4R4ICnyi
bALd7fYozvXQEZbTvGqWpLMuJ4h3RBz6IlGbwq9xG4qUAcRCVbxeEfo4NvkadDEvN42SZsA+eadQ
QWNLyPCcM9rjvwMXXvE10++q/N/K9P79wvFrvofxlH3xTAXgbrCIt19zJZsTRCKP6hOE5jjGjXvg
hBWWy1Y63WcJ0IarYhrahksPlu65TQkTz0PsqF7Rmj5psop96hbPYTV2uXA2Z8RlRc71Kt9v/fBx
E3jS6BXPbRFRfsK6hJ5G1DB+TK5vtTKn5RIBQQ8UYa6kld8c+t97MB6WcHdRRPAD+G0aKGXw1OUs
9UxyMHY/E+b/BtFpcmXkMFF8XObDQqcZRSSJpSppzyXVF9fg5P1lgCCSO9aCC0ib5jaBXZYGGkIS
+x8n8+3+RBT73AUjCIxL5rlwB706LgY0RVJpoNkERQJ//mWCgoDn8apdjW1ruIZrLUbU9GNOD88P
KKqQzvUJr2cKg8VTUFGMgnkTNoRMeJqDHO1yXOfw4pJvdyQm4h8I1XhL0ySRu83+EDl09QlFgF/x
9EmMPZ2szWoOuqjdQ4JDVKAwo6t6ezMm/GifK1jUxcbWadw1XhmMuvTdh5y+p85x/e7nk/hIYxni
I6On+6XOP/iGj3G4BOOFprcHgBgK+Q4lIUVAnGldZcQ/JINCh5o2cgGORYB6MZi70dgQfNTxiyue
m8jJJD+bEk8trvOYJDqQlc4nOWKx85UBVOr/Nzzux/r8piaWyqN8AYPqxxKluKsqF39oZy9Qk2nn
iqdpxTWLN+qIXMgnydR1bKzLc3Xn6TUVEAXgR3Tg7Z9aV5px4VcIFZ+KSo0KC1i0ji5/rm69Z8Qi
chkQsoVOoiyGJeUdlU3dtPXwDCFs6DOYccFWrx9KnhFo4f4lbikoqDyvms3jNlwNwxheSZcuHRSg
OSj9dTrSy4rOzLVL5hxyWYTLtNwHYs449lqBbT0DYEnOHrUmq/CQ29Ps01zKCwEN9VpefW7jex8W
yWnS4NB4qZLNYThd4weRU64ZbWmzQ00JskgSyZ6HsLXzrGt1fuR2ZwDF6OHbcqcMfMqF1YP5dh8r
4HpWAeY8H8YSHoVE022UBOO8ae3kwcX0Jhble6sxN6LNk2jN8HLBkInFjKd9F9VwUpFQl/cI0N13
y4lN6DpHhfUJW75tvGdYk14Yhpr6krPrhgMUKe8iMRCrvjcFrHEQGeQXG3U01kI0FnF15DqdcIz1
y8u60g1zTBnpjvWvvKVjCKQPv4spF4n/8oET7URGCwunFyjPVwDXSiwbBpGhAN2aFFucxkbospiu
MgUNsHw7Q1JzHSITR3yTN/iM4jpkglkbuvY3Owqj4+82CM3L310ZPGa8OCPtp8Q9eSKISsv00gk7
thOAXHJvOKmz3CwoVJ7XDcxADOjCFpLHKlAlEQMcMFGk6CI7LOA5qHmEDMRN8gQb74+2RVQpyOAO
sgL+kCJgB6awjLQIPXnGBhsnem1GfYPY5k9So1ufNWa27/OtM2wMVCq5Dox/UnzJKWWlCXOHY3I8
AVFRrZwNGNLctwgO+7zPRM03YE8r3/OvD2SgwOmqDSiaicKO9rCdRyMdlmeMpA3AH/dqpFbppTIc
yFkgLp1RzrXHv75bdT6gW05gLNCn+RK/v5P7ps3XYoMAoOoo7PnPhcs9rCQqL4/zaBjzWMf6hCeq
YtwqPJhtedrrluI7BNuFwPTwF0AuE6jvqEiZNfUTV1RxTxv/uPQWdUOqupmuANko6FXg8mQyDbXL
RRE+DOi+GHF4SZTBPE2Sok7uk5OH+rMYWyym1nQ18TO7KoW9b1EyIRvBg8HQBuOaMcPnd6XyUfNl
chaaPEBFFd4hIG1gW2rjMzWGQHGGmTVRxiFs+Y+1Gt78fGY8PxvwD0YcOX8CDgMF+bjuVdwakEOU
XW6OpiwEZuL/jE4dQJ6cyB93m2NH8GRqWq4eXLgrwCLd3VSFMST7JSGve2BDTuRPuoRcIvMk/kEC
Aia+ngB8qnA8qNunCSuc/cfkaThn4s612IQgFjq8vCIsUi9Ov3BY699Z9bMe937THvhvdLn8Easl
bOZxckRh0qQaiyGpiq+qhksPyy0Oi3sPL1nsKkPFD1ukw2b+1MfHwDgpojbOjpAPEhP1YmQ9723r
w3mhKGt68CBAtc3MNddN7bP3tRWMtKCWNwlDw7KNfVlvTNPz6y35YUeBm7L8WGaGWTcdZ1vjBcWU
PbumyIQ2zCfBwqpE2cQ+IulMdvxBIHKcKv7fBy8dST4yyFIjpSUn+WEykkIrAcDG3YvpwrK41La2
GyZO81Q620yrK0yYYndADPkUYNq1937lf6NAB0LkJZtepaQqJXOi7BcEAKTPJjgnYEiboIytnOOM
gwS2sor2Oljv1eCUcrW3rKfpA4jWagu9GIfYIpT74YE3Wb64NKzJBBBGbBeNIPMMyn1AffuVsvaO
o/1zlaCMisiL9Xtb+V3zY5G/wY9dkUId8EJTA+7W4Fx6Tj+jBY+pwLax4Vhd0UUz7dI54Ys3Rxxk
DrcONkR9hcWlkcor6MgLZnB3rfj4eiCaL6jf+NkypS5oOLa8DpfxyQZRxJZoTwlpGT9Iel9vocl9
bvHTEcc6PtKijC+2BmXbALb5AyN9UYtFOBngQGkvffuch0q6GMxCfCwOHARI3bCc907uEXeVD4k6
CTScTvl4xiJzF+j0te1nedJLaVu9JdgdLwNZyadavjWgem6Ck8VjKbZOvqJrbFFBzZKwrDTdsqYj
2R0c+/Yrx2tUXkRu5uTwFcEabnRaqVOOktcZlC0Sw56U6MtEjZLX9sK2D3M1TXmsKDKIHITohU6v
LmMPe1Il7ufeeYawQ1m27naumLjNwAcu0S/pocAf91Mf3UScG/RATsMHyAYRh2t+ysefm000T8V3
oYrE5IwMJTBmJam21z62AT/HbmXbNLlnQ5UceXLJS/96B1W1gd7JMgp8x46l8fQAqAdD65Qs5qYu
+6fFM29OSYC0AVUeTKdVZZovD5tWX3ShVqiHOA+6E0WHVTwMf3Y0yOFljuTuOiY9vXI0a+gREkE9
X3oUBhdc5cT+7/l+RAJtrgaxIHkqhyZJq+kbduVlozlB66HJyhHD/4PRIoapydX8zwh00i/bnlBh
1ohm0+Z04SgwO0GsypigHnH09XYkRpP51LxCtPe5LIkdTuvffFTW5Zz3SncpND9mT/v86Qpc6nrX
+Jfbr9WalUxUhv24D01FXc84Q/64nQ6JDppPJKKsPCbCkme8EHKT6+pLGolRI8IYAiU7GvJ6h0dh
m1OASmsg0mXOqCp1RrfqIFiRUDGn+oykbTxm1gz6J8wO89bgUU8aEmOl8EEAxiDGgKA9nlu0XOL0
47hqaawA3asXhKJDUcRA0sPetNV/2nWne+Sp6DculuniZaQz6WMGn1Eed/CVoNGP4EGQJ30a4cOk
ZsIxYiOxruDcBH3srNBNM5tOB/HKk59LLPnEFIe5lLjQdcuXNstC9GH88a766z8TRYsvi1ajC4sx
358BiauWy7ghz9Kka8FUozr/1WJ8Gmke2pH+BtyUDGM8OYsZ/oUHREZlfINNoc4d8bEIpUy1IZP4
DhF+zyazPRR+477IfkNxM6ydebs6XofFhFkeFgPg8TQH4FJ2m9zGL07rIOr9VYzpBvR37CwuCfHH
oO77yOf/S6enCpXBUGGTFpziarg4rC9jgBXXD2aPq8XzaDk5BRH7e+WBq2sjAofgODgQtxBRSbhm
pr9pjUGLkoCGH8DkbxjIH6bgkPWSMjkqyHXFCy4fxBB/QW4v0A7NABAN2+BmRKU1SoSOyO9iJD7/
kb3RHWM2pQPdjYrHF7vG/m3ewhgnxUVO5SBVg0ZSSphnUNEhOXE6mZPY6nYJucOjSCX4JD4QL18F
otX/XnuMK3HKVgUGj2jMTkAwaHgbGi5j2j54Hut/LRlUzW4XsLvzn22uvZJzBwZ2fcKSOhq9db0Q
EpO9LCmFWP4fvfSaDpB4vXLlJBzFJK/B+SWTmRGnT23bRHYy5P3YBJ2hbN5X6/0GM328AZr5H7If
93SFoSZJevzy16sotOjfvmlKgHNdppPUSj55SGLUusmnvL881hpqQJb07uouk3qa7sb+9VCSNkQg
sBNzhkXvAlwXfZ/hfX/P541ubBDKdsh8iBmokBr6w/d8nS7sJfvOgZAdmb8zrTJ9wyUUmCtwfh/Z
shIp3Y0yjzsWrK9GrngNgkbySybfw0y3PhIKqR0dGgn3LWBXyvze/4zwSDkweUFyVBlJikNc2j6U
UJyEDJk0ULo16/FeQC+SWXibut3/QkJKMiSIAhYw+8V7Ovt/KZ0z12xAUKiXS+Jq3B5dNMYlVQT4
wKjDy+Caz2mF0ExvYosNAYoeNtqKyVsjc63HkaSfG1pexIO2+XTBk9iEF/ZtrNxILr0n7GsEWvLb
WtLk+7gAPFieRpomzP7uhkI6H7nPxm+Fdw7dMS2TuancjJXTd8NYYnsVP8mBlqul6f3HZisFe6Rv
5r0vYQdVQAjph1zKkAR96KelFc+z9C99FxiTdIEojhkYnurFkj0XKcMqsMnk4Pf9BTyMIaMnjOOi
CYOUi5499O7UuAiycYMCPdK4jmQ3r07YeJ46pD8/8ef7GkW88acf18cqkwk8jEZSwyn2PQae1UUO
e2TSwYEp3xNolcz6QQvA3oW79Ov5YNeo3Ld8uqCV8rV+1B9UWJmQQ571cVdbOq2XxJbzrHdSwevl
B1jnwNMNNCDjHfHR0LLLx9RStEIvwBn3/ioChNPzNCTwJFvUZXU7u5lNADO5tSPArQ7zBAJGWtkF
JlhCCXUibF+9YoLvKrbkTmknVsAvaCr7keaydfpziri1y2Nd+i9DaKG2TGgFDD9OWjbrotMDXJLZ
bPkh/v8XlvC21eOxyzMKUfKJGSmxTMspu+/BmYXA3zBWdbZ752HqwXmhI4tpNmfEct8iAxL8aepw
x1p7GxG3ShfaBDVEbxux5zAdPv6bt49csXO37Z9FrAbekHY8AxaUl1h/nVJv9LJd/3TqojDXSzBK
4KtL9KQ78h7ZcnTC0LWX3iFi9VsZmCDhTXZGRgxbaPCfquDb3elb9m+1LCVHpR/ywZBbw7AloW9E
jyFqh9QtvQcHeTsb5iWFlV8Tticz8JzEABupMpU7AG4VmnbLWdUnOtnA9OJ/l4RSQB3FyRhDWVIu
1eVgLlrXmOOmgNAnCrB/Kc+iof9DlRArgaZjrbcGdjBdpWXLLOtX3MrrKx4xxrATYNhkEesceUmt
JGpfW7vjGrNc37op0FkFyjJsFfA9DnR5OrreR+arLjsUIKXcDD61SqH2bcB5oOTBLtk/iAPgdFi3
NqrCwlDhyxB03jUJYTpvLI0OsiqVm+omnCaTQ5yKjWBVdNpkAOm26SFYlmpfxFl6PZKdfvMEZLWX
qAACRcRKRxashT3ChZaOEQYgFKb/NVrAmcnhDQWIVpRkWj2KMrg24u/l1rtbhwBaI31cxC8Cxpnk
nmi4GsMYwOgVMtmDHKTpCpej5a1uFxi/UPMLu6u2UmAmZhWS8YsHozxqLYJ0rRmePVUtQzviGmjW
0kN1/a+rr/tbu9wMsUUpg7YRj9qnF/oxIR8rLiGoGT6KMf7OrT0x2MRz4zyBjuZf71UHsIg+Vyx5
Cx0TutySD1CwUGXQ17I49PEGUJn2JuH4Wv6WlcJJkS7JKxyTzf5x1GMBM2ytc+hc5cSZmeEb+v1K
/Dq4kFj/Uf1YKhtYihzfZe1nUSNiZ4y4GaPusfZWDW0eJU9L54b/9FU+iQNBpQjEXnWTisaKyEze
/87dedux3AOtNfQgSEj3f0I+MXB38Oaw77m7raBjMHLURfreVnaq34Q5QAz6eO/veIv80hm3x2OS
xkFqwL9Vl7F5L+JNTcCtIvZoRC7pF/u0A9uNfbXrLvKJhGw6cF1qgJn+wqYNxZy6ndU7CFZHCot6
REH4ZaJyIWF5bApTLiGCP/0CBltUy3Ig0bjVXoX9d4ucEERzxA59OVQCwUdOaHtCtU2tTm4yWQTS
2TYzSGY8uKv4UAQTY/YJu7EEonWniKPkbRknbmqIcTqGZWYgOg6Qh2rpm5t6xKS5BJJy0EW4xHJw
k+4T2ZH9bKAbtU49vNMJ7zPe7RqddRoIwkHIeUdgQvl10j/GDzwbFANci3NMZH0H4cv1O6CZqjFy
DT8Z4QMRvbD4yWpvJkd5TqSR32Up6TuaGey9eRyjKABOnWWywwflqWg1xkA6sfRiRNQ8+VpIPCDM
Lss1eXjzDZeMPo6e6UHZP4Zy2EC6anJRvf5jlpOVV8vwM0q2bomjylAVpWtGE8VbsVOKkZfHgy/p
UODYjvKfHUE2C7tN3Hjb3SCcZphY3W+FiCxyoLSvboUGyo4ig7e+AORHeKuOnlzCjrrjrTgBkYMk
X8j921PGWy3NDOcOdiBK5PRiN4f5dcQOkVJ7LolMk/qcGQLcxLcKFz3KjXSZhBGuCvUaSG0bb/K3
6dEjB2yK/cGevbmye5a/LL/S4eHKwxn79wP8zO3kcfegbd/9fsl//gJvqHQJNJaq0bncy5P0mrj2
U4lmkRgQyO90Hm6XKfP/SeglJclHu7OvVcNTruo09B5G27CHVzgtoO3MGbb80Rcza359HvsTQE0g
pfd5lXiJgt7c1hNW7N8TRHmnIM85PjubwlQMll0fmSn3qahpvE2pv+TvjGovCYWOCuWclLQIAQAU
fvDfBW8RktPkA+wSUgtVC55bV4yi6azrdZAkRXfDtRpAKPb67Se2NmPYI+iZO62UkeRPMbmRr30n
MFourhoo1rNzOPOk7PQWHGGKcYhuS4D9YahFh6/g1Gli7dMSNiR9eWVNhmFT+qElY6DH4ONcprnt
LL2NqM7B8OP4HyMAKIVEZNrWithLTD3u4Z2h7wNPUltBsLIVcgTRKEpTdtB8GbRjQKTv6/BPHQJ5
94IyiZgvTdU+G8YdyAkcfoDYF7l7n1l9gigXrXm+rSLSy+IzIXrxq74uDbcM3Z04KzyG4yPIVRLk
spK0eWd7CCjp41DsunLNaQ0EXedzvlhhWk91bvStxDATnBaF1k7OnBPB4TFg5sJbMlK18cVa4v5n
hFQBynBSQ1Gv63VpG97fiEUAi4/fSbdUU322iLKu8xP4BQAr0v4mzcend4sFwWnrFj2iUPKjXshE
+WIchpZuWnOkrl1e4RVZSXRZUNn6g9BSkarB32x3YgugILyBD55Ciu9qXYHEEqtQc+owFp2+PE3z
8lECRK1aKwFHe8C32ATi/meZkE+XZC4xH1BdqOwC24knCqgL6Ptv5tO+qnD6XAoZHnhcZ1ma23Zj
vakkycjOYPJAdx2NUw6td9/p0P1j4OzpDRZaAurDEwd5He+tIObsOcQilMELhKuOGUBV4W/IJ7+x
zHrth74b7NcVjIs9olETMl8b4iTnFUyI4wyUUMZemodWDGbhdCYfJivzM0eL91urQQInz0W26ejI
97weqqBLrASXs6Rd+SeYvLvdfXIPczgXDxSKBMKMt82zmuFH9aKKCHLkwKXRbO1+wnmYz/2pya32
SrHtND/sh3zwJHsmI2Ctpw/ZMz2f7EA9Dp85Q64D3wLJ1wYVkiNvIqJEbvAL/tOBp6gF4NhdgQ9W
5ktgBDo8FjI+i5m0ehlbUrMaJN1dNleNeERecYXvN0i+FOTf8PmTgtg0IFM+PvpmJt6nmV63jmNV
kbPAv23YCDuEVLlw+rRUz+mAg78Pv+CONao/HkuxpcUJuJ873n6r7L/DSXHdnk2nC3V8Pm7l72sQ
qtO8q4R0ePQbdfFMz7nH//ZbPkw6NdCu/TRilONlYJHWaxkr6vlb9Su8SOXqTDr6gL8hWKJ0rnGM
rvSkhRgCJqad2eFNE9WuY0cqhzmpyCBdGspS3yJ7XzyxVpsdVTLQV1K7IGqN6IBUxxTPaS/MxwSi
gp6MloG8jCA+9QmY8ICIHxDLgyCqJZRWRpxamcchqid37kBvjBjHFIFqML+3r9seAShKwmgcZB8X
imtD47wq1VxnY9HtC5R6vf4hAhCN49cbQ/LmPRaU/GLco8EWGDvITqQpxllzx7xbhD0jD8FmJKNd
hWcNRoAuCRcUfvODDwCRkR/nEw9d1eIGpDYfDtI830U4JqGFqf+b1T0xgZH19MHEY4uS9oy1zf5V
KOH/wB0c/LqrEWtZNEy4lOGSpQc0vvkoaANWvSUDk4sUvjBQg46xM4oTigYHWet+QP27iYJ49zPZ
BnnoMMbP5757D9jOxZYmjp0Z10xiMOHu6YgpDbswWDldvklqPp4BJA9qK38oRCJwtNaeuEjT4/02
fGikjzxOP9ELFtR7xgE0YApbcWDqXpw7Hx03xBmfHmpADKto5E2GLwxl/z7cDeZ/mnxPKCyxmmeM
2rNEo+L3S4UQITXdneYxV55sHkB1PoNvFn1PmV6NuDMnTyvugbjZXXvhHjZQTmc5iI/VD0f9Ad6h
YE7l3mRruVhULIwKN0/3vG3yL8yO3cWw46+rpaYgUCQlxuY/zlfulPzqBf05rLwff5uwgK3/d40e
arnVkWkngrvgpl5ficGHfLJ0rJLUDHNkO2LxWs16lPDEE3zCBSPRUh9y8IF9NoJ9SZGFeazqYpS7
OaD10fRdi31NLDh2k/lK0bMTCJ/1/LUzXpIvixd7sNDpDQqV4n+jNiHTBRlNQbyFcp3opLm2SSIF
cjf/tbQMnKzX87D3kpQ5QM7bXAI8MD68LjIq3ZvMkPR2LppXos4NSghA/64A+GcQqtZD+IIRV0Tg
WI6xQPu6Sc6+0xP0UZJUyOq8gh1t8qZvwvvjghDmtkFbb16ATpZS9utwNldpn58H3t009mS34ltw
ptjQxyPLPdnI+7qVtP5Gg4qpzwpwL/hOzoM89WbHkD+NKv3ToM1chEpOFRQiLlI8b6CwvRBC6JXr
2ZkbF14nMYpuzIS2KCmaZHPjaMArb23elMBvirjCPdO1YfLXjDzjCUZFj7dTs9k7ando0gXShUlY
5d3FWDlu5m1mojfBi1kfuMfddHJH87SBlYxqaruow/K4xv5Tqf31Q/R3LNr+DEbPEgru2hrYWTzQ
+qIo5dWQE98FO0II7YaitAYvg8Ciy+IV/U5oOH+4KNsleVXDMrrnZjX5PdGN891NI/cASlgX7xk7
jVAWMEUTj/PLQRbwlaCSirFVt0LWDHGW8kJAO6A8l5IqaTfVU4Mrs2FHsdlUkk6rfRPFAOC2VhbK
6s0GrE32bCjV05DCrFYHD4ftbl6+QsM5R56IG2Mlmw2k/dbmC4GF7eq4jjPb+/EPyDkYpQ6q1t2L
nYUbHK5TJ0EVFEcIWUYlCvnhBACC+F0/FshX+tnoxWzGL+C0WchxH35dYxPE8SUx+7k+6x2SJ+GB
1Gpqxr4N7ytU2Y+HG4vXlAQtaAAlnJGzdg2IMAG6wOrTICthk1dmZCM16ZROOw50qIwWrMyR5kM4
HRnWN6qJUaQyBN3N9Ovt9Jb2P8PJSA1htufmauow8vFW++2NkZaK/r53lJ/qaZgCOTerCeHt/7O3
w+tEyBn/u9pOn78bXNP02JjzN75Q8erSIlydQ3s/8RGEa2Wt+eIqcxHu6h0F453a864mImpPmseY
Re+iB5j6LjU4fZdrQk6FfOEPZrQroj3lNahf50XKocVP4krSLbkbeQEgWI6qYOXJ+qmW17I2o8BX
m2nBTfqxiBvbd2dPgVBZGcjgQB7kyjFMu8H1AtEHwEPZsApXz7LpDLsZaRRbGIWUQ157rZCOdluM
Xez+SH7AAqtb+KSnkHcM2vdJBsF2OcvTYEnrqTEgnRI5lejYewc/e1IRAzSG1VM8iMa04i5C/Scs
FtvvKhlONzA0jQ2JI0hNIhldwD8BieNcc1C4M6QrDuKH1f7MYC1A+x0SdrT8/gbkMZP0DHLXxQ3J
K7C4+Vo0TWIARK7ShcQPBLETFVCJmeKJoTDtt/kjHmxHVnVPxZpzb+1R+2ZEeaj7/8PoUtspb3an
cNyLeHto7GSh+dZuNnRMAwI2OSVPhH21cop8U6hR+Eqj74myiX1h2ruOP+9F3gw22yiBLx+eoWJD
gG1g2DsdBqRqsPChvBAbVrHUpEgrghRl6SG+AKgKe8Qn8SdazUplmUaWpvSnTXBdRrTtkoR9Aa7d
DoDd0SIaI8ki4Q0W9eCUv9XA8sWFKXV5SwpoMKe58ksF/Uqwt1+aXIJOy54ReKVUF/WAmiTjbBaN
lUeq6MOxK38ZhIad46PRBBXl5pWRI8mLl6fTrxbZBDVcWeb5EybbV2VmQIrPOR2CTmGJ/jdOgW9+
Jh+yi6cAiRsBsHOgFlAKTgznHIuDfTGTK+sTQXRC+weXKlGEuXyDUv9NtkKf4V8fs1nNJQHBrgB8
h6yDjk/av8eHtYsP4Nn7AqWtWipA0tiqdc11ceXcHARu3ktgKD7KNWofdeE972A/5LqlctW3GRRn
Nt9dfYm0NOjUmb25NoDBGvEgme0W+/zATW1CA2oal3btSQwHmSSB7qHkcfuN2Q6OEgxixbe3cFVd
hAw/R1dw06+Vc7KZ59ZPAdpYyqJjOvQmzOqq7kBXdRmCTM2Q1ScO2eiOqZvMZsvhpN6wdZiQwAti
XZFGZlSbzPJOMbDYxxkQydmcDlC9QlUEghwtossqlvCvjY1F8l66g9ntaVtZmUZfQL5w4Ka3XIIw
kNIUBvoNev0qLan5JtjgXvGyMYkAiOkmBNzMu+ACRXvcI7YOSXDnGFwFqt7zpnj1k4K42ttdm4R+
g7JDJUsbouf0Iy57LPd3NolMjLrIjaYzZjBtmzJ7aSaa+7y4DoYEoS0NF20CXwP8UVBIQBKiv3CR
fVBlIZVj54n3+hrw475KLTvQJXyoLf4JPzuqZArm/zjHvvulBfT93etPPPfusY2/hbXvWHviTKQW
NE0qW4xBNtJiCm3wimlMikD1ahIa6KEyRTyWDArX8TMQtXr9NACw+o+C0beWC9AWMe9EK4x2nvNI
BNiwAFK5IrF4PDPLL/5e8K8AkJBAo+pdlHILVBNcYvbzzUynJ+DwknCgVs5GKwbpQmUFjtNh2v33
BufRGxqD2Ea+zbYOYjQQs7e40xNiGAmO47Z4SB5R/96mGJzrZNhjXAhhpP7bNJp/6t+q9LL+j9dU
UGMfDFyjT3F8BhR7o3bV3FLvoTPnufvRjit6UVyOTY8X4tgIBGQty+uhzGmyD2jjCuf3ZJJvWkx6
SWyrpNs5qU/niOlvsr32MtsQ9mIfdlU1gj8qmXDixUEaYJF3lpnLBhOL99AHMTtrenbySimGepuP
9dp8pH4Q5J3ftkfmjH537GKSNP4o2pkv1vBiyyBtnJWvuwcrH7umK2snrvAJtxTvRQRCqRSSIg4w
F55l6mMWRJsgP2qRmHtX61T4iMU483V4dXpKIvlspixeQZTE4lVcdZysPT62afVLbgbiESHNmFpL
7jw5EYLg5luCEgRB3umZkDa/c+bGZIGB5tIT2mu9wZX9fCLa6uBC5o3tRwXgnObtvwQyzui7dxvC
ZoHvNiqMzvqdgtfo37936JjiWtQXX4AfJOnLDvd9+PYo1CQzBPH/yWaCbKQiBeADqFLBYHRPn+sy
+MrqItu+VWz1Kbxi5ROxTXg2il1nIolq1bKnymW+O+TweyEx5P+d6nTGDYDh1zmX7Ud+/a6UlQ7Y
ollMMxoqUelCUm/DKEyr6dUnMasNBQ1Z2uzYuN8MTVjhlSeAkphcKewlGhYZoDkdJTRN75SmNh1j
u8oNfrS0I/u9fHGTjf0wXlhaEu78y893THyizriyetIz5++lx9fWyfzAkZb0aKn73hXOZAf+UDxn
JDa1k6niiC+43NdK/kZYx086QPqb4SJcX0mIF38df4nw/YMjfvxz4yajNmZ9qJSfxfuar/6sxbmp
RJikUdul7KUrrw/CD5TpZuy11pET+VBh9ylZuJL1mXy8lq6K6CXx2JvmFzfP7O97LEltqctdKdHE
P8QkzsDkiT4vNJXenrw1egE3NbbvD3rUzjGtIvbb7FEaufGNMWoKD0JSjjKT7AvZ3On6q7JCUDD4
mIoAA20XbhOztBkprANMDwDbga7IC20tSR7ce5p/C1NN/AWeM9cP2XoCH78E7iuXvkXVCLKksdfC
NwzwairWa4+rSVjH9+5UJOsQfP2OMldu1vtjA6OzVo0CwEQhe0KFX3fnxScczO3lRL11YUlfFZKc
RqdAg9Lld7ol5sD+8G3xGS4C9O2hHk1Zr1c9Nm6e+GEqh/dsKRzqzGwbPb+rV6u1b96DhxfHYj3U
421lUaENRw25RVblr/c9gpFRrftMDH1J2mKlOL0c3Egdee7MeVvOaJmVjPX6hkXBqQbSI1SUXRC9
0/v5JPDOWF/tO+RWbLlepAymu+ql3zwwnCCe/9fCHJtkEbnybqZtyTe0IBzCfFi/niPSm16AHNbR
IeQO/hNcnqbbOsLy1vrAwwygQH6OQd8Og0tf17EQUyVtplm7ySLmbZ257WguhW6xfp0CQDO8JKLY
ii6ypj9/DqbP3Dx37IXjRdkKH1YtU6qVPIY7MHI7w9GWVHHAp9xH6z0cq2YnSwTOfyz8IAL19xRz
NfFko2rmwLm/Fuu6C0k4m6NpWij+NJdSG69GIx0H1NQ8jLLsAKIa9M5c2mKASIxEtCxzGqiVD8+s
L6uD4Ipzllgqn1Ec5Ga4OYeEae5CgRPYu54VMmsgActJ75HOSwhR/Tqwt6od4PahfWxb6aMXWpBI
dIMz0RxGjIkE1D6nGt7DgRjLWLgychz0tGwLMjZHVXQZY66hSISsxlzezcaI/MhuzV8bWsdSI/LL
zDYa+1A0TrkAtOn6iCpliQGNYu4QCcYTJkH1N0ZN8plvFaHL7WpAGTMZcIzq1EnxAJySgsTejQj/
GInzu5BhOJ78lfpI7muQONTFUeOPDa35tgYViy5eM8XLDY05lSJUr+YOL05gi3HGmrML0nqVkn9Y
DZL63vq97YlN7YrbO8K9n2IkOnTq5u2sLNgc33wQphKftDhJtZUONQjUbirg2/ZL5I+LYW0mGWn/
7ScvxsGQ+m2gCSy4WPv6X/3qymmjEPfKIkYHRB/ZD/XvuMboND/qXjkY/IF7Ex2acYkR/r5sjQTx
J3S9l+EVrljft11t0EO5IvZsMb+wjW/2Br8de12r0lAxUGLuSeHIDbytSEvcWlaYMScwhnpniqFW
/g4LeEzpWN6e6JQ+LuabqSnOsRdLiKEDOK+e3z8cLHDTF9rQMkoHY35YO1eIRR6zP6lmQ1t/5a2C
kAGgBvAMhssQAqAgvJlYkW6VFqlEB1AtYNs4E5X85XqfCvY3uZ9kuDVjO1ox8XXA9rZTjRG04SlN
xarY3km6DHqFJPNbn4Pbcgsw6bJ3cLO65GtEYCtmjE1CVhmpQKGVYzdOeKz+bddm152lH80cojrv
qo+g1Z51jS59+ZdR0Zf2Z+C3I6I6g6+7/VlXjRs+DMOzZDc7xBq7vWSMM5n4AxMHEonqE+Wj94Fc
j+LwfkYm0HltX6fIIK4zh1XrDldieZW6RVMhqRAtgdsD7ZrOCVYOMRvqsSSS6JAsTRRTKd2grZa8
ml4aSGuwcJjfA7zZMNSFbltMrgntXLCZ0vOqICbd/Bo7fo/vCySdXVEwelngGA3qnmgFOQFhEhEW
pFoHA5K7HktQ6JWLx7cXqTQmCBihQjK70XZ/JNkoSo84TWup8NaKnMJKYswjayXofxbjRxRof3fy
AJWjyvM7hkL67YJLjaccuT4jbnR+l+eHSO68kL5a07bjTwjbHxylOy8NTity4wIeCOlOXnfopXZc
SOkaIYQP7uPRkrXKIY2SEmSwBjnuQBR3KQWwMAV1ncEvsBj3FAL48A5na4hd0piyktxfcvfS1uoE
hx/BzD0rD7uEGJfmctr5Kx6vQjm//symca8gGr7N42oo416cD1BXfHdRKsS3V/hurFsxAnhK2/kv
pfFaKy2AZtfKokkdqQxtHNk8FsAJvWuG348lRJhB+rKCymSLcC4CZgHUUdgy510MYDKgDcYQZYK+
7Q5a/Sp5KiJokJSIVgD9yFGTS+4lBbcaxwuAgyvuXaTyFtSl+GSu86QtnvVylu80mHTuYhMvF1Qq
cSdBJ0mF8FaafeCDLSM3PfqHQZNuIgTqMDx9Ur3cKIaBEiU/Zyay+rZ/POxe/2gCNErWBV+8c8wy
tC5gwok+n43TzcHnSB+hONAzWVDNmdO5rjZ7Z348loy2NiK/22CQC9GYxOrpjRLZD4vSXR1LaDv5
E/TYDWIAnuMh+W/q+zeVpHrD8pS1XlR1cukk5+wa570/l0PzV+cpjrRUZcC5Huvk45FNZIKlg6Q+
zNwuEWEeIc6UNk6WE7RO1hHy6cGNpwsxo/tQUNiBoQ6sLPgnOodMeWKLT6jRC38RIP8jJ/t877ZQ
Wb9mEPwVDtjgJys91ISsL+o3ehnlGI95aR5oiHNatiBkmyi0JT39poUbwOpjCO5UexLmKBivrtsm
avZ29M1RTRQJxNC6RwUN1o5jFJdAhXd4mzV7dAL00b3kL5ZxNs3wDJLs0SMTqDNzPF1Xc5XkTgxa
0MBVMxblX4+5vEbvNsP8inpCOeBsOt0yCyw9ejB3ljM33fzQL8fA1bd698OetUvxgRqbZ7OJ7LnB
l8Kf/NTmzS9VvsM1k18LBh/RF4+0JaZwUekJnvuEmTPVmmqjsXoBQu33iRVkO0f6oDNgLMw+yu8N
JoPbpBQ7AoMCrCTchaWA5US5ZNRqgqz6Pp2mBTg/tWFCcczT39xLM0aFBP/3RDaiz9zrWI5w2nuT
1nwDI80KN6HDteruSAbZ3DGfsLU9Vse6lvpE3muF15OzqAEogMq9QBBx4oWyAPtxLKtHHVDI6HCz
yOhdUOH/aTbmpkm+4UpnteP65Bz8QLhJXiHdZsHH/1C5OhYLJlRKBzlGUB1SMT0zyNgGTpJuwrXg
gCvAHJ/cBKDU6AGNr2tvZPAMOAR/uCDJcGaRkiTRJRLBUOl0Oign2VsjIWazjLx3FUgWmbJkeneI
AXiqix9B0oZ4nfxYjcV18w/dI8PtD9HPCeOls5EBjhU71AiF1DlJvaiGw0PjYTjLDSTskKCbjHrz
mg8DAckZrKSz4Nrkj8KZaGldeVhReXXIjarXN0F2uWevHfe7WQLVH7oOi3KymB4+mEI6vnCrSJkD
Lx9ezl2L3GIFXFCdYxKOKvxauoW4NM/ireNvu664P4p1GNbCYn83NHUiQKGhNWzL0uoTVUI1JpQU
voT8KLM5ORxCKTMcCfFSEtxRIF9eq9nktupf4TCYA2Qw+W8WEuuP8LdqR4Yb/W6n/oDt9Ry2qs5i
nAZvtUSf5zGYuzY7TuyZjPd3iAbIb2h+aWNM8lONKH7a6FEfd4Eo8542OGhlXLOV1zQ7jNXK6Wnj
9oRAdaYvDIpxu8KksfiPh6kGqC1upXCwY6893pmuF42sDWLu6PosthmSPQD+SoR5LqWC5ZB410GX
4zY9vyn6L3FW/EO45pntIdgZfV3yJm3e1VFo4jXfmoLUmxw7PcPdvrInF7rzZTWaP+UerEVR2aG7
43OnkJSfdIEBcIyebb2D9r9NoFlzIC1KxD0TLJ7GNFf9UjsONGIZ4JqZvwxOPpwYUGmVi3dQFShy
UEhuB2afCHOhJzTU12lsbKDZ9hRA0SiDD+ix1P75xJnAlFtY3i3yiTZx83L0MFnGfG4whdDybaZ9
ZkOmBnR4rvAAHsrcOlUNylAy9EDSVYRDSjI9xQMKjVqAkwyGLaaH1rIzLwDYmx0wjKd9YtLKYpC/
oXfrQHSRhGLngNIZZhHJEyJfliLLayDBQt2DhJ5hjFoz1K2upPnpNGHFCXC3p6BpYIvp8z8CAWi3
Zx9CdVzSJUxijIpck+7Io5uHfg1G9q+59GeqXQxbYp/Eh5+Sk7Ge+H4lsPxejuoQEAZEfELd5QIm
88UpkIKatkOyI3AW8ALXasFB1cO242/DPWcS+2Q0rt3o0wiIfXRhfbdO7FbuaXDISRhhW/9c+zyf
3aQj7A7Q6KyUQ0NSFlYPV3dU8dZEoIo/mt5M7mYSuwcooEaAk2jO98o+qIdEDw6AmPpIOHpVvoHC
WztZxGM/ThiUJzlPjBwAbf0KWQl74lSd0r9sjeY25xRBvJvZc5S72nlLD1mlZLivDcWEfvr1Ck7p
IQI65/ITBEC9wPYQeJ3/sKCbsO/ZJdSd5wjwgFj77Tupcpu9gWm2M3LXQJJN1DxsJoBPwfZ0Eix2
i3Tpd38GPM8qp81v4JmkIFmAAP9JpdfLfUhfAhH0MaeHBc8VEazl/EVPuuABoNoTUyIoCcpRC9wn
znpumTLzRwZoEX5JvgXPD6zNeqmQAE/o7V6GdvyWINvw8lCJbCjvdpSg5QobuzAloeuJne4AjQqa
EHU6JW8+F1sJ88EsRJSqitI9HhrqL3Y2XEBePpwSYjz+6124ff7RTequKlfHRwy51LF4kLMW3uC6
Ie7plTBzxy4p3c2o50ynhU36e8Suh2FwFglvxmS8gfdjMmjn7fsXJylIluKD4S/xsKzxwPawkhrc
6ZubuXLWN2I+QFVcPti9nx2ZvOFVGTjNjQSc30eSZ0TqRshiR/pKpzPkOTz/zEQ/Ut94zDxmFE8Y
JG1Lal2FrtzDYGio+1i28PgkZH7X9DXwwpPPOdJg12Vpq3D+l8L07dayfdSAMNmLRLUUnlSel3i4
QAcCQPH+xmJVSbxx0P6xSYGPW7ItNdhQBYvsmqtd7MhQoGtF0u7MSnxJ8GzBgtRpPQ4oM1GUeIZ8
Zo5f6u0ylwjPFpTpfqgLvPhECswbozKi033n5/XJS5LZ5Hei/HpO6IZftoZYqq7GvWPolR3PCwhn
DkCMOZkgHNpNGquOEkQqzuI5/w/G4Mj/1TTeZsERuljmLTkiQUMSxaksIlQRlY+oZcXADot7+OzH
J36ykY3EyyxDB6qArlrGtpe9rUdTnOTZd1nW1YfFcNqNaxES0IvfByMrc0fJkM5Qw9QMuH+QbGX0
LlOHbv00UFK/i7Uf+AMCnYzR7qXXdgQoaFjYdk4r+pLLIPOWjfiSGv4zW85xYo47UaB7OGmViwSW
TkO8KUiXTJLO7ogYWFNZaHs1r+yC2+JkXf/z061a1TIgkHamQ6i0/mMkzBR7ZWZpq2gT8KwxPiof
q2H+MW8OsVTTUelVoz5QV+o8c8FfUgqsxGbisnjrl3Y4pa8zmeFa8L7/PVt9Vs3TbrActTCND82J
jb/+xyLMqtzv+mJ5obFeXT4Hb+0pYUUegteUj4FtRPXhSb6K959MJ/lR3PwabtcS5zKJmGmXjRTZ
JCMncdANgLAcecnlbubIdLm5q+0EY13zdi/T3lVmC5PmLaorFCVUaUT7IpWN1A0ZZ4ECpplDKCR1
ddxDF4vj381QmBrRRiEsPN9WcXAChMiKiZ9kx/yX2pjAyLonV8C4Wl4WgkRgCh5/3Az3v70mrHkd
faHE6Se6HLvzH/pBlu5Y2Ye8ifQ1OAqfAoqUJtbSA7D71qfG72BUrxEAaLlWCpp0uPZ83JmxJelO
v/IzW3zWbsg1b1jBsHUx5QnOr99X1SFwAKTsVvFn5WmC9iPzbmuKxix5p032Trgz2ZoTPzgnbjDm
FlVlXAXIPGjSd0+XrjwhlBSBcwtO7AjTAbdBCYi+08YEnbgrAEekh1n/bNJP+8CLkUyzENyvxG6l
d2Gg2ZeV2qlTvpcvzxHydDDIhFOG55Up+U6okuD7NYsOl8R2ShOlD+HiJ6SM3/Vqg0ys6JyZqgXF
Fu/gksxPWghjVhanaNtMjJGZgpKTLH4JIIRx9T2YUCxJF/M/+9P9FjMlDPMHSMQn9bQGC527wgHv
R8qXLjJ1yGNOkMmQ+pGeXoOn9iBH1NkECft+/xEqVOt5Uck3tKxqTqvA0x/dmlIraFW/+E6EY9a8
VJcWnW/xdaUWy2SSmlMpZlhgc6Xq7+dKShG0AA3ctW3VQT0+UP4c23ltDbYxM4c5+hNVPQ89TCtX
H3LrCcRcDbnF6E5wcCIDnchYhYz3+CFv/2JdQBkzdk7GJbsqqIuY+bVYw7OaE2DmQc+IN07EdssC
vFJegas9fPoqC0zrTzZaFXpUXKtDmZt782FhGxwg/nQ4VhoCAt5Icj/JNfeKzPC7DHcB5zzInpD0
zyvThaGUyLry8hpPCo9+tVbRBfXJFAANvs6xA3fSRQD0FIMiVdOy2Wd2SqH0yL7PhWbWT9GEOerS
ffHsFmZIjITQ2NgnQL7MAh93puqNGX1omaRXfsdN2WBjRRkqhL5/olByeDwwwJIBvWHXLSPfjgou
MmyFgMDWQKjanYcZngt6qjQS4XWyBIizQXw0BooUQMgNKAS0T3OBZeRnIBPqfItk25AJ7bnx/Ff+
c/5DzKpZF85mz2rhIIj5UOB+9Sa97itMYzbV65JQUVLkO3s9jKMu2zDzuK6EqY3Tn8KUOuHW9sH6
RwWKHDm5Xx248BZ9fvfqja1fA72L2WoglLs651kpYawd1+DmHFz3jOCWEcVjwh7d6H9qVcqgsGtJ
Joy/0dknk8dosodk9SjtgVUjS8dhfmD9UzgAZZwZ+Isw+rrjHb6qym7y9A27CBSMPQPsgPYV4WGm
CyYaUAf2y0V7Uag1OgIEivR7g5pH9jA9cZFWH0ysG1dEt333mDIpod9UTlzrgHi/nQsYhgmnUy4K
hNsG7aIlBtMfk30nIMttiO/+jjmSzWqV2GV9+dFxPcZTcIQ7svlRWF75NMHHpmhOba1r1IIrV8Gc
AkUkuLUwoeYcUDMthiRl2iQXSI3MVja202QelF6np0x2LE2pYzXLMkJGIZbwxcsNY21kASj0nx2M
ZnsZlSPFDVvVfv3F+RE4Gx2wGOKO90V3jIWqpoHSxCrwqV/78xQUUaNqAEuIdcyZv4uztkFmAMX1
J06PBC2IrCa3W5omNiePz0pT8HmyQJlttJG1fk95FrLwbMA7EvHUOLDJmadrPYkjOB1P+dNBah23
T0ChppTvUg/sxXNbdp47/Ov/2MzoZVnwwUdpwp/i5dmZlG4Kj5XbtV5PvhNWtbKC2nDsFLr9MwRC
27nYObl7gxB0Q5AhIC7/E1HJzONIDvNlq6/PEt6j94FfxbOi7nUxyVGVFlWeO/H8mHGPGvbv3sOr
gfZZXnyfSMUdJE0ZVBRZGNHZXpxLfJUZJZMi8qgE329Gr5GAHQa3r6bk4GG92yYqhMCZmSDAf+Mo
mtDObt8sTo0y7cHuIES2ItBw8AQRRNoxJbHC8NxA1g/fvRDJ5AFKFr6cBM3Pjd+nFWnelhW8kAV7
kyP/UQlIW7gU348OMwNefbZ2bAAJ3ksnfD7vW8anunwOuyYL8OOn4eYN+WpYlE2ctgQlBRNCiBfv
KVeGBxmSaHAOpYoKMDkenMRHGQGNaLWDQV8AqVREBywWWijHkTcK57zbtubd3nOANMOLbthOOvIe
MR4Tu1IIZNdBKzEsdoTbftoNKJWHJvt2QTv5jafC/nKz0kjf76Dcv563WZ2NRVG4tuM1ekNpoolm
HMnVtpC1GnCNCfgyWCzmMtbPF6sLUO0aKR67uHL75JI8Nbo8FAXyaAHA3aiKUuBUDnZNsAIBf441
QKkdz3QxkT3X4Ry/cgDD3A0TS2LDkbQg6Bkd7lPG99x2mWTZ0/t2XzaFm9NtcJVRDebGUkfmvRzq
3rewXG/DBsSl6uGeVfeDdNmJixT1Yo0q4rI65hjO0DDoD+HBGTJdaixKqapWC2M2MLsjdiXXLlRi
IO+lfHkG3/lcDO2Lsmmxh+6HZM9vCrKDJh0Zi4GmUTtgpXKxd62B5S/2STBrCeZm366JxDnKfco8
8Jn1xLuREAM5oL8ZKNcK3cf03vdwttwbpQu/twLYtD35bKeS7o9js9Tl3N745eRqAg5YnPBoxdiG
Hk9Zh0TPNNwJrUuVNN57vKKeeDHSoCU2v1Zh4c7UHzGYpA0z9s9A7xYy3wK/DGdV5mqws3SUMOQS
AVcM7CrBQbFenBRnXjC3exRSrY8DF4LFnIZXiyWhuCPx0mrJd80VcX418qCtn/DWR7OXo5/QKhWX
Z2+gO7QMQ/rbQ/ekN9fFsOFR5pCwTfuAhctOuEWjkTZ73yAbools4lp1XQZFPQFxqsDxgXxbFpyY
3n9dnUZJd5Ds/nAEPp9RlK0nSq3wVyOJZdd5XHuR3Yvt98WFQ1cDvUO9xkdtqYJSVImmUdfVDVis
tt9Mz3rKVXvtaNLgocY603+2UazZLPYOWWnzLFdAO3WmY7Yy+ssRvHf2sP1pY6tZG8FKT1SPGvnJ
QgQ9pstXvsUeh41tyID0nt8I997C+tIDPFPmGURDzZacWXhSz17YORIVav4pGOOa/MlXWBo3fvE0
aEbo6AMv5XTSpI5YbpRBUvJSR899M5/dVwGqWhebKmYOUA39wCnY0CPrAboLPZsd+O5KzlYZfrg8
XS5tXiWJWsSScFQ3DSH9c3j6TG6qY34z0X6MqlGtPUBO+KxhEgk+veAbAP/fNtZkb0JAgXa6f7NP
g41mXh8U1L9GpxOwMIURgpRsZ2E3qXr3utqp/VjtM/UkQH1tgM2mJQnTSxfxcOl/5aatL39MqmaM
ZGCUNImIaP0hwRmDjt8dY1scZ8wvPb5G1S/PdAGEGrBCEbG3+xwhd9BcVo9BKGUhBJIpI9R/W666
t6Dmjx/ysRbEACGMODIJoqgNaRrV+FMXT3C+lsGwiGz+QRAg+VCs4s2BeEwMnn/uLwSYvrTX8+c+
FgLZUKDXYmxzAgz8rL+vBEV0UdAcjXF35vllLolVZKSikSdGCq3Car/K4INMNDMpj3KIb+Dfl834
62NsbSmqBlN1LEwPgpuYLaM9B+3t7b6awkvk0yLw5zeb/Qc0TuBnpRP5WZNiOjxyC14wHLGEekqQ
P24aVdEDbbAEOQPuPdaXgY6z9DaxpwQ+mHzE1Xk8DU5KzLembbJkRAg7dtYCM+2tgp6SOcGIgc2M
w3iFAnliBN9mMPUWf4uUmyszoOLUazf3g+eRfujQ6nnyyhkU4qNIyeJhyaWnlBj/Go3xoVPVRpGy
mdr6ZEiGWBJhgQHyq2xZmET8jDzspMntFJb/L5w9LC3xlno4Dk/x1szehNOEOtxVS165EQUvgP2n
vikgY8qq2n+J7Dwp1yfyFCSwdMwYWhKJNki4rH/eRKjmTiR8BwenMpLIDJ6VgWquShqdWUA6wDJj
ERfBFvuOQdN6byZk1K/Lqwb2nO5VEmNV4zviHTZ8DzB+SEF45aU0b7wIyzFKkNj7NMlZ72N5AuX7
lj/b9A0V1QW6m+f5y1t76mScj488I/QThw0902ncy5wlSxn9ltcKz+VbjtNH8tui+Jqtu+qTddc1
Hj5ndX2ZSMmruC7yXSBZavBd/zfeYsV6ieCZwDfQ0A4cvqRM9WYtQsahJ7BtgsbLvKjnduDqoknC
pH0/hbl5etySiimnb0cGweB2OpgGaPPL57RvF3TvlNLWlK1thqp8JkCBKZ+yNn+ocxgSqgvDQqGJ
ddQbichLuDQ24ABvGLdCieAlK+ra9z/8T63a2Tk1d8U7v/QtCO/8Z27pjww5ZDAapWQflzS98qtw
vanATcEbPFXqv0QkXSRFLOWBTi7jXf+akwKTXq9VrJvynAg3jxxsFSLjYrETUTAZV4hAlW6uxjAq
6UkvmWow2gHlavr5+0VKGT2lv2vYvS3IITAWDZypqTYSBHWVakYfe3NzLAmCsRKsur7Qdsh8qbln
PrpIUIZAgturvpF7aKVAkb76RVJNF/lrW5mEj3kJteyTgdEDvDqam5oUWNW7Z/J9NR2TiSav9oZI
P4JKyDKz5SrVwiHbGjWcEUMOiHKznW9NpZ7Ry7vMuUP23yP13jt/0HlG91rADi8RnOsDKQ44NtyU
c4IRIm2P0fbg6xNHQAoZk6hNaTUS8K9OJF1c3XuxyOWwdxCiG/go64OHxxkKuYedyC7q630ptXrw
zyWKQ6MAfwx+cTDblZtPuzlTUKElUDDUupLKX6bUkGdsjIjd09/9gZFJDsByr/gNwaHeJzC+pGbS
Li++l03/rrAEi5AP0YYAgRb41OGQdwgKegagA2U67l9g3fXDbVFu5Fnq1uw1t7J3UNro98ZjBE8k
EpJpWDKbogV1AwGLgFH2bk2A2QEAuOGyS9JB/KlabqRsaIcGtyZLxtDr/IcN4SIBuHNa/2MpD9AT
tjQEuuHIbFFBXjTAmUg0sokczbeFA5k0do3SfZzvrG2NDjlRGN7wKp9mv7Cj2VqjeMq9exiXDf37
QvV8oLH8Ddd+y0CZcExs9AjCTKQpnrFkw8DFI0kLsPfalN8BGo2t5c41gBHylFSMJcPEuOTfSXCi
I86nATaTBkbnnWf+UxmH6dSGkEuFPn6sq5EQXsT6WrV3OeL8oRnvjm5W3pwInwQpCAqmtK80Nlkw
mDkvXIHtBahfPti1OAInVLFnhIiBuQifvJiUSL6bWI/Fvcz+FLalk02MODDmudZWfqvjfxVe+ysB
rpAZquyg64FR4prnTokFZoxggkH5nzvA5SP4plwgv3LdBmQV/kETZcyHV9dPUEiKL5RNebrAQHNY
D7YFDHoCPY9yxwmf9Wc6l5aIbGSBIjUqYrkMar8Y/95xmdv0f7xun35Tfv0hw4+7C4L8cjqraStT
tT/rCvXAWikZyqP1bEim1CFPCDWW3DiEH4gLhXrC0KLLfE9myzOO9aqD68aKLl642thLZE7+GcQh
1BQp6qbGdcXcfBD3Sebb73TcOCYjm3V3ya91trMK6GD3B11cU0Rw30jF08U0Ae2leSRdURhGPDJn
oXiqdW1X/O2A7h53/atDrrU/5WAXjLTbgzK4ucrpdVlmn53YV9/mKDQM9+oYpoRy7ut6JvzaZxiW
09UQhbqcom4CsgcTJrgC8rgx0Q1ZyqrCGNg3RNXjq159SiW390/sD5l3YcPk8RCg/Gz2XEJsNbUj
6UQ6Baf2txPBvNtbgILaJTVi2cYXMdX8ltDnlczn2uadv6VTUpZjDkQ67z7YpYFYtDif6pzMRWhQ
gTNSqVHRurcaKXB1pWj0w6f0v3suATYSpBcp0kS6LDuItMb7ps0rxH6yiCc3+PzTN8Vei0XrYv1Q
9APqymFxZohLkxsh0gzOSuYfoVik8WfuLhUPozg+r7wSs9fU48jZj+P6aq13wzFnS3/uKKJXYixf
r8VxX8fNcVnwXL1nn7h/3V9BwK4F2YLbzQ+VbZvd55KSOFq2vQ/z+E8H7F80P6//bYT7hF0SiAQI
uOocCm1tPI3Wasi67/I0yPNCmmDenwTuuFszZMVVsSGyHViOPfE/EjkIkwNKNaWNqq8JYJMrijJp
QoFq2WKuJmjt9AROU3y7il4v4MZUvYwsOCcalRYzMlfRTMOWPsal4gH22drXB9eajwFLRipG89Kk
ZtJJqis1lJRbi3ObdNf4lm3xKMssBHSRprcORRvYDLQzMnB22S8M5fPIBtmrIIxHj9OBkXirlDes
L5aKLcKEzIFOzgd/ITOsqxWLVnwz9cpX4/fET6DW629EG8WGyr9zAOsNi1dliMnR47F2l66W4sva
Hkem5CkpOSJmYt4oI58JMhL7eenrDY+M0GXhWCbv+F5B/1Th7cvVLls8YDS5fmPwat5tMnfE+js9
nGprw9S9XsQG/wPZkJRoHxgI90e9I73ScsWkqymEahXGZ3VQXjxxUcPb4uIQxMRELsYZYbVV4uNP
amaPxiqpjf6ibGMsLBj9rRfg9XcvD++NUV2tKHY1x9SL2UBzllidhcp+oL1ufuuo6whd8xcxx5ZM
h4TXsIA5hojZEiwsCUmtSXo1hx756z31C0uFG7V8aNBS40VvsyPEvR+LHwWMC6uved2Ye7aGLDRS
8hzyDVA9mSSzWYlUDU38MDlJMG11+OoB8fANpT+27x/7pdGyVYydKT9nD4wg41WkDtjTfCpDHSkS
JPL204L25yqSNjrNswEMYEbmw8HKQPgtUDcHlethQvv7kBVOqNj3ghu8kq9SfnNw1WkD4I51F2eu
H1umlbXUivXOuWhM8h2DSjKNCRKupQxP0IxFyiZWjINzI+wHSPzfu5dRqrxbrzyfzqBLWT4P3WAx
ASJgBR0IatNVZvPpI7HYBRQHfiUWcFYtKHn7yhpD3bW+7+r0U2zkWoEL6BsU2NE7y/Fq2BRvhmsp
CRchIN4O+NN4HBMu4m7lKXW7HWhhu64FDeqM4XkBfgyM9drqb3xCiG1eI/hdziU81ymH+C2yla48
VDtAU+alwJJ7D2lX33XAV5EmkmieAhswnyYoPvlNu7nl2iCu68WXy2GLEZHWW7dyM9SCXdM41Htk
t16FK4T5k5kL/Lt6dMltNDiDqo1OGQp6w9Klj4H/nAdwadzpX9+5Sd/wYaejEsIuEErXLIP7LyF6
1Cm9PNw2yd7weOCwvBY2jnKNOVqMggaZN/eIpU95IUF2aMW5yfvCfXXYrnQxZlmCkRaPkifke/uQ
7E/ubSvh0+FVDfqUjbL8nDBc0qGxhWwAzRKKPD8aBuYKPhP1kRF9A395ObVUgYV1JSV9EQHr6vIl
3/5eKpT1fI7I92EaVACZ5gGgg4wrpA8Hdoq1Dhk87PdurQNS1KZC06HlHswsxB4cJzGZlrxKt20f
ayKgF2rCnOC0ux5V6Urv0vWg40X7ZMo2cwlGn8bBp4jB4l9XURutBBJfjujpIl+FA5rdQVB2F4Qz
+3T3DP48HyxV8P4yVC7xye583p8KeRfGrs5PEQhsYUZZ4nQU+LNB/JMf2fcR2GeNj6UPY7rWbHOb
GJU8/fplbbXtQZxldsicdC3jnRg3dgBVgkO9Cxekh0BQ3gT42q0m+YthhJbegXFGHV2qgX3dhY7S
7FPsbwn1TJVCqwjgvkSOzkeSpxVSIiHBlXDcUjGnufdYecPh0gfcQ7EhBJxI1exNxbgm7ZcDDm4j
7mIULz3g9wsEiwp+/9Z0s/+LjL5myji7QEnkR/0ks8FwFoCeWosVvsmdzJvuB/ruynZApocCKVzH
17CdTNAMY4QI1iEnotm4sSqGGBvD1e/Lfp6mgj0FTHmcNzgYbyeI+4oSYamAf2wqkNxnY4axFjSD
YdOJmE0eQahyVGTVLmRCkk50zKp9jVlDehVnluB6QgRo2sMYUyIHqkyE5yOPGcH3kDbLKBzJd3VY
Fj7C/T7omm6NjeD7qg+kOGyvBDm55EcvSkLbFGMpELA6p5OXO3Skz+Z1agPfYVTFkCaAccrDq24C
SaNY2oTK9h7F3tIpyEiAIS33xfkV9ElTHShaWm76ux+sBdpv80DFxB39T8FZsMzogsanbcxFERSx
hOAxbZN5JBug6WZ8xxqhdWQ9p2xIlIvpKOsJX7acg6lZWmxzIFIcerz6g9O+Jk1D+msykUNyhJPM
nZWl/qAvPzmsh/d7WMboFxc4573zfXZCjibEyqFD4Gn78kgPhnkWT0g53wFBOeAcsRc5L9XttljV
Y1Bnds1DrmajgYee5A798H8omObfkl6AkIgGRkGkAEK3BjnhwDX7mgsXUxALBaXZn4D2YkcZ7uAO
lB09nsXbbd35HVCoxE43z/TJABjfTUh7AHMY9Nr5l3kYUx+R1dIFrsyeQJh7AOlhqpuESHCSR8Ly
3ZGOxvJLDx7A5DmANMYvgs2RPs/2ZPm4e9/WyQBBwp6bQl9FR8N2VNblQfkX9Qym07dv27lgwEHI
KYH7VK3TKLn1/yBDj4VEsrXi9pdDjFrkEWcWB19595HUSJ0xF033eYpbvLEqzhv10PbHrkhMJJBA
9cPd2XPS0yTb1IiQAwjUGjCqYFRdHChd44IFjDGOVUhEJNJCnPgISOAXVfkSPdr5FtOZBXbUs25S
lAowhpzFJ02K6E31+eSoM0Q6EvehZWlcoxBb6Yj9TBwQdLuqAksr7U+TQx3KwrtyVDCc2RjH1lm+
WS/9cJVQ3xc2hKRzzJDWZtLE8Ir344g3nMBl8/tmPJ8O0axN4D2/tFD6eiaFLRCc201OjYMqYomb
+MIqNwaU3aFIvflCs0L0jl/INTeKOY6rK8OOZ0MlOlJKvzRimMJ3Nm/qYVlG1Kc+wyvJ/+y8/SNK
tU0aujEBItxeG1z6qYTZWSyaFyHT52q0JYoo3zkM3U+pRK9siN3eP+gfC3B+w0DZVajaFOLNoCaf
pVkaS8gmg7p/Xsgsdn6EcLjMyh1oqYa6fiEyO/u7zdcZL8sk0TyQ6bN7vHp0P1vwmfCGqwsPUMa6
tFhx+IMzMnebhbog93siFebHOygIQRshcZhN+rOx2xzt+vf3VQ32041ziZ34BsZzdRpfDTwKFNHe
gNcmxr4Wxix9pQ0uVU3TMCcX5SK984uXb+3RQ4YSBw6Dlf9Mwg/ls7AvAOQGVr8yZ8TVJsH4HLyw
fCnmC6JLn0jg87ULKPlEZOnDjpx1lgbGYCkBYV3BxgDQGtl7mZ75H5cdHIfhEUECx+sJKgRZTsST
aMb57g2o37ZApYRe4uk23/GK+39dK0HNB74habUSnWaYprhIDQ8Vsg7NPOxMSKYbhR//UxeK+e6k
kp7W5djrC7XufLLAAcHKBs0NGyMSMBmxhRny2A/bbYCvFLj53SXyDtQbb+IuwtT79DngYiD7Awgy
dMOHvLQPtrtzmT4ylYwV8ObVZIORQo7qIP3behXQ1899t/O5NoJLtMLNpwyRvXjN//Z55feFpBQs
CdoqNE4DCzAPY5WVXSQv1lFkM6O+ZIQ8sdqUuy0aHkWnrbq4p9+6YYyc5/ZwsqipEDsc7jcfleq/
3i+CFL/0rEWzyq9MJhNujNQhXBA0NunBWYnU2Spu4iqwv+iNJLbo25vxpYbtEtNDIbXwdkUrw2ry
BCOhFN0IehVyJm+hd5GGPsbQpHfyqDOQ7bBimoS0j5uF7ijlD65W2NkTtfdYQEKU4qnEMt7TWckR
WH4gGCT/ojh6KnibKyVbVV17s7sm9gFh9vneeuaUn0xgEMwWEaN5/Orm+FyMdcALMP/S7+BzOvOu
KTaIiQ4EPX8wPvrlHM+2nFiE/0ZMvXRAhaDIniF7Hk4isk723U+CRVQfMDF0df6GmqUnFhyThkVy
J2sxMRnHwki3hHNHK5PoqHbIuKW7S6fhB3ixCf0/M5X6Ojq7Na266YX1Mcw+labAmtKoZAQaTzT0
93PXl03facukSq9nPL5MO7mutWIS7FYR7ndQZcXjNGxAMfhHlSez1HdbqhfvkCD9WbOpOpT6KnaM
m/mSVPIHAFkKrP5mIMkWAIbehAl1IBi9gVOrkSbwR2CCsUiOmox1QiF7lYS2GwxBwwL9Q38OCOYE
LQXIKRLI01hV8y7COaf9KkbO7F83lXTqSsfgRhzpB58i3UuXFxdPA1ux5G6GQ69ssPshFL/1rpdO
SecQRzJ0hJnDKlKOnlYvZpcUrO3ENM2NqesHy+O6eGXyFrnW4x9Gb8s1+DCK7fbCYyalXsxDo1hf
LUQd6iB5Xu6jl325eVZKREna+z9cGgXcK3PyzwBYiZ2unSXUPHTcfz9XZ0hXOOo2ANaaWzdgcB/J
PEmiB8LbZSKGzvxjncM1vhbNKSYfMwxOyL5h0R2YNL6kKPQCfWgCYOmxWfvIPiMomJH5FHo0oPFo
6B9GeZsL4d8aClWh4op9LPImUpeWv52aGKPFbO2/zTeL3dYMKqdHEIh8NILXFMQwyVhtcFjfINRV
ukK16VrTpdsV1Dbzkr7kj/DnfAq+tU4Oxm53OBZomg5t7FZneYZpqqRc2rwaW0Ui5ZDzpU84hu2m
bfpo0d3AKpdLosARoSJri2vfJVTHlg0k19P0iYEh/zxLMlev2R40OTK9kGDPyVM+tVS0xgcynbUr
x5tOzySFj2HZNJ4EVnNrBLEjdXynfCu4Q8UzQxYj8h6XcpW+L+GWgUaoIVimTRClEEuKRpotEg9j
RXGRS5iyhG8a2dJOK8d+Ge/SJig7TmeYU389zvo16XyFgsiM1/keFn/+srIFj84giTzu1NJcBlwB
yKNXGfGUUyaBGWMmZ2DQt7cav1aqvuOckNMc6irzPGKpLRi9xIwDff4sKm3/UrGeoEMvr6kSbjnK
UEgX9ewcQdqurxQ5PM+Rml2saB5kdykTs1+ev2ibBxybh7cE1eMSfOmcBfZnwv0WDhAqu59pyU9S
D+g4O9BAe7xSDDDckPDY20G7oY+GOJjLM/gorIHO+IJy8P7d/wcr0AEA0D+zkZsj8g7mEeJprjYs
1sfAdgyONiikEHCG3T4RH0RWvLOdfHfQIJjOtdWZgshV6vU57TNO5yZ4NtR1Sif29v1ZCrzvJfjX
FNpUEf+oLxZTOiEmGM/zXt/X+ZBN/XwiLjnwhbPPBbNKe5BeDy4YoF4BOGqSNJM8nCMvb4ltr/XM
tBaq3U2SLPSZGsip76jnihvdV/iRMBA7v0HKt0hc2tS441VBkHJm2cMdGaKMTQMlKsvfgXZO+nD5
ptcXM2xsdj8eGCImoqtNBMcx9Q5tXIjNSu0YGo6qykyB9RwejuwruglV31f/pPrt+0JdHjaVhvYu
XhCABoWixF8pw5MkCfBXPdqE39C6rnyg8pkvGTtz4fnkZIKz018reBvFXBmppvb529VLMqoBkaUz
XcZ+aAhWmjLhqg2SVW08Ugm4iB9NRz7QJLiZd9dWwVnPGRVH4+dwgF2tOYEpLYknzyrC7umAufx/
AWEn1vTMYgWX+GaAxJwArsRfmm75mjfjyp9v94d2ho3SXaWZKHBGNm69AXQZu4lw5+08t2Q9KuFE
gppGEV6VEHae9EBm97sVK4X0B+FUE46FTmNeAcutymKd/Hw2xeaif+wKSXFhIxCkaIkAhGVBLXk9
MG53YxM8j3BlTUBA2EzWzkpCMZ00TO6SS7o6VwakqWfg78qzKE/bD5GhPQe3qq2F3wDjfAx2ZpRM
uoYzoU9G/rcfoChCNbd3/8w3wPYRDP25CJHAQZKPaT+PbG83m4GCORD5XEJo2tBEcCvkXuhO6sFI
1L48bvlotvMlSrZrV3c8QH73QHSl33hQpq/TkvWjoZnMPzlaaRhpP3sPNfq2QQNkUGl162Fz1qGP
BXx5ERQ9+jf/ZJGN6ns4kzs9q3wWUR783Av6uel0YUyxCRiDKJS1bvUz6BZjHGihHvmeFp58pN71
2hgQ+oZXkrAOOA9Qob3xpQbCGEY/wsEmWKqK6/1WATUUHlBzRgyJWucaPIjQXSKcwEZkGXOSk16c
2otBkJM+dm4sNpDduOxdatEObU6NrWXz1HHr9BMngsbZrSAWCQqMk7GPGa2bHhVRe8etMGN4XYUk
GEd3g120C0i/Ht+BZAx7HvYAxWYKz565IljPnVoeH0yHoybDsFLcBeFMFoovGCoQylN0jH4Wbi/4
C7kB0XGQEYWT6fWk4m8qoBcsHTegAREskZnyx5y23MLWDlnrng+ANqcOtS9lTnZmqXt4ovPyKZ3t
wY1HdQusaEJKd0WMVwXgPoyMRVIa9dROQ64eq/tsSVHxY5aeD5tueWA3a/IFZUWQ9b1bndUh4Jbc
g4QJsQ6ijw56TNa7NrdrTvSPNz+09PM2Lgww8qcR5rhszqwtAZ1EAjLyit8oQeVtAna8Cq11ZRcy
ARGQ/aQFM7ms/CV0/1ZamjoRbzdLiNtxjKoo6Ru+/KE2QJDbz7TF7K3klqfmGRZh1KxO76K4v65k
q0AkT6bsXL7TTOaSQWCl8SYZftPVFaHc6eNgD3y7L3+WKpByWzp2+UqwTnY+Vi7kHB7PkO4vQIMp
KJyncaJU2ohhpandAOFpchzfP+KHVH8u5pzcJTtIZ1zOqcUo5PgthsGOJZX8iZiSdnD7Rbqh9Tvf
1vCI6Ng6aA09c++/xnIhUsOnnfFoPkVPFcdj+qvJJPh0fgG5ilTQlDVck3apWq1AiS82Teh3KDos
p4yAaed5WeX3M2qjKeYbQgm3mb8qOOd2TFb2jtvfUPf59dQgpt22FeiT5bfgPFuCtF9fbtGfvaz+
j7dCW5Yt5V+sVK2MR7JUvKE3I7zsujLj1xg9ZBjkVQTbYac7oupo/ffxhKH7jqZ/vH1PKtpIBmfg
LieU+LZxY6g9tCUMinzEjHXtVpmg2clw+xqbhVBfSJTpIqbKAn93phUWteKIGbc3+W8GRK2ZBhUs
SG4gWcWQFqb4fKpZ0/2OmA30QC3kQ0cpU4Q6aUkfCYFT1KXsMZ27Xtq4YxtyV0Xvzl764bIlDc83
w0+GXCZ7LmFTCHXDlRbiRQQYHqcduTcZ18+82ECTNtJ7ddXdBxNVpw94IZjNFiUkH/vUc1HoExHn
NKYoF+cA927BzoMvOctWEXkGGHmnUS4w3QhZ/qDoU7hWYrrUuy+FAMXz7Q/wcILBmgb3TVn2AeVl
HKS1BDw3olpl7Xq1pMz5NE3GC1SXDOgy4d3ANt5vyl9xcsWE+p/VZMVChf6YxhOe9fwQbjWjPVuL
S8cNNHEqo32WOuliGmE3dvHSNoTd8e3p8yRpq9uNi10zOgRhXY+fvIef+WMK+X1v844QVCiRSmVj
5nCswBonchFJ5Z9TTTn+HGLhX76HyykLMwdtF8MN2BrHrdZNiY43w5f+kIblsoreg2j6ee2NzNdm
9srGvfoMEWCDxpe3IoC/YGZGuiC98H3q2oZ5yvUi7WztElPSogqyB981rl4piFLk95rJFevmPwZq
i5/p7tAYPwIuSEc5yT8NY2okaok/0CrglBz7Ps4iersD+0VB2GRwqTuvFbSQ2oBEuOSU8mkVM2YK
uym18Vbal8Ias4vfnRShYG2Ejgpck4t5xAdQJVnTf6adAHX+RLjc5u2St03sbP2sPprg8djT8Inu
6dUzSg4ZbM4GldYzAk90x4zZ+ygqY2PnIIePoel9BWLxKi8P17C9ZoV3zGJMy5yB15EfhreHNb7J
5rRGc2rq/Lp2Rnt/QnjzStTtC+mzQ3MJ787TwvglrI+udyGCLnqaAcMU5acwpLETVG257qc3EJdM
if630Re35sn0GnBy6RZCKz2WrRBXG30VErWBAuN5p+G+qKkEzVjWrQYEGLQ6oxC5n9A35lYXZhbe
njLcAks/WpyyCes0eZx9geNcoOQlNgvj2zHQJN+B3ddvfhCDj9L2ZB03IxDpZoUCkDHhsSCG4Spx
PLun4AeSD666pW+C4DcPDvuAI8TVLPkdOaT/xCwF1g0jkKUlooGtT/xTTseHeQY3W3HbftpoPwPM
5g36su6gMh+gZ5r6FRirGB9ph2IXHQTPkXPIJDQI1IgdG70ynaYMFmwYX7oIwtUh+HaUrga9Dm20
cbnN0X+6GtrnFvlA6h/+Dn0/9fshLEWFLEvc/GZ0r+8FIAzSpdL5ZxKcKDoDTJThdY/kEtMSkntA
Jm2ewnybwW35s4So3F+FrcriDicelMwLQ3gnMwRulWXSSyfVNac3bCmWXn7rMzANbQqkDsKMBCr1
LLi3qWI5cADtIndt7BjX9B8eOytk0NmK/K+h7uq4yaBQKAZe3TIfwzqUnmhOf14/RqoIzBEAluRg
HoOYBTw1OyAmpbF0xqIa8SZYdlqoitkcppYB19TZ+Wradv/1cKDzFqZzkN1a64l6WlDQ/9weyI2B
3KlC+zsw++YcUXlGp8ZgQeHZFg4WiyIA2ZjMAmR/WUoX0o5Rs056j6tonhyFibauRBH+fdUn7ZBh
ln5kWzZwO6SaZS5qQBW0fwTt//s6guw8DUgDZ2hTwhrRuyA29vBHN8Cegk6AyqFDSb4rfD9rB4HB
1q3zx35XdCKBG1e477g4maYQchWJz4onvP1r/mcUOqT7j/WZZ9oY6i15VkCsOCVqQm5Gzyo2EH6K
aZFEinO/Ksp6chYs5kYAGRriYZo+g+YiiqyDW9dTYTG0zCD4W1NUUI/RqC0/N3N3DiyzI1z8nLoO
VRqlrnTzbuDxGodFVWxIKGhAd8IUsnzt7Q6K2/ILsCsWywQIjcN1GRdbX1Xo/cHZIAG4lPGE1AfZ
ckUw7nWbJJhz3OOJ4MNuR667TAvWZGA3Qgo2mNfsJPrY3ymZTlFf6RrHnZtRtnMe2CjfXoVfjGzm
EBpIMZwYhaaG7ntv8qRCaLeyOEdsfA9oCtKoJcLrPloIQz3X4BQ8T6vuUqkdt5UuQEqjHw51K+3t
FqvaJpUtSuXLG1LwmhaWrabBO7h9iSTs3xVAEMi9E+0su/iusq/y9P2swb2lm4m27QCDp0PvxXSw
TrxqoeVg2Oni5zg7R828VKu7HoiUXhH9RVO7qiD8JRcXOLmJ+i/v2cFfIC+pYHGob7Ioy94/uEE6
s0kjsB/thx4cmvAQenYnbiKWSpZ2VTMQAOwGLd39Ir8gzzaxpcNbkB1iJEnUtl2pjI8zfez8ug1x
KBOgoPhPhNzzoyU9JCNyK+yG/eOaZPVLbKFEQxsVoBYmb0vSZa6U0V3DAqbI2dIuaUNAxnjlBarW
mqj4MIv4t40BWJUuMbWZdanDtlfoNF+7CzDzQLh5yYdZTdAH+uq2AXgCsF64jFHuiI0oWKCHhVyi
hAe9k2AT30pa+/n24FGBT4P7qbE8EcH+lZ3Ub+8xyCiDFyfQ+OY8Zw4Xx5HD7o8cwWweIHUy9wQ7
HaYklMIyx1VNF4633MeZSXVcxSsbpaMEQz5uRZk2yF0BuqSxHwOHPC3w7PU3xdpxuk5ySEhDXL8p
1mdZNNAUWR/8oQ25TigrLp1ElQz9KtI4ClMAZ9/ANKsQevietLKyFwrVDXOIWIM3KbuPFINELEhN
Y4XdhLTaHdVkRYY9slQE+JBhCdT/+C127MHPx6Ho6oF2I5rSYKuIqKK2hZypWsqjHtxY1tN/2Va2
Tjwvl2rNKKQsTK2qiJEq5/EbnWXZa8vw+3qfthCUFSeriazUIn4NVNtX8Fd9pgEDYe5vqLQuVlEN
gLu7o3krA60DjSgPDmtFnGn3bNK42+/sGoi116m6+p6znLrNKtkQK61S9c63LmHR6ggR0yD8aUjA
FAW8T+k1yfxCXuZbv9NlEie1E1/0No0o3PzQ7c8bycuElR4JOPGY5Wtf/pCSH4mdv8425268mOXT
AJxyRUFn6ARKSO9AdNt6wwQp4T4ntg9D7WcxJR73czqzndcJtOhfeADLs1FjpLfvEVIymoNZjfwB
Bl/lrIgMJ5JGtwR8O1sr82M55gdAyUTO3FdShuPNXr4HW2vzJBLOiyxVySINASs92L3sPqZaouaA
IetrgF9OoXd5GTbKENG8T3rRORbgRFrUWTBknfxL1XzTHfjPMHMuQQ5fcdkeYCjLP3I6s8BOB29v
BHGzX+f2AS9iktc2+WiIAwnt8dvbWnHSAR4Efabt6gy5mxE8ICGQEtQAK/HMKIorjenA3GZ/hPjc
ntU/pq3ngW23pUeUxIojzKaivonNqfbNg2VlrOyobGQkTvhAmfTPoJU1Pu2o7votFz9I8I8lINa/
qpsc4RZnIjW0qVutt3HbVljEWq8Dxu9lmZgRzwM/gEwjXV14pFQISjHYpdudaz7SrRHgQViyetBS
26ShDfF7pzf8F9mflLmC3ZWD1EjKWVrjzqh1UcejFH7UZa7e0H9d7LyHKJvQpC80OZUQJfJMfeaE
FU4/+7D+n2ePItjTCF8vBeM/1mXy255qmXFGQ37e6NSpKoF/lIrSYYYiodxeyu8jYZ0GfYHmvi4t
m3mZbog94RJS2fkQnqb3J+dhKZ2tI/Wjl7Q3tX5g9Dxmq7YnDzjxqSct9x7DReHXkGTF7a8UCDRc
76sKb4LUvjB/lT7LarzlsnlvFY9Yq0z5Yp3MkYsMVN6AaqRxOT291udksYjwqUcuyrSFZc3aytA8
Do3S857hP4j4UVFXCvzH037+aAHT1iaHiia454b0W4xOsmuEjol6Q6sblAU+dahLV3nkPrMy90Z4
cahNv1CbQ9SP/jM7clYmTfyAs+cyN6opx2FRbP/lE4AdGR6+RtQMGcXy7Uz0/xNfx80rYNxOnpoC
lOYUlnYKO5gvEwI/IGqnMg8lNLpiOGtlHH5SGkgLMnrQUe/B7ZPI3wbOHaDwDJMWCmbFKzb5LxeO
ET/PvtxvCEP1ifw6a+vocl7B85ytp9ZkK0gCDs42ck/uUlx1XmO4v6aFKSmt30Ab7FYw0UcJLXcK
DK+M5khHSltl8gT6vPSrgbJH5Xh2qpG4AH08AMNgQ9Jj4ocz7h4Jqagkd/ZjG0wsMKhmssVlCD6r
BI3XinyMHUvGqGnvpKCH07PCZ+d6N9Jpr7gk2AENQokch5cbsuCCOrLB02JtHkjveNd7zwChRpGE
EN67pJ7FtW7yzhV7GHWxH+HIXh0wwZd+Oqi3VWePgOJlmBFZEbBbBPCMFcpY2hqp1QH0+uHA5pQt
+hxmLs359eY/9nC5O9QbAFGA0zQNVmWemVAsxsR0r1Jv6dfSBiHibaOfFxeORzSaOUIZEZeQ8yZL
rg31mMTnsyc2pFpFnEAk9hHrdqRgn5bIqmy7vAKhetTnjGrVDIduGl6PqM3ozeNu7BxDtPJBzIGz
1W9AAaZKBMbGCNG342CdCKFsHBVx0/mpj0DAFJbj3h8tSTHi4wF+7OaCI/oTU4bpmKqGVYN7/niw
AaXDPOhR/R4mAHVg8Wg5mCEH3i1xEa7E+x+j3HMsMHaYDRjRtXdVO96lU+p3K49YqCHKbxaLxyoG
qTppa+qTNtRH0Z9Cj1FICL6LcEjzoLPStlVgkCXLvApjHUty/Om+u+jt4k/MhNJ7mEnkVMRiname
ouYUXNhF1K+jNgsyKKbQQwtDHH90lSWdeERwSTiz3asE3tD65+Np/SkNlDMCsNZDTPg2i+O5OWVY
E4EwLrPWQ8GWutyxiSgoCOV0Em7pVcy8Ohb8UzypoefGQHchYuEZl3ncAiwQFlPpG+Nv+iSR4wzT
EqWv92xObBylDOtrDeHt8yBpiVyVVapbdCzYTUbXwSIm0PTCMAZwk1GI4gctzgZJuugN7huQ6UBc
x9OWVi2R6F2C1WJGsMUiDRNYkRLVdVqr1ybA+dzXSez3RiIX37Kcs2W36ULOq8iPRaeIFQmxrZnp
PGyegWGNtgM5Mlb9vRfgHbajA13/EfVH5G7eqFur5Ntj9b7vjBo7td+k4yxzrQOlTlsMC/e+hRcL
iuB4DOebHab6C0Dw37gNuaGh8Wz8VSbQXMfWSR2NhGwjCHjH3eKsNcaOhGmeQw55LB3ahyI8TAbx
agwnsbFDuAkZs2VPbN6/n81TkCAH0Ik5NAv0iRrk+tCU7+fuS7odtmguXSTLUU+zGMzuzUIU05z6
4pCden7ARdGk89ZlYf82hdxmvflRer+MfPEGhteoAQsaeZEyU1neGe3dyzPrmwxrwntwTU3h3gcL
AirstWW18EFV4wMtOxSIRbIlQU0yklDZnn9fVk7fXkwEHx81OfOXbIZCJ145h0XW4Paqpe6Sk6FQ
o7HTxJhtWnLoKyOtL6dfJFTQcek7vFlzhtz8Y6C4zfp7GnEtLrfUaMc+QSz6yodbvIsAwAxDCVJm
6kk3jSMcbfsE/UrYHraW+L8QHxKBFvXadmxeuByzwAotN8WGyXKTY/ShpE/ZfhzipMQl2rLVDkom
wpS7Li8+QtlGx+pnoNRdCWxwMymE7V6og5mpfj6fwzLxLuU1YsDDJYrqIU+v3zSkBSFcaWK6+TBv
JPGDmyXPNzxt+bSaoUA4/qQ+Ag1AbBlNVK8HKewB63c47brsaC+vss/9kRVEkEw1YKDGaccaT83I
fhPv+U6ojL2NW5O8DYwijWII6jdfj6OCvUgVY0qkve1bF3lMfohATxZK9BemZZXTi1pEakYG2EYI
w8McpnGkxb6urO5NuIJ+TEHxGmyySvSyyCF3Amlf90DcCYm6YHt/FniAEIOSTXKU08l+AbUrlAu2
RLSEJJEFMg2rHXakjAnlb7Tsc9CHznlTNW2WPrJ1eUURuNKZq8Z36FbYk/SMiyTW/5VetzwoJK5+
DoCuiJUa7x7wh/TYtNE3rsUOZjHMIQeR2GlRxfmF0Wn3VCNu9Wxp48aW1+sy+cITmbW7t1LdzwaT
hzPJ2n6q7LqUpTATuZhTLX2zgP3cRrEkGs6SoMgOaUhdQ3WI5yEeDTuPiDG4QLPUaOvNGG/rCO3j
5lZ0nDN+bS1a4Qyz4qEZ7qOQv89+zJRo0uEtBQrXVcP/CiuzDD1VcPL+Rag91nlSWVV8CyudAUsI
eG10Hc2BnqMFTb5gMGK2JYGORTAvSS6LFLhYyQms3j6pA0+ATMKLS+cXa71bjlAMN8+BUMK/WSFJ
bdN1iHi7SAs6Tz77iKRKpiIm6bTqFWR3wkh/mOD9Mzk4sdrbex9NAf1BHIBycUyDT1AkfcIi7JzW
9hqxE/YMmSPV1mMuBTY6Qg7LzYevDOzMbcgHCaaTZBpZmWF13yF10VyQfecychmDihA9Aih6i32Q
DpqpSuotALeglu8gdSGH28bv/1dE/fBlYiQESP/XswVIG8SjMRdU6lUd0Fh1rg0z1bt7zTq8Ut6M
4Q5Hpw1XUDUFbk/cJRELwLPJ+ToKoav3UypuJORMOXYv+X0Y8gDDKBPxoEHCoQgLrLXFzmXA/iEg
S5fFNvU6OGX9SeaND2gRcQQNS6LB3hNrrju5Gtq43q30dy7uaKlapLxL6Yf8H10oRD4GdQ096ASg
ceSVfbmqBz4G5HiJwDstMqLj3m/S3pjVx8wqLG4WiW+DXxdXOGKdX2VPK3k2fNzagONfvsy5ww7G
+f4qFKzD1qktss3fQ9eaVZ2nVtDz6ngCZOeIzpfZC6apbD7rCDVtKpnHSTtkloMyYdM+nP5gzuFk
MB1muc7oj6OGA69uM3IvbGXk9ZG99hC+X+CG/AZiFVPX3QQX1kFULe8alaIMES88cF7tM5FijTab
uhv5rBYNha1YlncK2wloTlRq+iWssM3NCi9wER5+o1droQztQU/RNkYtECT4dq+W6MAW1YBKXpbr
9LjbdwRK58/eZmiJTjFjjXDeGnTHGJePOcYM2dlKD0ldrEtFoxuIXuDWTk6KjWg8F7dNL9UiIpxE
qMd+RKBPZ0DqUIA8bk/AnZSRVW/+Z9sbmtvmy0sTUSKby3drS1dI+7oaqGLeIfJgryCW2OHoxn4A
EnDvJZvuue5f+vMn80DQLH3PkURIc27DsIPINmk+1Ds/MVbpkzPiFdPIGTQ4ojzfbNYNUJenq9SA
g0OQddXS4CbooH0Mz271fwjh7WxQpMTVwBAWP52jGhLSBwqh73oWhkq0qIk7oUNSpA8A018dVHd0
vC8o9QigLr9e2z2UHJexYo6SXxk2Cbu6vzFcoMf2SeQJ6HZASZZLVW1TbGJBbpRekNAPn0Yjg24l
ANXIk+NFu2oEYkAOvtVfHC0GHyrD63NFtWLO/mOryVEWR/QoXmlAaYJX0xXcwIvKdzOXK/3etzzY
+JQxIwBIZygxdqnuuOEED640K579Lr3FXK+KMfM6zLfhV8kylACCDIGy5rm9eR+gwpGCNcYmf3gU
6Uusm3cT5A1v1elI4LvA+jkF8e7Fxh+igtWv2T4AFObxZuiEiMxPucTvkjdHw/bIDAIGtC6AlKKV
XXcQrlbUtuSdxjhtP3PJKvcbmTTEtbeMyQWmLJayLrqywMgq2XhjOCBsJTqQtcIvJsmYvS9oDyeQ
Y+kCtDqxaBlHHt+VkIOv/oUADugVP4TaKrZWzvSYCtXjaEIeJSCpVWlrToT7WwWKs8RiGHcrsOVi
+NXe2IQqrSYeMl5zD7mjt2uzU1x4hlfOoYO70uv9/EJoGox5Go37q3mYrVnsRqSJdg3st4pONhMF
bG/we9AnnXQnyr+wTW0EG8MQ4Vv5anCUxMEGOba1/Tdks4c9+hCEzAJod90A16Nm0lj4YptxPZt1
Wmv/B8bMsmGHmj+QzZqUlqGa4GpHEZA2R7zM8cUylZsDUKP6QuhsEkl/zIdWRsPCHXMS70uxIaF9
onwngX8oZNOdErIZMmYD4pSr53kY7QO3MtUDt7xIEljFHuSvVvauvMoFzHGQ0Vpwq3LnLTFiyhCF
wUWmMYE4Z7hzQmniMZSJYSMYaw+Nir0klQourgujlC9pPTV3ars6f3BeXNMscnnXj7MB579Zugp1
K9AVDygBb8PeZO2tZ9bblf9tpw6EN5OBXYKnnwc85Bs/WPhHiLXeJSCyPsb1sSCrPLSir7cmVi75
q9HgPJ9gexcvEAqtXZFTr7eWk6sXUbLzsxV7GCHZGpPF7LtAwc5LhvknUgfKcgBjJQpBrhusn47L
ZyJYxJiZOFjVOAVZurFcdQkI37oSXoow764p1w0rBhXnedKoVC/t7kvDzb46k7HyYTRlDFvoQwKh
BcF91MkNB9gR/G6ZfyVEVS5O2rmv78uhglh4uNCd14/BsJiwgFpDyDcahgZcdV0jU7jrTkegyYWV
k5BSiD4qggJQuXCW8nvWYFbIjgmP2+cyKNYUOxKT0dmcOAA1TC6QM6eTOrTPW6HWjDiUv8pbZK2p
2xPhtNPUYcoyf56iBCtCY+WRrvCOpxBuj3PRao3xgsPuCpXfetKpnSDVJeNmeXt4kVWEys7Ta0to
BsiWxReGVE31mkrR9k+RVMWM2bRtMCK2x7GfC3869fNuEOmMLnEfjpk6vdk9XOT0bHSXCKe94dEq
RjMJDrieWFfwdFIphQu+zoDjLJso8iECIyjUozLSjrPhSIfuHFV+9a0Wyb6YOIk+WO65OTRTKTX9
21YnkPFSE/OLIOFb/OjWdCXMYptgasP8yk4sQ6xOEVA95bsga2UPiv6N26larQ8wn4+fiXUoIa2+
ovd+yOMTPmp/C+W+reAm9XzvIJFPZJfMkJnUFXKQYwIItYONZ4OHaAWxAL6DEqsJe1DwaCMlF2FN
6nw7SF+9hrQ/yQjPWSFm8ze4jboTYTGU46JBpwYSSyTGpgkMEDPaw7nMj6xDL3DYHdllMQk3Vzj4
z8j7QDxBB254Dyh+l9fMCWSVk7PlwZF6kBL1IN6Nalnyd/HH6mxp/Ow20wZVGWEsXZJnQAHw+CF+
FEj9z++D5sygO+vMoH4anbF8X2adfb+zMFW04qpYkgaMD0GkS9ReWiwbmhzhvIkLp4BfqvUKDC0w
DCeZcyec1xjswg9m0hJne5tE704qdcFlCrGV85s/IMZiHAUHZGAdC9vgxaMKi2T+6MBelOodo89g
BUuh4TdMmSM6MYDc1ccbzg3hkUUHfwwCrriPhzITRh6ajM5xHOtSxLkfFRhoWpOIJbWeIpb5Q8Pu
RdxxeNpnOsHegYUzWXRn0zt9LVyjFl2hAXWS7su5Hu5EP9un4dZ1qPrN8k9gvrb+ZaSI49rdqbqf
pPhSPCEBITRTpa2odxtLfA0fDOAUvUYadvIJca2OpnsqhJJDwnbD+xq600kXkpOKtZz+c6DtmnY4
wzD2xTw/v137vAg0APL3S6nvoakkY8c1HbvScf06SiZhj8559xtBAnnbUUX56g1kLbjJg+uMCrTZ
umUzmYcHI33mAtUX0X9U2gTcfAveUnzOD519JXS/n8kLCc6+AyPK6fCoImLhJ0aLYykhfp72ECV0
gw5yYEWO9LokcSw5C1466Xf6QCbHe5pn2uc9LBBROUmoT+RgAeciQ5S6BM9cFLwXy9o8IkjKL6vx
ChJ5JyHwj+l8xbIdZYrxZm0TiFlSz02CYAnVhREZ+Izg9l8ASXmkIeLL4j1W/sLoSFcL95/UJFG7
uY928wcpDN5ZQUGxpA2Y4QMxBDOl10/iqqLsr7U1pAoMTAumf3CBVJsXHNX8bxTxShiwIZQBj2IW
jgNEXjfa+LBnaSdfZiUY1/CzPXU8TAgCVV3uoMGbG577ySnClw+HVV0iVnvhlJIur7GgMsMaQ0X+
haPbLwQwaDsFCgnNZKv8dzGv46nVhDIRz11z/ub8YzE96q9P6GcWxcDkDnoO/WDF4mQ5XA7Ax8Qr
6YrXF9u9ns+5ycfwxKFIdr7SYdfrsjBAW6N/sst3MIUYYzVnhHEZTQw/+/c7pxqLN0yQc+j9etVf
Wx/8iMHsP5klO4VvyjtRZlUM4WRPl8KMV6Z2nYzJMWYj1xWGy8EcntHgZHXXCnPoEfdv7l5CL7ry
GVtYvwJgmhzmdDgg+oh/gfNu7lcI5tIygZUq2NDafjuXNiGD/c7op3Y3jXIlqrSG+Xy78EC5uJlF
M7CQEef5AXwRQnViTdfsF7AiLPiygx94c0pBfhWnqtQ1CjIOzuAEhmIbT4st7hmpzN8XS6x7Imsy
AeTGmbyf7LsSfwF0hcTcZQGZy9K2moJB00MHT54/e+N5oGctfcqyhXpq0FSnHVBsD1FUUoqfGD36
gazVYT8zrLAx14MIjkTfumWYMjA0H9Sh/LEVDPnU9v5OeW1mUo5BRTWKTyPV6MzZ2WwtmEBoAhG/
3PmkpMPhumrchzECcOp0MV52NB6ipYQVuKWJWcW6SKwsLUknmwBXvgj5KemeoBq0swvKwkZssypY
SFgsaMnRqGKttHt/dw2LCIDp6wI+FpRbnpSC03f9EERe9SWvvgMq0TnHeJsJYj+PBW2bvLi4ViFa
Leq6cCZarXWhp73wxf43WCgmzzNr9mJwcNjZCqtAORjQB2e6Q7fNLFgWfL3OwaFFQTnGiDpanhuY
rd/TSR/J2MyUG/r+kewsqFwTsVE9m6K02RK6G5gm8U97RHT47UqG8YHQF4Or2vNyD4C94EjI8g4m
y4CSpnxHd8olcjY4W0Mw8vQgRjnWFU4O1qbkjJY/7D2uWwqWjEtBzYk2RTsQ1RxI0cONzHGJbO9o
klK7olS9BOw12gtWqJ7JndWOFI4CTs5+oMO6TsMgVU//JhqRe8kvNW9Vbe4xUJDQeFNBUZlhm0pB
gsnGzaJ9dgQJX6lw3+H7Ws/0OyIodTYTHeOAtQO8UPAr8r5zGuVcWo1Ohp4ErX3gFr7BStiP1Rem
Tvm5WFqyNVlV3KY97q2KLZhhzPSAIybIfb2jn5JF4cTmry27oMFMmLW66YTZPQfAxvqs3u4ZVcOH
K6poa3Ixc39xtm/oqQrln+Jbrx7CPS2IqUSBXZg2v8qY9h0z5LLUq+Xrvw73l4RSA4ZbHkCPdeDV
bf5gtlQuQhU56rvONOhurTeIFrOwEcu94NBeHCnPzegM7VJonsfsHTMDJ04mFQPQpALojP+5Gzmc
OWqGdeeHUvOkHcE7lX35LJ9Wjjkh35kt2vdq87LAB8o0wu5eVOqX9PQY9w6eXvktcs4RnHFZmtkz
iRhvx0pX9w57HBR7gtv94cmyAfW6dBsjfHKC7BmESiNtbWKCkQNg9eaBTeTVITMLOLZj3V0eYC6X
UDJ/YhO5IbsVaizuACdfcBfHfLGpwcF0JPOYOUDqeC1bVSNCY+YSka1/YD41TsMsHJ/TVS6b8fi8
tOJkPgGqDQJloCGclDhfRD1GHIvAcTxJJu4fwkYxyRVpvr5G+qBPWfcTE7jvX7wS1+vGAQKsDNTy
ruiRO3LHhE8+VeB99bMh22pocPiPUvcm8AYw5qhA4b0ecc48MR0RhzraAzNHTfF7Q7IXxAzO/ylu
GRaIOP3JsUz1GfP4YZa1UpDwd0VM4wJCOSBS4kRmtGM3CZvC8EG4wAPXfViljzc0x+YB5bkRUU6k
wr5qgw3LgU9LMMHDXMjp01bHv2PSgOWv0yyjlymbFJleKB+PRV0CjJz6rmTnl7qRVSPWV/ukcsCh
hRa1e3Qm2N8agDbBa3EG/05hToBpkqK9zX2iThPbHW5ei6vOmm35zlS4aCjklqpQEpKXO906OMNm
1S8WWcYFhMYVJ2ELHHRr0yvSDMpG8UO9NR4399IPkExUN9nUf9a6j1g9RIyZ/BZYGv20kMRhYxqk
a6A1KCqFjVy+S7S9TVO6igC58qAPs0o+Y35/U+JWchVM9zt/5q1rdWh+tihn7a5zeh6Kt8OTMlRY
ujnNmmWYfi0MQF6tyrZv67Z4hNuzH6juV7Z9htftLYYYVYuVU38/OAWMf4yt8VAemCXrrCL7CRPp
hokjf5FckBey3BeZiWGZkeKfp9efXfhrz+3bhyudf5HmQAWmDC7TJogEms2jOLXKV7ZeX0x51ZqC
FhoLJh2sQaYGBpNsXdAqyQN4KZtRTsm+9Cu6f+GTDchDVcQXOJ50ovJo4OBNN9JRVjDwoOlimRy1
exvxTc8Ohmkunx/lwg5zcnglquoesa2R9ovRDrfN6c0yE5QVVuFvFnzyVwVwcSpUnxB9OMU+x99G
4wf6j5v+YHc/K7Sx+yDaqindoW2SLOcxj0fx8VBxdujk6broitSghSIC0WSlcBLEUMzeeLjr+gUf
CumYgq4U6LANQYRBV3JnCpYv0XLBGbkQBMntGTrvaz3H/M/ulxP1GBzkuv3sD/Eonc3yW6mKLIVb
piZCjdgn6EMX8NmFEZ4kD70m699bMX+g4vMaKqa75/oI/yx/4GV9hMowulMfSwM5RjYa/KoqNBlR
e0Bji4WMbY8Yf0+o5mpzB4xN6dbTBQ5vM9khdtiT7gj/tO9lKqhj1ylDf09I2pSuKd0rjcGgKwS9
cbWwm8hPDqkJEo4iS/s/sN6RW6TPwLkA6PFHhSiLQRSFl0lCGt4Zq4iypkKxvNU8r7haIP7S+nKR
f4/eDaDo+6DjM/X2m/+VJiSqZfGHWbmG7DlrTEVMnb+8a9qs9I4tFtgwz37nt6i4Pn8YNq/HeSZd
hlQvqR1hqZBYxSzxGKq/OvVw1NEJBC8aDOurcTfH2D+VJ03N2q/Nt6GxPxidKygYoMXj5d4jvXCF
MBLfxf5Hz0cfvWukI0fUHZ2PIskkB7P/fbgY6dmGAneB8V+deDRNcVMYvTq0DmbyOr5z8ZjzQ4fm
l0nnBORiJFJ40uiT2VF4Prou66WZsmJ0bhSaChQXQ4Cwi7cIgozNaovZxU7rAqI9nU4whkrLhiHm
UBBuMidjMBygaLknhBO+Eaqwbjje8HRO5EaiyZ1PkkwEXpoQRMvnLSXaFWHEn4Ko3wlaxb696Nma
Bi+Whm2y6I0bqQ5CgdcK0sh+Bu453vxdOcF0igNQZ7ySxgEzAnsL2qpHQXlGfkeaOEHspgf48MQV
gcXAx2hw0e6ejD2Pqo2cNyK5r+p7NRhnyt3dPxCIn3sj4KMnnO9s6gbpEwyNYaaB7bhVwc/lUKzt
vD/pwq8DzCU0qlerS+MeIArCMQqUPxp8AM8jwWOlRRZiFMLWJP/DLofRtsG7mHX1vbemhWmxF/C8
5BEWCd6PvizjJE0ltSKj79CF5hH2WHghamaA3lm0Dd2gf159oqPpQWzR6iWeN9w1hcHc/cKA3/D1
azq9FmrKDkWEZAslaNXbh0YkiZQmSvbpiKqdwdWJAH5aMG8ceexTYBuKYyUOwRtBmK3E33ciOeY5
TLHNuLK33fSbgar+6HnkpdTPW5Wlq9roLjHoGyou3y75a66Q1QhkaBJeiydZyFT2VYd2N4iCM0KS
aSqUe3kr+3QDeVFQjwjjEfVpZL6IIxw0X42o853CfVXlK/clKu1W5trlcTkciN2Z/++ZGdvAITik
JG8WcbdB8hwdGZVBSbzdywYz7uPMTSmQZRcGJm1pply2I+hoESKiizyPlq2T5J8KxtqJ9M1UvlQd
QU3UXMpihnP047Gzcfh4OuOnvGtf8t5+af1IjQPImMqr5QHgQyLxH+dQs3D6uNim0RUFH+53ESX7
59vgdaOHN2BPzOxXjy8C216wwcge82O/uzgJUD0du0oWYNhQKpr9HxnbrYqCjLL7UiPBCy+Pc10T
muWgAyDMcen7ILICP1vj90P+enMeuBkTInyHuYVLNRcjierwILbG619MNLFcsqEDgMqtianOY4rD
+RB9Q+Ke7YvJ9PqnMshdg0n88DU/XHSfdrg31uaO+eRvyc2+HfUQ5A/FYdza65lOoI6rpACKlKfG
U22ik/a5j9XwyCx3gM2ygaX2cvaf+EAbB+PSUSzMV8T4H5gIHqKGvkv35BClVf84/1do2kegEe9N
uT5qTugQ5K59iGtmM7vxGmeDkTX/CpDSP4A6zDYvMd7gFZJCKJeLf3ZOog0lCVE6ZvUYEnyTVVkY
J52FQdJyHY7SsGxz6XIYfLTuc1RykUJGVrhtoEb6HjqQJhQFerJ6TXZgLQNBJIk7k7Ir1EQLFps2
WlZi/6BfsmqXRGzhXeJZE1fnYqILt4B5hZ7fXJkCtwptkP5YZ3jl/tPfhJeQVtPWjSs0XjWDTs9o
PRH4ZZk0huxEolzYGu8oJywpyWMLZhoXIFuu/jTQly3Ou9wXiYpp36v/XnkdbL5EUPwHquSpuUfw
eh3jAQwV5NJAg6cPRVlQRGkj3vJSdIm4lmeoRX+j0cgHeOAEG2BeDnN9kxFzbdioNPgSVWpE7B0B
e8hwVye+OGZZeQgpiQaptwXSSLFVaY1xv9HE3YjXuZGiYR5nmA1X7DYjHG9vI7jXJE7dI59fthzh
tWcXrHTJaXOE2CuXiGoAf0t3GAH8zg+eH49K7FdCSlPNyMJRwm3lXWmddQF7mRds9pCYcJckMOdj
2XhxHG9K9fQ10KIl6mTFjtQZ9UYpBtA3wtcf5hu6mNiMIa6jEU/nqI8nqiqYPWlctqPbqUhCk8fr
eaCug8HW/LeJnJBguR3x5u+6iIaH0CCtF5ctLavwZg93YhIxclJFAqUv8YxN17xzPuTXd76ZMUyQ
qO7IYhvJax8JvN6gbw0/bLFGTgOH1NhhDGZYYBXdTFwvpTTnqLUWOqmSgBlMQXmK0UQELQ5wJWkO
TLGiV4nmW1/eJya5EjJ1Q6Cj3WMpuDGIICp8ODPCGXPuW/LJeL5+nfyu9nMKhjbZU0gwN0JmdeLj
O0bdXZne9Xmxrz/BNb2p9bzfqbZGkJL118CZ+Hmipk0zNz09Td38iEp85QIdhLjYii3uGeu/Yr+d
znxbnX/0eg4uX/X+FWpc6/2Du2vy1X3hwzoKET7hwmdV2E6PXe+A6MIKw3rbr/azAqImnNnX2wrI
12QY1D1/Zmn0KFl+ELvrTAnibZITCMeB8GM0xqGjX6Us67fAPuPMsnniukxtvlc2S0vF+p19XNzx
HX1FalTfylBKlqm8JGy8osu71/phN6WEZFEwW444mLRbLWhoU58T66SCivw14/+28LgFh/7u7lLw
vE3qj5KomlTOb5yafBEO9OubJNYUBIlb+NgRti9HoOVHEiohUybTRRMccTQGrMg4Hz+TwVXmZpKU
YyrXG8Ke2YLtDCIsmYmSWUnRsBJwpk5YaREHcH3syiGvD+eXPjeaghcbsUIjRUuHA4PoPIKq/0tk
DRXk/hxujPRX7NfsZSRH5tkYJCjQQSOhTMBMYqwCDavYme5hZddr6spIE+/M5BzJUun6BuGufiRF
aICgvpt4TdbzzB1RsyBzGWIT1OBB6bSgJjtvlmc7/DhoA3HNoNAKCwdZ60cPAo3C0BW3/xrct1ZN
oqx9VdW6Pk4IbbrvpWWN8NSyrk0UrvBd+yCwsvwU1x1YTMi2Jg4C+CxS4Td0dcGMR0V5RLRaggg0
Pb+DMpAT4YO6SZQIDQ/WFUpSlgtL0cvgeu4d1x+KKs1ZfjGk6nVNJJtSVeYGuycljbu9+C1r0ef9
YB50FOb/hGzENp/gRSmwuT56P9CfvhKo3jfAS3BYSgMyNXzogwCc8jJgYcI8y55vZFXxAs82fRhp
ptL59/hnxAHG0qIqBoIaUd/e5BiYbFoieFKhuzRJoSXY4J+UyEuflyAQ0nJJ20Nrwxlql/LQ85db
aW+EeOEWnsNYLmrdEoZwzWeDFhG4IM8lZN0+0Smvm7IixdxLecjvEa33wANG93ea+kjGziTNel+o
XKOpDBRXffWcoOmkdRFmlsmHGo4MVYM4A685aryJZ3rMYuJfYX69IEPe0VpvUrIjQXldoDR1e48P
EtH3WsZXUlpO5LpEnVhsJ6IPuQnQXX3uBUJqvPYHg/9mpH33B2Ihk2wMugi1+kKijl/qyumVQ4hd
EU595SDK04n7yMy++4x5KT0UlbcFWdAsKOIw0yBRyauHDT5s6yp6LOtpnmNvjrDDbr5IGR09gsEz
mxx9bN26R053rVHdX8xgufphx+5RY0iCgLQOsXZZJu4FLOEnl2pOAfRJlFNgsQ2ZemtY8Tm4LWPk
0DThmphEuNK6sgPDe7+OMaO9JUrfNYWfg7GuZQKqIvQq8LAaxk5SlHZSyZLoXVJw/QkZyj/DXCz0
XPdtHiF3Skci6uKjkniJS8I/askgTSzCvmCNDzv8MtH/cRSwIdjZscvTuFElLkPK9Swrj3t6XYrI
cf1OUAu/9h87/+w8cR9U+jPVKhXW0nFDcLKhS0AzDVrdGsglrcZRRr3MbzDM3ai9KyruynuHClja
2z1kxrXmpQ4Q7e/8hp4JBgzG2fPPENKO1kI4nEHNa+ndBkjm4qJyYynKgV09Di5qUhRvYhtg+scq
mIyyp/uPgM4844kwpKTbaiEDUU0ZYWwuvgxYIIIDneOT4nfuW4uBrlATfXYj8flQShIgLKvUlnj3
G1aq7zHQtJVE8Kwpuk6FmMDVdprpEjF6AdSiThdA+3UOm8qbTD0bMr1zE/gyVEdaIfRSUJYLlQkr
M4oIhOFUycUhTtYUvIR4exJJk920hXU8pOGLea2M2WHI4pXRXIlZA7jgSvkF63vrgFCsogpSWxRQ
2WoTVoXgaftPJlP7JHyBgrW/ZBabd1J32sex9mEVsEPCpGtsdWQ9iL2jle7NSGZ8RfDU8orXHyzF
Odz7djSsBsOXsiRY8AuRnqs84F2oKiHeVGCzHQE1/6mkxvGfJbcivKe0Cyo/p41F4z96uJ2ZO1uM
OO+PUeIKpS9ryJAbEiECrXz7dAKd4L17RmkVtB0FG6SDAh7tP59SrBaZrDQGzrn1OwtsFPWHwjxB
GvI+UtIFhHNIuvqUCpfLi4gPN64ivv8Cwy4f1EsE79xtiG43KThgBaYxltuaMLCgoxPS9sPlBFoa
A3xhbYxb5Cqwjd+u29jnRhSF7+CrVJzNrisw2RraI1io3mbRkYQniraPCYKZ0Fn0qMEWmqrC8wgB
wMrFFFuQgGkqPIPA0hb1ybfGpaQNxUo7194wxDXzWWBr5xz+65UUnWqmfAu1adEYxNZd4sQyLPCS
3QIogZXhCs3sWN7zjnq1P2KxTMZwKELmCtfXUFMcjeXrHtBd9Hrt719ZavqKHrcL13AgQTT9RKMY
Te+L5JeCSP2SRQXOBW1psq6z2RMmuZQtSacYhuUl91Ua9OzCUUeMciqTshT7Fae3LWsSc1qweUwc
PDiZ0qSj628o8dWUSD1fy8YieG9ZwK4K6Z7K9FzjxWctzQwm7E6ZVBxq0/Ei2/w4I9W2+iA+mpCK
dfVZsnMA9SfNVZIKNi50lZRZmRMor8r1Jz7VCqpmrYwV2C+so5ncsvqcdIikVs8aqLQKgZElxNje
n8uQLZbl6U2Paaw1Xa/cqbPFNBHQusZx6UZe2gxR8TvPdCzQpjmrkwqnTkSCeyA8P+GlpEglyA2C
KYKPWIqMI2e9bHs+DdIVOQnwg5QlT4KjKRRDv1ODLsR1y/I1ARKm+Xg+OhySNtqSnijTiebjBPAg
1Uvl/276OQP9uu/xJRBrJUewppLwj5NASH1eB23CxYTtHSV/gOt1uUsxLM3ZVLiUcLDgoYuuz+9h
pPQTq1ds+og/G6GV/wUUEqRCjghGQvjy1uru6+UqZ5VfzVLa3domfzj9elfrewRXA36hTZdUAd/q
H9lwQ1UdjV1DY9d/l11ovpaxv0UqT1nf2GKthRETnW5RsFJ+kF9LrCurwurMKrAXOInFlx7IxaPC
W8GMXwZJ3PgaL+jTv0n+9jC6qmNMOVAgCNx8r8S5Qf5Tx2xFNbduFXVYo9zzhS4I3jtzU0Jsmioz
4Aqk5FlS+HxuNIxU4dk+jt4zCiZkhQUFL+o1qjVMiA3VX8HPqnexqO6rceIs2IWitNYVAWJSn/nG
jxzmJCI2GPJD4exuCWWqKHNUWDb8C1bZl2DszyD9TA1avG/y6WeyvXZSesUcVBWgjPo6a8a6cSJZ
0dAvZuqJmUUQ1yu/9DU4Jm40hw7IHZluUUiXj9zua6zAvGchsIu8vEynwVaM1YRd9TX9ZpAL7QYM
hcvf2MIYxBmq3d/VCtccNTwY2aLhHeDq204w5TUFn4t/riAOovQm6Cq9yvYJ++Gu07OL1xpDzNE1
wOYmLSl1YH6tbjkwtLf7iX75nuYvc9rnLwGdcCLEU8JHhfeHk/nC1NdOK06IoxwO+IHPEdCzSntQ
3LM45htLytjMZsi3M1D5UumSRscOe3uhBGrK4P59d45fmDLbqzIo/dblT4lwK3TKyYQX7JPDS1Xk
9q2Bp+3UPEioAMZrEPlRQbnC0QZqXrlPcIPJIZSb8zTy0rj42xh7Y2cST+To8i/GivyXdb4E8n0M
Nh13HCqLpskypCxbNuvxlt+E1pu/Y11VyP5jvVuBJ0VIPqZKmjZUCxLR/M2ucIs1nteKPt5aiyPW
Xn6fAMwvjobkokl0dCIGt4FqF2lzClds/ktkjbHmwcyJ1VsdFEeS0wkLkqyX8V+933MlbMvo6f5+
IDPaBWndPVUJdXa5ol0r2PU5I2lZ6NpE/VSP5FumtYejLZ7aN+Voa/n6FNqMko5MFD/dfEIA66ZO
m3MI+R1gELXK54jbrQCfaU4FYKagzYsEQMPKkBLpBZt2GQc2SbEBtRKTC9FPd2YEiD2yzeBHcHIM
qxLdd/ld3jSXDcfNXZMC+VjDWSJWl8Olv93TWJTOuXGD8mYXkMXfJyxIkbDEfBggpVW2zAS70zCx
VNkOzwDtXxc2zk3jb7XfBVjOjGbc0gxwv3Gj19ZkXk3vjj9ZjJqk1cvUKIFLSkTzV5PhQIGvK2b4
V1QducFMyXLJGcGQps1rM7NSJoUbSvf0Pl5KNBs3KIk6PModT3RriCF/S9JxYA1JzvrSOHQBm4BW
7wUk2FKGRrg3eKJuV3MQ+o00tY9ldpOT+AsQe0fFECs+iIusgrs2zVRS5Gj+PmEAhhjgP1WvLbGN
JaZnfL3RlJJvTinoS78hS8kM46dBF6MBSt3XYEMiAIcrGeFmHxZrCdV2IStZAUnkEH1dCPRXihqw
9e8N3bFONIu9Mr4INC1Jpd5AIgOLO2ta5l2qKFxd73UeB1BgYlV2D3/nDr7rzFC1YtK0K6vHCS3w
0vGK5Iuw1ljSfOFDjrco3RblzDJSvuH1qzngC6KpQvzJW9uEuToyvxBViF+P3YmChpcfo5UmDHwC
l8WP13SKYwPknuLsNAj7voK2N3lYUMMAUBSj5aRtFOjpV7yN/+vXtgJxi1Vv1hMf+31V10DDlnnj
QFnO9UJvRrNnglpOJeuRYL8YNQl8WpIzXa7yfco9Ys/2vecRX7rms+7qnGo5VhNYo6cYzD7dbe5K
5MrapkwFMiB309N6M+cd7FYHlZx7h7AAAzbJHF4eTua0Z8feZAPXn4aucYE2DOYS75xfuBi4eBGT
9nONowMJtddQW8JXg0zJx9ltvuFuT7wffXvKeAE6SncpsZMbBxzvRH0uDpWc4XAC3B5KzNUUF7R9
D9dEUN8APHalQY9H7+cn0NrAIKUCgj0g3QZdK6k/zTviM2rTphFgpoaWBl/Wlgjwwzjb8iKBMLKp
/1boXBs+8bz5UPxJqV6GLTv30Mf5BqbdAboGf8c1BqO7cq8itoOA3zuhYm/oDCeRsgGkJHXhd9YU
ZWPQc+Czn+vdNWpzsTlR9AwkcpSZQEzD6EGZD7sTBQD2uvoYPVKlrruxba0V9jefasEuQYFIhh55
l+cpTL/pzIDVIMBsX3hB2yj3npi76WOyGcbt5edjNqrLj8ZQgmkZLlqkQQ5ilRys1lAMCjeumTiq
etg4dQzZg86uqYeqENmShfX5nZeboKHwKRaYtYEKXLnnfnPv/GUribX0PjIFpTBGF/dVl/fUj5J5
IzNGORXV9nSW040gQWBwL9YKrsQ04Eu1XNYQ4nhCs+E1e7AOG9tegX5F7Mz2/i95NwP0iAZ4R7kZ
sEpJklCNYYXZ0nJJJCR2zMbVYIjAMb7ZoK1BG7686lAPVbn6dddRgNY1XakM4gak3vXhdiGT4MQm
ZbOhOYX2JrGd9g/cUXxlhQbBugDJwIzxC5D90nC+cojbZSZlvEydGdI5oh4c6MOOKBpiYHtVG94R
tzIr6+iKeMedjyM9k9PAICw0T93L58zUJv8/bsTiJRsdGGubPHQjp5iFO22blMsZFl/aRpPbwZly
UnALuy5SXPViAN00/pWAwdzgogZfLGRnDYC+4SGAgSrb7FjUJk34vUWgXzSh8Xb/yQSQLaqO2+DE
AWs/bB8Fp1i/UMSb0n/UZCsfe26Vao8gBTJTKoxtu+hUb/pK9Lj7ey4o5NjvvaZqJAnIV2GFQ/9D
lSfXqzAd1ZVMhNhy5pOYYeVaLDK4WgpVhf6naGjk5I4DxtzTHb6pTg3ZTQRnsCXnX2e6Yq9v599G
Gbr9+gB1YHvp0w+dabSbgGRyFeuPARLGclHw82+Z/UfoLaN1U+T8Tw05N3LRncEPC3+Wv+dj5Ppa
WBdCKZdkWtowESjtlVnhLX+kZ7kdyKSLf++SVpm0H1NTKaG5POiC05pA7oZqBuThflPo11CzO0GP
lDpOZ+EEPxed3q42WTsucq7wBaz2buwv7OSzdLuVQxEvEgqxtuFvzzR9MZkNgHYJ3xHzfXIMknpr
mvtrdZM1NH5ib+h8OwfW0xeqsBLiokLlbLUy3/1NGGWrjrQeS/M2X0TJ6UzFTpHYZHYex7GXOcXG
3hlv7wanCuhzEvDte7hro7DVRN3l7VD5EpDqg9r/TKWas3VL1vhmAXjljtLRKKT2zyufIGjwf+Li
n3EfF7/7T3LpdYG6+XkTgwrGdNc3/Qy8eoHq2A4GRxXNqpdv70s4+wfctKt2dstpTmJFV77NMy8N
nPu7IGExQVPB2EMtFE7iFJ3jUYTjnTbwNNu3MzpBqlsfYRJGEtXxNwgYOT1IbFECYILrA6/ed6kL
4Op6vraI+4H72c2eNePsE/Q72eEHpKqP8pGHCsqoTJW1HTCepJgVvrO7lq91FcmqBvshHWMkWYYd
gOPBLGY5dtMHC10OtaZpPRKsi8qpoSB+EsO70DcIivr7D8adIZkw7zjlUr+NyifvsLp2mIIxXHpZ
/8g3RFFrSXFnCba3ZuclkYzu+TUF5KkYDmK7fecBDenZLfgw7pKUfuYMZtfvBs5GKehJaEdTBhY4
bc6pae0ZVRlcshQlC5pd9uCDw96D0wx7gbeV4Xy6aqCuY6o/0NbF0YI/jZmsqcT38kFoU1gf61ak
O4uu+HSKgPARxFlOuIfFr4S21KpYekTVk79mAsSMeZyQTf+l12HP7wFs41aGzwcJaFZIZ65KR+Q3
jnSqPkAAovrIHUMuWrs3OXeQMvgICyQLjocvPY6+3tlOUC8oD/GfWJ310U197RXdqfQdlKqhjKPn
HBup1UzkDEapgr2ttOUCOsYyX2zNR8BCJXxHx9SUTa4KE87pkkQ4R6sE5tDFJJiM1AdusMlZplNt
YvLFdpYd6LfSi/bKZ1dLs0nne/fcBkL+e9QEYhtn2YUohkaRNhoN2xd10mRs/pMMIIMHSDm9+okE
UvXR9pFF7HZuPgbQmeiF+3MKfAfjS65zbVkS/MTJyQAtbJOn0BLjObhul0a0GlAyLlzu7eNHxn7X
XSoZkebjTIQi/x7L78vFN6W5Pebg3SBHXzfyKogxV1vscr7QMdIEDYGWSQWU6TrGa0UI5X+yCpsv
7tjFuqg1UWndcsN/nvJgjGRMhj/Mk24JNuoRFW+neacvcsc7R3Qhh6zT3Yoo4iBNlwEJ3I/zkDpg
+/gM8uoQqcHOzh4frGy1o8+o/IXCqCzvU/b8BfEr86LG8KJuWNEvFoUxcHElOE8KKQhZgpv75lLs
Q2gxtlELh0GJHMtEQ8R2hBUpXaCQr9mOtefCFtIXzBoDE8QGyH1z+XhNkpWjFkDbQZIEoG6U+ePG
aYyyOdNOz1pm9zriKJxmx+f+MATrm/Ukx1vtd72BRD53ATLi+R2fq3iJc9HjccmKWAfA5t0M+zka
KpLzLrmLvgzslmiZbYCm0kOEPph4dsYz4E1U/YSmnZdDhH/w9d3wCHTobJC93OGjhXO6bzxKF9Dt
hqS00tkS7Z4Zpp1ZXKqRTCMYEdQLHqoOjDltd8cJ0zZvWThBlfH7rMlj/JHdH+3czIRojz4lyLY3
BwOoKDZOY6hetHF/UNQQPbqFiXfWU1TTUEfdyXVC6w1G09uR/Zx1S+xj+rnwvD6DVW65xZaVt4uo
36DRmzVGCu/WbvJD1DvL+eqSA7qUNWFSahTnqVPQAfCQ086k9qLVltZMkYPD+Q2wr5zSHQg+Iwyy
pFCCn+AgXgu7TD+Sl6MCZZ1X7QQ6eTmnR86abLNknSo905UoDBMICfa7tTbzWTO6lzKsLQlTeBZY
a7T6V/e7BGokiKulMQuv/dyZ5HN0QS9er/gE3UFs2WetSHpgqxK1S20bNIoWI8xiG3OIXQBLihQh
iq48elLVBDptliJM+acKs56dL22hGUtUAhdCNpF9h8CKTyn2pfc7/iMZxS+FcjSmBy2avh0LZiQo
DecaO1dxZ7Ed95DL7Zk1mowUoPU4l5vAOXTE9Lc6im0SkoGj1Z1xRlUF8zPKJ9hKNyahsOuet9mN
OsM2qwx8N92gh/juWIeb70OIhRNMtB9CYkLTjQMrQ9vNBOCMdxmDW6hQN3tOXNsUd9sT1HoK4Jc6
SmTc9GVQPhQFofjmRN6SE5xPcqrDyRUiLwJNffS/oX20waan4afuLtCaWE1NJKkeEQwDIcgtrfci
WiIGEsJfqq8XYmtze8jZhl1SOHNbhROyicBn+MWf9YigGhQ5nliDTTBp+UK/+j1HTGeylmD3hTAb
pN4e6urIXGftofomyaWraa6tXyy0njKrc+/wl+kajhLmGP6dqUvcquGsL1sFHLBonQHJyii8e7Xj
tbEHtoRb2qUlc/AkEszHp5h+1niEF2fgEvkjVl0EnzVAfZyfSTSmsat8bvpIM2+aZTjaw1Gvx1z1
/jGf2OPNZz6NZ2lCNWcL6AxHeJzFHBw5c+I8sVSrCZBnggO4EaX2225Xs+YEo1hW1aKNWgoj+gsS
UlBeT9J1fR/hfGChsvF/ApLoA+exNUj4XFCy4d2HM1UOHCiQr0A2TGRIjtw2zmKyqfOncDsWqX8D
ApWyN5ExzgsWMr+kWCO9EFbayum/Lw0mbItuoFmgcWqdTRBaLXWMjqIRpQmtfUIi1Y80KH73tmdZ
upbzESutyKCFjpSGW4CaO5dWquyOYWPKLSLjA+VhV/Hx5ALGa+3IrcjNzqjT4YxLR4TpOoDVNwfB
CYj43pqIH9aZUS4bpB6J91k37d3LdxJ/kTGX7qg97QNbEFyzSqRrrdUBcnKz6Ev+AyS9gBsovsdH
fKtx1evYgp4kcirGZqtYQhNuHP8fPKUn0ZwNbIPa8H3580mkoHDDG38RFyc81Je9nSdTdn1zCpsD
q2k3rGZVrHoHO36qALz8jLTDBlXrUGawtUJN+bM1bSIU9iNahbSYCq5e91rbwJhzTiaB8W6x+skW
FiM/fsA3W6+0pA6JX633ZeCBfzisemHB3G/Vljle5ODGATSvUqR8IycJKkfpPY/4O2w46NIElLBn
Kl/PyKChE+c/SEjpsnRCnxTDxuNYpIR6LN/rU9JZhU7+6AV82nRzwxbkmV0p4ngEiCRhwUZv/T55
h4P3rbAtAXVNo23qu7RH0Fb40Ag2XqpVWb0qW6qKZHoZ1w+DtYv7G/DeeGBQDw44plTjM562lt9/
ujIQRpS59HxaSosE8IESjHhfv6oG133l3P01t6vxYLPekvt7zaAguItlFVidH1TwGTsCvHZ78cOG
e2dXhJd2vAyBQNEIyjAQuYb+p2nreND+wziExHi0/2Kl8fAX+0ifsa4Nma653HeegARLxAjPIDK/
sEDFvhpFUNVFP3twlGyZ9OpXzZUGE37jEj7C0o/lKPJ8oQJjvoqazMrRZOfTGQCB/IkazLqJ9Yu6
8ZuqWi9TEy5O2+d6GIpsII7bL7S1FVI6F6NEQecibbR5I5IDtN7UxL2QZCzraIHw/Kl6l5Ix8c64
2FUSLeEQ/DfSzkpu2sN3seaG+XkLyWLMMs/kUAd7J7oR7n+nPV9PtsBa0iUSi8r8i4zFKXXUlVD8
pGv1QzMZcJLvxO3ALTe4SqwYaR5nQNTP5VLYc6lMavEOnenKCdpMLUOSRT59/0EHrDcN8tvH293J
/4REtsbiuD4oiVO8kIPnsi1iTGf09oEt1PO4uNqYZqVSNAO2tB3kWl67GrvzaBYKz5RjqEq0UN1X
8UJRbzwuhzItbCGR0PSShT20L3S9pIm3sYasripfjAw98qqFgNOD6Q4HXAnIBjz/HZCHiwD3QZ0B
GXgNma5rtXFLiwXPe7IHlwErKhJetdalTmMn+fGXh2v6zenHBwkgVsjnhCZ/72ul1n3FlE1b42/q
o52ohTduVyX8tFFnb00xEUKZd28j17zbHKo8AbJIsRzPfuF4Oa4ESiQkVq7j9XQbpL8SaZ1kYsZn
93w/e4pmbDtig5ywId2dZmn4HNzteoC+1qKVsmUBOr7VhvGPZ5nvto8h+zcChnyIR6+fDCXVWG+A
jUysOObUqvjwYlFn4XBOUTvea62vKmEgOLdg8cseJlcYSN/3ovwELSOwoXGx9VgMvH2bgzjQisiN
ninumz7EI0+uhF1JY9Bz3cVJd4zWAPdU/bew+dWAKHupT0TY2kuu1CQg0WBgubr3y4nBeFRkt1Qy
fPKisRYY2xbgvK3ob2f/GnvLJyhukeNaT+RKPDdHw/AryYtZX0pnzXcUqhFCgC4ArY+jkayiJ4vY
UHZeQLJr+mqS3j2WI+0b6S8w1B97+5bxk7cTFkHKExpIcMJZOi9bp0YoLcqf/KXVjRq4juJbMlIG
E2/zdhl7zJdOU8d3IQAy/nm+nZuTaMypausx8SAfOxb/AHqkvLdIrDBB9bA72exSXxE+fBNmtIIx
gIJt4sUe4/cEitDQidt0KZgHJgOzWalOKAX1MRaKKrrrgmKpy84CRIBryEZhIM19nnXYwec/2HdX
RmtTK15O7G21Lt8USq65tW/cnA5u7SnqJqvuJJCKn+Yk1wrO7K6iOYiVgF2z1N2xXNBg4+qiF2J0
f2TTOLmMXWijGnHGZjCn2U8UAlyczuZrXVPm7PkBckXIYLnDgvcsTZbyqfz8MOYs5/1YZaKBLHM2
3buc8w6JWQ8US8UnnAiso5hxhrq8KIWU+TyQfGlX4QZpo66RANBFWkiqHIsjEejsegYgtnK//9qs
8NDhCyw3/6NVaOxXMUW1fFg6WeKoaiOBUGrWrPrexTybNMkF941W8vyO67iTHsBmIMTs1KhwooZs
OMo7PXoi7zHE74ywlYdVjFF0Tz5KPggZ7amO+kLGp9Z4OpztyweDbiytTQNUDNw1NIcVowa65c02
DgBYZOL4omKdIU37rXuNVSC460Ez4lUmwN50EScYha8oNJrYSrQLkYNLG8p8iJP+YQoo0JwMsJS3
a6ncyJpHlyOan8TRAyfiWa8jSuikJWNZogViTPqG2B/0pbnXo/tvFNcaehnX4JMzaDDWrKtj812l
X4E5OaH8ZyUu7boATJTHFedi8nla13mSayo2dxSoIe8F57hqpl1DoBxNcAgSAO7TON3t61atc+EI
Afro69qYZmqMwBYZ5Wit2GtCZWGSwmp39zGj9oaK7ogW132Oq+bcNPKU6TYqrANgqQO4jpez/BmQ
T5ljyPaT2In0nqYIAYxqtw0yYmqmYFjxxHqwB+IWsFZ987Yk5h7wRM3J0tz/0rwsqw4Q9kX/8u59
phys/ONUUnz8AGW5VWmj1EzBUV2Lyb2MS6uxQa9dNQRkBYEOdbz6rbXbTdkA3igPnWKEJqsnrcvc
DRVSs0Mz1zhsQ9zmkCXF79bKJp4ewDOQ3+clJOMhuqKlGw0h4aHyQdWypMNUFqPN7TZrQVul+z7W
LveOVl2yBEmQd+wOqp8blCJYtStBNR0nLHTHFGwREFQo5OmGCHF/UZ9IxUKUrVEQLQE0t5EjWpUL
z4ZnF6ksN6Vt8ZzFQZCVD0qNttO7e/i4fhF3ddDB17SA55PT4RtSfAyV9aF2wW6YZ9OanME8kGUF
U3tH6vjw+snJmeEPBdXOtEKYcLQg535fX/BLr5wnFfU7JibadDZEuwM7LOL50kv69YY/yGLzyitX
Fdzy5JkbwW43Q3pTcnLF4kvD5gf4NAcqNAdGVtDuTUwEPRBdxp0vjn+ZKtwSwAJ73oyBybjSkcFT
fRXv1AVDgMxWmtGC0hc2BPsvnktDJ0MUjlUYVV4wAranJUO85NRrciKM2/hbzWGozUe36b+C5bMC
+mV7nLXXzXyzhej4K64zXj8xSUe3OmOE3SjpRzgi+hlHfWPWZez1ph8GIGjt+Wdi7YPhQr4nbU6M
r01+7B/mA4wJnJbZTazK2A+r32cqYuIh/oc39qR+VfVl7FnGYB/fkKfYTOas+/X+y/1QqH6K4BDS
LekmEbtTJG2Zn0E9TijGx9khVeUFVcoReUiRVXDeMwVQOn60hqp0D2+B1Sdiyspz7Sbd4S76ssSh
neM2AP8CeFdtXVEQGSMDuSoRyNgq29y6Uu1Iya7zCDCKtU7VdVuUKHR+wFMH/2Y43MR4yylOygg9
DdxqVFNE8dbDzA479R4UsCCuOxQ/jh0iyMcfu7J0pKyACbINzYdp13PMCsLzPc3nU9Jci3Rx4rRo
81GAF7QwLWnUZwDKr4iM/oJdf2l/LeHe8agExUSlin1vTRo2rKI/yokN0Pwt0UfL1/Hl+IGww1s7
SAcUqNfodBYeXsRLkV3F5X5MS3E2aMQzL4jWAZJxwO7NUvdRlUF9Qit8zzTs+8IDuEQIjQCir08G
+uLh/o/MdhqaybaEDDLA02kuZg/MEM0uLkGOYUWlSivGmMfKxbiACnnj9uIqKyGnIMErfPb8YKUi
tcOCY7G7lxkYMajQ8HvGFI73ex28e/AJqjRObswxZ4kK09/zMk6cpLs6+0dNuw4N8g1+Yo6KlpuE
LpY8ObR2ykWTv2FJjd0mMEYFZV97bbzni4zJn56dNsfZzcAtoyj9pbENzMQazgS5U+qJknMxTmvo
dB2vXVltRm2D4bPOZ24Yzet7mRSH5cVZB9pCrR00hExoujZ00yNIoF25VR8d7NNu1l3rzet9mRVn
/7bn5ixHUbbTGmWbvTYjDiLWvBYTFtSKiC2eOvDZ0hOGCChAqTFAwGNKgyZ4FmSLEJtBrNwJ/q/U
cjaGt6FKrqGWjSSSgdihjGPNX+2odN6oDBvmj+qz6zCXKEWFcH45F0MxbkgC5vI1RuY6lZn4Lx0c
hygeuLoV23W5KwaHPv8MfulBe75eu4Xwp/jRse9dmHuaH42G7TOzfluRLm3MjmavceH3HJHdXHQq
Rcn6T9m2sy1diHiXnrcP+3dbQuyjUgyLqs5d3pGgDRBTywo2za9EHn6zSwH2pn4OJQ+O8ZA78i07
etduofulPEITvzEJ8zFBuyAEHcV7oogCw1+gPej/H6DTqfGov8V5byXpH7CCWffJgNNvg5mPCq3k
g4U4qmcFyWpxoahXSXYh5WUDTDqku8w52dOY4MvZTJU8xw2mNCAKWaexZhtyjTae23TlbYtYy4nJ
PRSuOf5LmLNq6P8tpBfNbqEMdyYWt9W+s0XNAbYWkZHOwnzgrEVAg9uP2wl0aNMBCMpWo5vCXmbe
EqM9Q7/9GMsBEPsMhcQEXMzWXy6vxoIdSXbcLa97viflivhqf5g3dCQxcxLqQ8pjR5dPbwWiBgaE
WO6LcmO/bprsw4Nf9zakPnNxYu1Fo5tX9aIC/yFGXEOzoWf1LOw+AEiJg30c06RPaTwrtGoi7g3b
ZR1wsvKGFbBBs2w+QQs6iAuxScbzphRyvD99Ptmi3LM1nQ7OrvplVW5NS4naz6j0g/fX1Gq4DBdR
l9R+oUYi3TSiX08tMr7efPjc7c2F5osEabbRr/KOB2PNFUG6/ENhrASo+fakn49BvIKPvPqITdOR
go0/NsrgPHzqtIwRJpmG6G/OTASvBJMKW2hg5eVX9pY6u7oj8HzUL3tUV1srbT5JeV2EiyMLsv5p
k86S0KahpgI9wLDYg5FCtUpXj7lPBfGtg7Mx6Y7/8U9sVyy7PibCZtc7KQxYomTdkDLnpUM7cHjl
UkR+qh6Y6vV8fw2tPRP2a++xg65lKOB1q/O4/nrV/XikzNIHZXGMu3T+XNBGCDChGyPzXB27F1+A
TcX+axyz1u6xJGYERnSRkgQ11teEnvDDk1vxL95ROFCQWa3IRYtIDnAFGCSUeETE0CuXNDS/RZfb
6D04l/VeYsaq+7IdAijnckpVaOaRDkSLS6aGWeH374P7PNkLmKr/Rb7vg9eBpSBvXAkzApvKM0n6
KYQmGImno0NrVze4Ht0/52fLFAHqle1YBsSM+RU6yz9Cb93G18o/rW8aUYB9VsRPkF7Xe30ZsSHL
ppZzP1kUQrkjVCuUzdKSFQGs2ymilPja64l+yvw2K4lcRTKf/9GbISQoV+Eg25nRKgHfFnpvhL9h
dWSB2+v8UpAzWdWMTKxKpSL8k+cKpUbsjPiM2FZMCP+I9A2j0cm97RH2OjhB3lXUzbs3vf/RvTIG
fqE+UBvpqphLeedlxKVMcasRdBeNejV5/XjmGPHXr/3WTnthQz10gbFO9e2e4l5DvUm9NQPzM4Zo
xgWKUgMk/lmvcPeIW8DrwV7g2AwoAC5yed/CGQC/zdIDPixbMj//AEmNs2zZX1VxsSM9VYQGHKMx
tq4aoMovE9EMiy470MRTyJET/0ebpkcoh57lSKN05r3PaF+vV+kWjKuf8QiEvrs1EwseJCEWi5u9
cMm/P2G1DcMbD2E62UPn63CInTpapHLnF02iU8SQ9d3C4pYxnarzGY2P0iu49I735Ydzb8xrQWm3
1vcwuw2az1iDlV/HZUe7RN0QhrsRS9GqdVuHMemosw1zwudJFt/jG47n4nHf3+WSWZHgsST+6YBn
HTbN65ly2JyZRI/v4bN+I6rwUJTGMhC0xH+3ogDur9995mJ3U9IPskl6UJwaEOhXA3R+7Li+n+FF
HLTZ6+IBF8Efwzid34WRIRbD6oOctRt5o+oEbE+NhkUBJPe4KiSRK3iTIeJJm8RW86Ou+GkUYOD4
dHZS+oXQNfypeqm9OrjSCqo3AlAe9PQDAjcmyKklGAcKdUUp+yhmM+qjRMfF7DmFhK77YvJ0Modz
bvEO+ofricGKnrJWXRzhZn4ltU3X1Uhwr88cUjqzZFg+RGYmllCA6ifBxKgifhMG/TnAFdablS3B
FhqlSfi1pb9TFl+icrNq7tC3DZpJIvSuOXtG5RhJJklEhtDCq4ty9NJnI94IJGpovo4snM4E6PQp
nHkFg5QtjSB3qbwAqYiusysVSvBfs3XcsQ8GmML55t3yKaV7wn/lPN70lv58e0S+s4wcBNyDGmF3
X09SH9fxYmWp/DJumM54qWV1i5BQPTBayT/IXmC0IfJrLujv1Lzm9fYD9oFmlmHmgJ8TxpOeu5sN
PunV7rJJEt0Tc8PB3aVVgktHAU3BVYW4Bi5Upr7pO5Y9jAu27Ht/2cda4bH9LR9miipdocXbn4qT
KlQb3q2w1sN1I75Ci9kjIACabBhMROd/l7nt76ez6rfkjWS1JPaBwqdb4lUrreILFR3xakyBf+e3
ispbP7isE5FeMKmroWPRavqxLLZhsbtYusnGu56lBwzOSo2YhG/f0oRQeSTa+LxP3pY+XLVS/3r8
nTviTcVPDly4V9aOCexUOCdNWyal6CdHU9hkVXWYOef9jc5I5zSvXVCZyUNnz2PwcuHWmcM996y7
Hys3sboL3nTTmLeng5V3E3kNkwb0gfQjaGkfDLz8rrDlwmN5yeAtnQhzDN6OaLr+DGCyYhSV7rxj
WhSim9e5GH8bsZIxVJf60ZXLCac8C4BamedTvUJUFmZ5naJoTdmihZrx10P2YnP1WWj7TsAy74Vf
i6gNsn5vfSwC8uLGOmtWtosGLpExOPQjKRuI0DcVF8sO1I/3fQyxBb3Dx5s+jIYysksyX+ZIhFuY
hP0SLPdtGkNEzRNHhcoTW6hZIUe+o1Vy6IaN4JKif3sR9dfxC/7ppstZX1QKJg53NTzFWdTovtY7
Mzyjs0mlwl9VY4qbzxgAlK8TdXJ2FOR7puS0M2oTvctYDK50XoV4rEt1dsNXBnBJiq6LAVWCxny5
GS/kv+cfe89Y1vPQ9hZMFRZIe2CQlkIOIfdZctHOjFB+m8XwCzXXZUK8YmmHrQotvfkDnwIeBoTW
uDAPFGFmQ7H8fz73OcL6kLg/ndd/8HaRIWgw+JASIXg3SPo1nA/IsUkbNylVGR0MK+bKaq8QNg7d
Iw69NBrLBIcIK65rJRL/hpBAwDEukgJTpqB6/bO99kfMyn/Yb1So+18f54g4JSHg3qYkRzqyJ3Gn
qZPJoBtEmFq/keKE9HbKV0Pn+nPqM+HKmT0VkZ5zQ28aWBJE+5+ilUa/zv/uzR9GxWUR2ZxLEC2D
AmAeLK3lZF1WtrF4em55Skciaby5JsoH5vcbt+iM8K5kAkpDL166BSzceqs3ooQw2cIPlqhRNNOk
Kq6ru+dZIEmE1LymW0LekeuDeEjVEiBoAmqkyEg7jHhl6WanKClsuxqmnGbSx3BN6r+Ukxe8LKK7
WV6nTYbCNds97QMgAE8awW4vFsBIWOyJ0qujYom4/OLpkO17vEUE7zc62zUKJqNTDPfHyFcmTL4a
Mj11ZrZo9AcRjyGFZCJ9U/KIZvxA4SLQ4OVab5Yt15HE0YWu/3c6C4MIHe7MXXlqnEOiQCaad+4n
7U5apo3JTfm/kQgbemMilUrOI21Of1N/jP5JSIyl3XTgm4Z9THKdTLHJ/zG8QwFBkk8uCFYc/KAC
BTGnbsEn3jvNgYvxYr9eHI2PcgRy8DTvMWReCXIVRHJE2V2OOonZr6V0aSI6fgOp90J14Rnc2WgX
Aua1qSw3pmmHsCo85z5lyT4IOy8FJL9VokmymUVnpyhCPnabqCmRrmf/3hYpz1rVt1Tq4qrsbp2X
EnDooAcFAoucsln+a/8GDbwYzGYc4K7P5uT82COOdmrERJYM9JyPUX7TXP9L6aY29xUH2GcQOQN2
dZGESGIgqpzQ/VLLznD4VnLOfaNh9D5IEE1O9DEAfl30ZkV4VOsRpz2nqeXjC8PlQqr1cnGEaGUW
zK1GJC0coxBSg6Gp5bple4HxCzLG0N7P1/me8lLpZN4iLERVLIiEe1BPX8aK8uX/K2il8A1OSosy
RPMl3zaHGWHP/qm1lX6rPaVPpay4eE/g4XlkTKQjEZPzp512va8dXqWpDF5BbJZWtBiysJPEBlSg
yPa64fTFFv+PNzb5SgckprZlz8MnuInsqmtoMnFeWK0tUgObDOVxGtkIEuKfkRLrUxeOB6fRqzIH
aqTbl+IZ0T0nkRIfXniLNc6RQgWTICGEmSP64ZdpTij0hVOYgxhVSDQIvci1GUBOBNGcgq6qIpXF
Xr3X6CfIrZsIea/U7P8S2jVEeQy33MLTHG76uySa8fDFHS9ue0yBwkNBESjX643AMoPEXDr38v0O
Kwx3j6EOeKAekKRExqNSnhlqS+QDsIZROHVV2mChJDO+0hDh7ytT2+rASM3vc8AlTLerUVsviMgs
w5GVP8rrJsyJAnzXh716+DbFql/rYMzok0OBHNZXDpMRVf8ADfVJgiukqaOMZloP6tefyF4HqF+N
ANn/2PlUHk11N/1QUBBXUjVVYGthZ27I4Aypfds2bl1E3W3D9Z6yUFZFcuVHUytAfEIlLu702Gq+
XZkijMh9gHss0ArfPBh7mGkA/ZBLv+HpCqcQpbp/Ue9fq6koBptE1WI7K1pNr5Aa8rfe/QCF6W6v
WFQmtCL+fsan9L9GiSYe87D0hu1SA/3TOwIZk61QFoxpdUQ4hH/CuIiN1HwMNI5kxRl0jfp8leKH
6aW0PS8/4u7TR9XkLNmutBSFFJi1sVqqyvjE5ecg8lvdtRgPe4m07f4gRZLcjv8LIzv/IM/3lw0b
gN8/AOMGg0rV1Hdfn5xINumGr6Nc+OWQYXvjNyrRH5TOgUYIRoZW3syiBfObCH2+iGUrsMo96vMT
EOXFzK6q27mFjg9ZuhwZ6IMG7pJ0+p8Uf+vhC/l+RE2hJFKUu1w7UrLmmwOPehWjsszA8WT97Qe8
+Pw0jhZDh8ygxrVdXu0d1hbXWS1dq+3E/Ocf4C8I5bhFYfSz1s358NerJmkZGUylVynK6V7ZGS5i
ip221T4b0xwXRmYGX2Mn7H6D0eAeavLkBvtQRpYZKIbcwlE1doQOxTkvubjsX0cfVYp1cbhT3pLG
J0eghxq88275r9tJuAs9hIwhNreu2GWD6fgJ37hBVGkNlvnnyC+lLi9uVSSoiFJefVozA9cj9QZh
shJr9rgIoq3GOBoht2vX4eNhyHE2b0948Jbj7r0Xw4PAwObrz/0zB/lMjVpZ2u8GwxnOGn/o2KpX
FNCacyWs5uEz96fKj7Y7gl6E/3grXLNzHvNWIYCXXDtCiRLJ4OH+Pt6gaZYnmw+m6XXTGbGwNQ+Q
vtd++j4dXHDnJItHlYZdHxCV6qi2Cva43mZxmq+mOjSH+ehQ1Y0M4OGrjD6XgEvNjKn/xfXetLbw
/zF86mMPHcSHgYhrwr8Z/yRyf9qFfDqNHrL0B4o4/k14Aw6jhy9MXbqb2j79O15A/PCCKtSLFm14
6gQfjMoMnzNVN69nSrffsdu1YcOJX/cmUCqxm9vNzRmXyL5EahF9aP6ZoIRirN04jrllqwhSWJCO
d/ZZLjuBz1yhGZYvEryjuvo8OhoyG9DikkgvadYtaeYPQRy12U2dPkuznyB69ilLATW7VBprpXLo
9veIhptDI/4VqR+34zbrlJumtNc8A9xEOk39tHG3O2ko0C295qk0rmgAqcUNviZXrUYJDZ/N7eYM
mEv/GuAmvkIoAW7fEfhZMET/24zywMExdiuKMQt1Sn/MVsOyB1kcdrHFxrsR/No+3VAiiQK9+y8L
sBg8hCqt4GqiXC9ePzF48G321Q8c6gfqMlZel9wVuSHS6vWjCsypnhkrSgCNGXEI3LysQTgBfBgE
eEzD2ft6JRcArtVytxavLVc/k+GaRDyXZenGEOPVn85f5OsVz12H/MHSr+RgX6W46Jt1yyfLrVzz
3UWaTCE47kf3Uch/OrTll8nY5WggEeJjVTHJYepNaOU9bsG3HROsARLNej/e3eCUJvSXThtJY/7W
LeSNZDc4Y1ts4ZoJk57xs9ClzYcM0SQL87Hv3/cNhuaeXkcCIS5LEXdUiMj6Zc3oBWwgRYFPjpp7
6+7hCMp9jK+QN8aUkIZ0t0svLeog8H8VZOMYF7594oknyDmH/kulsAJ5Z4A2VwXBUnK0I8+mdxnV
cb7RXZ7N0IHV07Qm1Qov59D92VTD3IZHSZW1ueTa4eTykc8laGog1RuLKE6w6FDHou2pVurg9ZPb
qHZtzJsDtvN63sMr4PvWK7cLZfCde/YRs4ojtzpo1um7PKqHWN4AjIrUBchHk0jDfa+V6H6L2YJk
a+dfKXNq7CpNv1exUrfw8HXaiPRVEpGWLo++zONjo3Bd6kdgt8o69YdwHwt2x28epnevRimXRwE/
VnEQTsT4UmOp7P82Nzse11VePYuN6xvhEBhvVt74RGd98pK2aFLBinUPDjQA5ExgL7DELFD7S/qO
tUulVcDyljQog3cLl6qccmQ8LPIRIO13q8jJ8gjN+E4sGLht/QBGRALFnPBuebD6JpHXnea9tkIO
G+bELTllfkFKp08OFFdFrI4XNLQYyuH6aWTSG03rW3xe8keXL+hS8nPOeEyNeS1MF2S6+0eVLb3X
dhQU5FgTD5fevhm1CEWwU0LFU2fSQaX0eGemLWa7UXdMDH4MvfAeiqcImAWfZSENrr0lqwlpt3o9
xsGdyVFX6V8UQkO8yCc6yroCg8910r711QcuYm200r2T93vi+Yxgvof2FfXWMTeCvyyO4znae1pO
5m3vlMR+bzzzHo6kGHU43AwZehS2RxDH7EjZnMmPjN3dTecGZIOO09rINIwJ+9JIxqqly2846yCc
iAa/goc8CYuhPQWQDa+QAHyjqOQz1QvLjK6VIbzgkyxFTQYbkTIiLjB4yNahAsPnzS589s9S24Jg
Z2hPWqyttISf1/osFG9Q44uc5SKdKZTRwD5zX/yirWmszNUgQ5whdKnC0VjP8j/bef0P2jhTQzoE
/qX7uu7+vHatFji/gc6S7xiLaPVheimVhaEBcRGlbyjbDDQvnO2icWhVfz754x573/HbV+TffFSl
XpGhhmzxhwMOajz5ocMRxtHQoYUvhhfzjKwtDovI4l5K1oI5YBq20BSGTCaKuRz9hVf9ViYbjE9i
+7zSoJQguLNkDWzSWq7DZ41uyDCUb3WeB8oWar5PlYwHhajCQuIrRw5xv9phkdeJF/3Ij5bN+fVm
p3m58zpP3BYtetdW4GB1HVQUCmyiC/CDzajhILs/1qudDPcyCVc8xHdOG9ivD0dbXf32+/hJKA13
3F11O6jMeOqusPArVkhvfDrSe3n45BwQfZOOowfkGK8mhfhgtqDJxuix9ns0CvtnLToRIvnQLDmK
Cz2rTQEqPmTPgxiWFS2iDJBKXao3IsfGrXojtRSHRV1voFAQDEjUQ4JaLin4wuH+i7KkqBdwEH2h
p2rmxJXJmAQAs4kQWLVTibfSOSxOwh+Kx2FGfxwuwGEt6fLJfS9SFDw4eiDgKNlcw6iSWiPSalOF
UrfZIbUgMSss16o/g1LHlAYorEaf1LK4RfzjKZjPAjfldMOMPPIyHKV0aqN+Vscoj7c4J91FjpYW
D1n6erTZZG3BCB2i3hjGHXvNcRId9icsa7+sy0gIElh96gXs2FJOANNgsUF+6WPoU89Q/0QIfwB8
pO6D/h0q66UrPKZVaniHViSxEDTkzwj1CTyG/J3cHXSU62E8qy6vNIm+ugu/7L0XazBEih+XaNxQ
eweWfAfid8aSX/HihhdvEcPI8qAd2pl5rbLzNZ1yBwKb8RGNGCeepw105OEYCSASI6Capo5PMf1F
+geR7zeLkY+l/4ZhfnuCY5NYmISBkQniNdxrtdUo8L0da+9BiVzhWAyuNuMwoVFfcU3m4ITOHYcI
FRsafhyIRO/uHMzGji5EIka8aUQoF9pgHWG+5UQ5xA6Ajw+vs3R8iZSp2G0kIEg+03Gx9JMjwK3l
IEVwdktC4rnpouwoD/PeX8p4kz7FoxiomGAP9bdpwLLOY0TyzGIi1OrShxRNoFUW+8vJPkfphqkK
eywtaJ3tp2XCoVkdA0zsY4dCtn7+xWO16CB/0Nfwq099zyusL/lmbAkUx5QBe7SGpLQw1DEq1urJ
0S/RAAmNRMlbgocN6Q2kMy4aMmTH0LXURYS8sjCE1/6Dy68RAIrdR6FvgBJgffr4XjmvBFoGXJah
8o6s6c0uo/TJk/pMmljkQ6kbfTt/7tuOcsoXlKDhc1xK5ks2VkRprZvd4H0y1eqqpmFsMCuV8Dc4
9/hpk+bmo90FEcXjdv7Kx8yO1WqcxfHhR81Hm763Oadrnj4OW68GiuNSMZVWGSUf3kSPTq/erajj
pTxHk2tI+nOZ+enVVPaeOP2Fb7xRk1OLbtNaSTh4qjXEW8xLvCk/I/lAeE0uL5XLwz01r7EDqfr8
0djamQFq2EuwntU1upToCB7mOZrVfg+c+rlWTP+RerSWGqYenlOIHvlsywqsqfehEXQVOP8GZaJN
sqrTV0UCvsNfceT5ApXyxOZa/il81aszEr/7EMx+xaQ3nsObthYumwhiY1hPVLX6EjSN+OFHBumP
r9Il64PYFy/yvHvNjDHb3zzVLM1iUBio9Qz87D8RJa78uq0fea5EUnRRkp6M6PaYE59oz2hth+lw
lW1+7efuMTtjUuCyVSZDRlndfKvuMoE4z6wJ3S2msU9li1LbAMZbJm1utfLDGC1S4Yc3V/+nGibZ
hJ1yJuGtkuro1j5tVcq066H9/fxwjwmbY5XKhEJxjTV9eVcqtzTmmUkl+Q0m+zCq5spB7lVdN1vP
XS7EchhtVuUTC54+ykN+JgPGz2jwY9yxhcoceaGzUgyRYSxh2VyokoFuFhBfekk3poHE0OKptCBz
Dq8n+N4oA0BI7JsdJs4lVz1NbOFyiVfGDHDwcN2zUpVxEP9/bbmmmY/Gm7ZcvVstkIFyf/i8TR94
sHRTrDIWPZIJ/E0Ni1A8UE3lTC5yFPDkIIW/sSSUbEqCkZ9AF5+ZHu1K04mDUlsJBn1T1bWYX24S
OZ0RA9FJmeExYt9ooeWwjx8t5K8NnMmidC9w2Ln2BgGHAwpIl2VG18x+PC0VYzZc6O6Lbx4KHWzE
P05RpaKtVH8l3bLUKIIY3d8F+dygApJx5APeqaxDw3sGablBYkauwBkiSB4mNiWkgw+rGOoYEYd5
Xqb5o21b0xiTdHBmb9FYemjt4hjqJHBEtqF8hdoJUx0dgxC/fyXrcvYhl4fOLrjGj+UgxGyZl8IX
reqNeMyaciCGpB8YooL5HVSVyrwVf3zr7vQQjfKZnp3wZhHuY0h6VtdRl8oyus4dSt4ns3G+Dkip
ggIb1h/Y1XlFfAw9NZcHfdNmGNesGj6exQ0Rdpiu1bLSLY+54eS9br3X5iewv1b/W6v+RpO5uMKj
0+0olFBjCMlg1EtXKN0tgG7Xq5Xsi+3WregJCg+a/kT7V2TUopjXwocwCjNBfyYjQv/l1ABFg6W7
orXfu0ocS/AbR4JT4JCM8hvT0zcxyQUCn+m5ghCAiufNXtgAlrMSv2lBtBaHAgSdgNVmASAXWgSR
e8JInIHVroxVWjvUQfa3vt2foCzjh19mFdnXQyExA2apX9NOWwnHEKasFUPuPqZqgimvY1jkd5Cy
WleTDx1Q5Lt/CmC/z5X45RfdMnkIsVWEU26RfQZj7dxGXA9ZKHDTVAmfzl0tzvsB9Ky/oo3fgrvN
9xRhy1UP+5EuzBtIiH4Gw4/AGShJDq/PfEPgFtbNyPMOMW6pufSRCn4UQ3RMYhL8YnUzc88456j7
C1mYKOu5G+02V0GZPFoVSBzueZN7M7Ak0kkkX4AfM5HH09DGu7MQzsx0a7AAxpLOKpINdedYIV3J
Idfg3l0ElUKBaeqw4sArVl3uAnMPdBlH0HVAdB/5Qza8HKEBxk6Lt5clUYIA84pEMB1iQFnfJvfV
bs+Uk5E5e9IWQQ2CG6DNb0Wdo8VeZjwlAcsHQFbvS+9rJLSCh3jB/1UkLYhhYpZvRFcR1vMq0KEg
THlKVVXfp1nTBhXM74UQrUXUQx4MOH4Fsjc3LXUE2tnIKw9LWu1TxWW7Nm9VZnXpEBdtv2iG0jrv
bAxNl8IimUoSxzmaQYD4kS0x+EXKHLiXX+466anFOlu9Qc+OMPRtfWtiHBxxvWhKNIYTKMcRbEDe
3FVP0zGRjICClfq2cyD2Lcptf2yA7xlKIbpPzcm6GuqM2ZaamMd6iqRd0dJacw93ObBILYnqvT5/
CGkpSOPoFluR3PFvdq3arJK5LS20HQ7Agi9oJBT/TR+9hFL1YeOyMDdhDZR7H4dcE/mhYkw975JV
RGlNqYMxSuCYvUarkRMDoTsN1fcW15BliwYyiJwmX4+BQ1AYqFYRV6YihEi53G3CQdEDl+NCgCA/
eegz/GA1aEfONPF7ClAMwN2QzVSgc+1PTBBTfYcANVmvNuckXik4JHYpsk0HaU7kKCqFlPyUATd1
WIuSexqE7C24zibkSKnmZj3H7e5Vp3G0iAi8webBfZGSqBEUqlMRHxuWGTblb5mX/0E0MbOKW3xO
VMfv109hD52TzZ9VC1eVP33bpMcyfi4ViSgEn/+nm5TvkJ1psVUAkeIlU/dYpyMTrZo3WudEFnL7
aSoXHPkrJUKy+sNWD+z2rPtJuv6xVPfmhAs4GTNacBkt/hpFnf+SnUe52CdJTm1iQbx0hOM1HrxM
LemvQbCstKfrZ0uYhlOMq/LAlFuRDbVlRvkno/hRVKaHQbPEkY1WkJ/I49kK2+CXBH7E2WebxMbI
T+D9G+B35Gg3bmizr/n44qFT1uILs78WV51Ln0VMirYCbhnalkwV0RpM1baUGtREOsdxjETdX3YM
D5xITaozcqVbKoFp+/tlXZlxuuM3I1ebBDJ5HXvnMzWPAyxdX2lWPB/5NcjTEn4BqW0XTt6Y24Eu
H7Cty5OR6KmaR20sd0qx+ZGXNqIy5/z3e8SCaNX+m/KiwSFLRdvM5XZCz5Mxho7f1oCnDQo5TJdb
vBKn66Abu2EDkAeQA7osrruLxTa8ZP5efomb/aLkGjC+5TI5uFIDtVeb55GixotRZ2BQa5UEz5w6
Ur2MM6RaSP4+zIfBeHYGTrULWK9dMHCYnlSeVm97TZrqO7MqG0hzhNKnD1mfPkQtqh3TjGhkhanY
0fM+0Brvb2rv4OKldx8R2vXX8Sj8xnSpsbrzasgOSX5nleBUCtykxzXLlc2al5G87rJaoO6u8sAN
14zOQ2NdqSo144AVDzjcqSnLoGJTWxeb1kwV4Z44BF5FPj9nogQHXGzfiWH3pKNhBWQK8gVRfJED
up+xxikA5JBIqjHMYdvMTX/VZOE5PaMwGX/EQgmn0iJStJ/m8ly+A02NdYJ2rU0+HWGdvFXAmXio
Ll7/syJyMQJJJA7v6JmN020LwLKPzpE5AfW06Tw40khuY24wpVWqUsWxCG+7toYEWou7b9mFOy+s
og2btu+0sOZxZZrA+xBvq24dByOWUeTsZ+cTfQaynJqQVcPsNFaizDYck1XKEss8E0wWTxKbDwUM
NJmJGrjCHGWB8D8VFI1/owKZ+Bqtws4mo/fovFwqXHm3AC7JGRiWI6Msc2QyihpIjQCFq7tkZzUd
3pYcPZxWRSnttzcm7IevMOrhxpovSeZ+hMRq7HlXcCre8Zyqua8c7feZ3W1OMAQOPa5ouA6FeiJi
3DXM+G5La7qwDe/xMoAr5kYhE16XHM2hVf6XO5Jc4siGtoEHq17gkHKL8XmAIxbJPokKKwSpT3Ot
rcrLuxWc9cbCws0ZjIIYxg9Ktq4Tgoee1+evJkWrH/DCN0pmpTQiqyk6Kda4U2CHYHUnRjrQcNiT
IPwxgfJStxWVWsI//XvuGPY5gazqpjIkmtm+aFKcVGnJ0rcoAfdTFgz9f7hsTDJd5uY59qMhUF1x
oZ7mNsznBk7JBrUbfgIcLyQpL+jaY9kXg/I8u/JFmAxr53HGc+fAHcRIImAZT0dmFnQsL9ydygpN
SLmMT0Wc43D3aKQwHa0vax5gRW6Eu+yJ9Kaq3rqKWeJGaZu75CWWHnTfD6254ke/Yz3vRz5HLzJr
7gO4Gub0lGlqpS3Uh8xMw3eOYUWRK1sI7Af95IHuO/juI2ffRL6CtcGlcOYTbHzAwBWGD1vK0pTu
EOP0XlgJDTQHyLv0sYOQ9a2NeRtnLznVlZd4XTQ1W2myo+yVJ/4IU0c/uC+nNFqyldLuc0pz5gQw
ChBikP8sBOapmShDFDmTTxuGP2dHob23C8GI3TK039h+v3iDd8vlblMEgKdEegHy3Mk0wv31l0c4
1r2DqbQg8/faIXU676Mz0SsxT1qSSALnb81kpl/39d+6vHtFGj7NNO8DoFT3Q81lwLoXipZPRwj2
J2kfBqQ8rs4qLi1z17ICk+aARAjVSc69412yjbgzdbz5mbdRO8AKCBAsqQo5Nu5mnJDgvfQlq6Gg
W3NWg481zbp8dG+uA5XMnT34q8SGed+r6DozwxAzplXLg9sYemmY6AgBmCVgzMiAvze98o7K2cm+
srPuAf9IhDUukCMz0DlFrn9yqZjwsUitUc8uN3uo1ohIywdhFmJIskPhqYPFvDdJSZkHnZYfjQNm
+68q15zqNdr6LjLBhDI0m/bz/PNxI5/LjqIuM0rB/TkMGTZGDyc8d3J5IeWtkzYhLHkQELf+pM+Z
pp7c7Sg2R9HjUf25v9aZaJXfEkI2BFv1awpotECRDtQAB28U+PjG9c6WKaKi/67ID/zFztvTBSjY
7tTDjCzNnBc9JQrjcln2i6Kp3uRyTEWfN95dztHAhBZGz41T
`protect end_protected

