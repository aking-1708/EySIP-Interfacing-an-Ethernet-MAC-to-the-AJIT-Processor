

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UTmxs0OkmJURXBOVdUGR7t0vPgcBU0oVnrXWTlGh9ogLy+aZVadnSNImcgn+4jLE3/0AXAxZXQ82
Xbw5u5ikwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NDHq9z13OnSHCjB5ixLI6v+O9siiJNJuJRP5KO7VWFUgsdEdfLm2msHdSHMZWHSOwKZ3fpyDnmNx
BgNrMCYycBeI/rO2pKL2N4HQAMnhKOZtiPFF9n2RUplezsx3A1KtfrZPlHnD/UnZMT1dsl6klarx
WHWoOj2BdFWF78jqP/k=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pd1c/MzUc/ohRsjBZ9c2FYMEVEx0/T+c02CO5nj1hjCkjBTD1iExW4b2fGAqq2hXvApptvjN3kao
diEYImrFYF0oK+4fJDQ0NDCFSHEPkV9IuYgpAy5fNfC1Dx9rVAZAI1tVIUXAIZsy7oaGc/ReA3s3
/Ev1+YSM6X62ouq0EXc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ds2lszdMaBUWm49P9ovDqEJCNyznNiiJV1s10TsqQV85Goa2s6Y0q2oK0nkUurPC2r1U/lFQ6UkY
FyQj83Ie6eOpnawKkK55JF60SUgc/KJzJ7bDwIpaZjrpb+XlrqrzZU73J8jBBHKLoF1/Njgvn5Ad
h9N2MGH8gaas+uT9uDuZCA+ii46LQ3K2yd1YWXKK4uzoENDnOnWVcV9omYQiZt2WoMmuDtnHiiD6
BU9fNvTDJc2E+yqoRZLq/i7Vp6O2raEB1EabQzrK+1rVqoRBidd5D+df98jf+SVXW4uK81yOCvMA
LOV3/ZU0qCRQoJbwjKLC39h49ly0sWjEpfW/gQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
df0vCAvcFSWs5BffbtXlfaFIBd83+wey54D1uX3YAx267SlsUp8LU636/ulbSzkGShRGyHAsajTQ
lak4/g7ql/uNS4cPDTprvz1MsadnxOACDABIUOl7lg4w0zjMlnHliJydcn6lPMrRHgqJ6QJh1Ypj
8in4rFzqjprqSxw1d/10YsZZxkQoba/tmtftne+6yGg56W2Fvkku/OTLhJ4+2k81Et3P6Hl8rQs8
H3zDC5jgcWutFMz9ATChQpuoW1Bt6ol0u96wp5xiZl1ORv7DkneMNq66FiXR7uQAikRnfSIiT6/5
QAjuFDJ9beaONJ/7PX0YKv+VUGzRFq0ZFYEUEQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nCZ8D9A90hmHjnYoY13nJu1ipj+rg1ZVc4+qcqLwK/I4sVkFzYXzOHfQZXQ7YKW8qcQwr7Ja8l+y
rmS/aej2Bl+/GBm2e8OPwXjYQfJZAcWrX3bukYUhs960X48k+oy8IM2fpLqIO5UjCHWUKDAmMH8s
veeZjDOkDvXS6zx4x9hZL9OB3MW0oK6L//tk4UtxPcVZEJmBR7mpHfQdetJlD12R2NEAOMEs9GYi
egJoRgy2DcxVo/qhMUxikMoNK8DRbPimHxnf/gi8Ss6Awc1pw8Haokg7dho4WvcGQs5jULvRh435
wbmLZ1FnvnxhHSbLJwY8aBTSiBsD5Jozey23DQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504800)
`protect data_block
5yyDy1WTby3EfHlpfofncqpl6a5Ldvu1f0W1GZGFgFZn6LkNU6XREFBBS/BFqrSnBLB7xeeRprEJ
Q0TSda58sH7ghuM/sb0LNhyGEqoniI00MBCaM3SWsku3JU8XVx7zomYFDyTi1z7VfyeFucXflawd
mENwtv/PRxLVHqWfsJkqiqfmhVv0rl64LYtXTQuUfqNFTAL2ZW29ZgQqoPd1KESSVcQoVsjzpNvq
SxE7IDDmDt4D3u24VcchVmQMOsUyS0avhrCfxFh4VRF6GW86X3myYAHFqWbUfUv47V/KJRxSAtn3
+BxjPCrGU7Gap6tBpusO2KFhwEdR72ytb+BmIFkfLkYJhnJO3CSBhJTij4lS9OzramJpxat2owD6
xjz5sEAhqHlW3CdN2yoTYcFur6UrK0uAD3sh157BMxwDT+cQwzRQ4rfekBUGi6jBvSCJ2iyXQSZH
rUjYCrklu/8RyQLr4bACFGicMK1dEPZQelUPOrq2CuQ8dBUwUfbHokFKGwGhWoBjq+zyHNHvcvnE
BooMVpN33Yb53tkLohFG4b7y3rcVmiZNHye2+m+Y9kSLY3iYbdrZnPQsZN2UApt1d1s3jDZi9nMY
5t+mhskTpznJofmzKLcUZHHjZXWVsDjqk2pZgGvefOAQqhCu8sFFi0P+tpfBkqDTy6iIn7OEX/gE
VPQ+JTsOcs65gE1dGHScO8Pbiet/ciAk8ywH6JSnonPsAMo/uzFlTcLqcePGXqZe2GK02NFd9zta
FvksCyL4MAIkK74cGTqE4P9dCw2VaKHIzdXMrkTtjabBo3y9GrKzDVdWEUgy7vQUq1/9zCtewR8c
U2y3z07Qezr80idS6S6xCqcyra+kHO0LHt55zxDN4XCQrLUlbvKiYVZYP1uBgVjK2YbiU1Fsaz4E
mygu1OG3k5oppbcTlhHPimvddRekgsh8HKI0VzA1AqZDOnklSDeztb5ea/6wWH2kRBKujFuNfzON
lowP5aqkyWkN0yYWL9gPDAJiB4iBdqTSBAIsjYBqcbScAORsOVJ2o2jr/OeX9bvqnogKxxRnsma0
FBxpNvWE6pZGPjDnxcr3pCr4lN9PkZ1OAdvrpR9wse4S1Q/FzFbtWZmTzbjCnG6pwmT2p0Mk/t9m
BLlpanuI8tGl8t16tkDpBIx+C1dINc1TdEZCvpOIrKrYVQrR/rEAetXsjkhXDYY/i3Kt4L8uKWzO
G2Hqemw/Ya1ADGSTZJjqGBifQ7KFLE+loeK5/Y0CXIEo6B/w5kK9d/k5k8/SeyJG72Ccw8Lnan95
vXL75VLECTpZ2dwv4XAgQ9xvukd2moaFS11dNpSG02pkDEXbo9NeB/SA98UWF8bVoYL97SOz4wTl
BGIAkpPFnPPUz8hw7elCRhuAQase2SW29qGjSQgtcr6NqmRuCwb8nCs2dAjT3ZbdICzuZzCFncek
c6Z+36ljcXmanGX5NcN1K0q+U9tIqHnOmybO/eToJDLZwcpcLJXOlgVwDMf2+ttQRknQy1r09A1G
QBNDpYlLF/6BVYsqjzUgueajnx4WfDVFI4oQ1RQNCviDxRn+4YvDKLWewQs+LfQsIPXLCC7yQuKm
WbkCswHhuel1lo9ChGihEzXLqtzVQv2fIVOMB1BxcBOXQIS3u4xy3FyiBM8C/4mCqmNLPezgqKD4
fLAg/bFYiEx5GD9jjvkWveS5wC+JQhUnaBS0DrWSM9x6n+MErAx8HNNVi0SQC2USUFq2nLAXudZJ
MiLjOig59HmzDS0+v2io6ZUFtfas3N6IMs0eyoMh/YYDlV6w76VcmBkMGGS1kk90b6YHD7mq82To
TPit6AvQNK/y0jNpoIWbluW/4K+rBfkIx3Ktj7FHHwnvL7hKv4eEoIUHRTeNY9/FH6JdWErwMkR0
wAmd0LJuYfpw7I+o/uNZ8JvevpYIoLHIZDo7A/81yPhql0sRPyFPiqgXlMNuwadPc8fg0Vu9ZgD0
1hE6b8wbFqYQrZ5KnCCZYmrdiD9I8hfjGLsPPgchWW7cvFtO45kcDcn6Mdl7//KjEmk9SZxyieP2
hBNIkanHWIzQNxPTkn4clX9oJQ2pEv/6CUqP4kmGIbT6HUWuYVZnD7ecPtC6WgwGxs85yLbxPqbb
G+qo97IiF6qEeAe0boBnGQfUAbyBgS4+62kTXDwaikduHBHSSoJu/XUP1/LNs8L03To8LMIbjaak
YNNR4Ip02sojecBRguCGvXesO1y+VCFuhvZSSTavBepyN985WvBkPi7cmfnbvIpy32O8F+J33oBO
pNqY168jz1zo59/7wY+DEsmM8Y04pZrY7ugdBymZ7irW+XbuKr4dlbOZJhnQHi8qPAw9L9fVTRXS
LjWh25LYD6uNg7fTgVUs4nJro7cgrf/HjmVn/EsD4okg4mm+dMPgrlsxYSd3qFYpJpv5WiFutPQE
8Llbm+Vu8IzgDJyo83KcPx2kUIPBXF4++n0KxYKTN12rbvRj8Wmx+ssTnBvEFaZM01TnsPa/yw9V
GZW4AQX7PEZRBl6qISyNKKVcQafZfGbrf40yMd6dL4cBjjW/ixcP3PGp79oNCpKQwkgNyjTF48nN
8hYsrQkQq9l3fZfB3JePOX9nv9ry8cJ0oMKU9i63YwQi6Q/Yjz10gs0QTvpHJ5/HX07ZEEbAtrYZ
SyVx34qGGeAv7L+CM7Ld+Qtjn0YfEYHKRovWQL1pe1jw98WgHrZJqb9Zwo4yif2WSD7O3PNGR4nP
O9BDiuFvVldMkZFLfXoskR5vkxHBloZpb1x1Toq3szYhCioEK2/0OmD7GVHYyjYsBeGVwRB9cr4W
FAQxYOA8YIKZqBXKbaixmn09drxpsqWQkw8xl/2Z3AeF71HMftrIGtfuSNgVKGsvsADtK5r/v29r
mPzpFrlOZr+wYWAcDZa0Hztg4L5udY6yaPhAdRPcb/INGYqilVh/07I0sM6Z2ij+fDY2KGcaS43l
enYFmxX65zzslSoSUb0QWxjYeWqnIXuQ0HuL9rf4xxUJxsFC0A/0Tpz6jEtYoFaLQDfiPOcixVYd
wKpJcaAggtbwI1a0w5wpCZnQ9gT6t3qmhzNkCg8si0zIIKrkoHLHG+WtiJGPBNOlV9p64egraSEt
qkhtHVce/am5AfntPvLLZEyOMckusgjYC4sfaEIzLgHHEyzahaon0bhrEm7tyRRIYMInL85WmdCS
k7CK6vDZPMTE9IfSNVHvXh9sYgOmlZqFBEIWvYByjKJIxLt82B1P8vSmFj9nwaq52uVJVO4Wq7WW
38IlI0hR73KdMhqkOr04NRiZJrDLmYAFTh8W4YRA71qlGJgxc37H58viffs59Jrc8NpTofzpVwGD
OXOiW8Alba6OqFXsNoDSHMhGsqOjat04L8cBvQiwgnjus4aAbp3/lN6el02C2Qcz1LoGp7HzDx2w
ULbvoXHE7gsPhb4tx4NrpqzlVwbABaqOy1QZNTn2sBr71Cb8MNL7TZrCZbpAbxLs3Y6U7MQKJxzi
l4cxDTWGWMOdNyVl/d3MTC7bfiADjo/rWi/wAW7cLYl7x5EcE9kLeXN21QzUaQUyNk52gaL0k84s
7BP3Dvz5lsr1zVzNRLo2v9DpWHpA2T/kRa3gey7uT3VOZ7fGEKIsGdoVXlIEb9vWGGwoZe6IFrkU
RkAkdBtpL3xG/39qu7D6BoSg5tNsQG/17xpiVCzhNk8abIb6hM54Fyq0pk1+6MdpMvaQTLb9xEHJ
guznE2cL+57G7MLv0NBuErTQNkleD8FCEyL67KZuOeOqQcsgeBYP8QmR5ev0TBZRKojMbg5Inw1P
IAclorTRbEFiY+DIyIHaBJ0wZ1LHjQBQ7grllwcd14KVClSY0dEBCdvBhzCGyvcTU41uyQAKHXhI
h847gr5oHhibEAKb87Ho/Fo8onRWXPOVggKuJ4GMznpzzl+8esyOhWNXUYiZZRrNLaiks5zhJwfd
xruGZ9AaKvwge7vqG4vBjxwTHtzrXGgMi+JBVq8GDQmG/MjKz5WtwNF1OTbt3vbqRXwITBldHLpl
Qof6E5+st9pMqOMge1iRDRPaURobyIsEgdxZqz+PUmr8n8u67PQ1L3SsyYTqY51ztqD9un/VEKSl
MDVztiOzW9hgpub+385zLcQuwYzvP+ccZBZGwwsO2spV+O+JCF4nFzdiqgfuz+8CmNxu0l03V5Pd
NswWbh6Vuo2mbEwfX8t9L6WArPs+QklqF1bVLTGh84NTKDXMzeZ1RZGi+0IlNMrKLO4M5mB77Ely
s+gsNOrUs0WmA7FTGgkiEjPWaPv1QOix3DnJLf3aQKRS04O4p+o+K7k2YA54fRlf7hc62mwMTalq
YIP2RawxwciyKUM8rypKFnSJeQ8176fQCdvUbYZvReMQC7QmyYN90gfRLq6BC4cgrLa2umoAOwiJ
t9B6RR6ithtxpG6rdtn1Mj4Ip6KbaOrxU0SZfPFvfgGi3NWwWf1VnZrrabyRmqdP3Ei4jrWquSRT
Ri7AsJapXrYSVOCeVt2+noiRKRQRZ91bDszE+kwJq84FTlZHPfQ98ULztwfl+I6hmzBLsxJqbmKX
3BYKeoWxoESQWT6qm3Cz5SFQny+g8BqIMCRcebf4vIlrvMFHxWYPGnPiRx7wf+Y9jmhSnCGjpqWT
le3QAsdkvYBlW57mQ+3ldSuRRGr5FnVn0KUi4RlPdLa8pIHPDOBXAMebHj7Y3+nqNPPtwP1gnsrX
Q7OvybzEemEIVixP9Q5I5x4m0fsVvgK+qmF7FxhnNKjMEssGfYS2bVy4v5CAyueWNAlOMjzM3i1x
vcdjEDFQbSBR8YquHPa/egZiX0NJkA1Tmw9hOkBl7wWGYy65AgYUZ3UL4W/kSwOg/Fa6sRoWlPqG
YAi/hEeVTJe5cNB4FEUHQo2+kgQO3VTmtymOv5iacotB6NfuQhbwrhpEH4PZ+j/6J5geWmaq/ZZt
gsgaRY1ZwstIAY/cGrLL+QKkDUvvvnqzVWNnCDof+6IuFvxAaKtI8hoqVTRfpTMLX70B4KaXBxXg
c+lxUEOz1y9oCF+T1BQrvWEaEL9z4gR5Ik7nJ1S2weY/qUyNE4HtN7mm4TyObf0FQRZle1vEJjDH
DowezzvCofP+2SDOIrZohNXDWkczG9hEGkqe0/LP7+a04LxHukOhoRsUZU+4mTFmYhDfnI4KsZsR
cqt8IOe/P/4d5+pFfk2Xq6wyeksjqPE5wyvRm68RjbBUD9TCttk6wzCS7B6SrMmES6/cSixo7b9Z
HucDzgcQKydgpva/5l8BjegYNte3Oiyd7MHGp7mKhdtbwMz+f+eTRj5RUsDb7ctWqbyodfexfZB9
le4U7Ms7deuY/MSthX6FL6iu+y7S6GsZRkF4Ueo3p1lPBGUL9FWQ8ZabCvktahZv+HRnHHux4DJI
fjMiJ3A3Jbu5BQaGm4EOOYxbw7adPH0oZ2y0m5/+kiQmSUUXTiXuktTDAbeqq4c35qJQemyc9JMV
oLugo3q39SF06V59H8OWehuS1qJSKvkFotPwXi4H4WVjLUmotdNauEraPhnBQiMagM93r0Zm2c/l
bPFk2AjAhNCAlhlyOPyWyZ+BVf93YnFHevDIemzO7l8PwqVjtaIoJ9SzZydkuv5d2arhssLvoN6t
thMyCdVDWwjVB0zsEKStIkpD/jVSdv0qTswKP45yBBF1S7FUGKAjTMmOq0D2ep5MNUXoY2tb+5Gs
x8W/UkX58Ti2A8bnpJoiTlPUcdyOrtmyTb0+arH5h7MQc9xSBo5O5SHbipJsqzvMFg594AaMQJwi
uygILaOpCHGgNrM+m0z0FxnJ6PafOZwDUZEbGAsnLyRQE973pCfDy5VgzN6HL0nsPooQ1GyZEZnK
TqtLVRZiJrhlrf6DgQgkhkQn5AkOcy8+xyIozjX4LXNy16q7raGXHXRQph7EMoR2tF8BVFIek2MB
1gDYgY44HULKcPdVdS5my3YBAFnL/HQkwgehASH7LIlXbDL6WXTV4QVuYPw74mS5sVcFxRbKAJfC
B5x3jgWEtEeWvgiM3E3vJm80BQ6BQCFe6qdjI7Mx2Yb+J75g5Wg49uo84SxB6KeNxAHY9Nuz4w/S
l/Eale/Tz5GT9c4w77G1n+pwZPzQJwTRoHr3Il9qVLJSwfPRqXqRuFDqANIANY6th/YX0JKf0BEe
LFn1V1PE0EMjy/iLn7JvXbQYEClwPOkvbk6ydVrkB4v3vwEfYGzvH4DxlE98aJvsC8S4c2QLDxcq
V9uK7KAyaGUNKMJf3RwwxdRIpRNBqdWfq7+FyLThKGZI2vODEIxbBwyOuj9bRqlJaQAZFaXxN+KD
haPzTKpe+aotWgY0xHDFyqAuUuTBB2DsQ355jDXRJLEUu+z3K45d3G+DcR7YT2Hu9O+PCOOAPzuj
rsiath4SWiuDz0kRaPfz7acPQ67Hs+KERc1nmehNTzaLsPHyEqAjNG6KBX1d+SuObBvUv94aao1u
qVH6g2HxopxOtH3arGW0pjz2RJxiqrQBdR2+8qAmyUYuNQ2FDcPMcM3Aw7cO4RbtNiao2MOs5pjp
742YgLc14YKvB4JqI1XNkL67QbcllX4aNCRxLoQMgsPuzqB48lwuu1Z7DYts+v0nOmp084DIWfME
2xSFKIJnfuMytldfOCSFfZwy0vt74wpaw+bThvBW+53o0HObScV6L1jggTLn9/lFCHbJaQdPYMX8
yHpCD2LAy0hX8FAysc2tBpPrXaEPFX6O0019YomVxUApjvkzSUKILUjwX5JFmBdcy6M+3iif3ZMF
NCaAAcbRGopjHh2W+sY4LFfFCAPo2USBRLR2Em7h5w6nm2CMaQhDSl9nBcmIrTD6y+8lP/Cz0FPZ
N1gh6nZab5UNhOlTSOJPYV0Q1pg/rfrXBFfh4RRqB6alC9VlA2bx2GfjsE2zAFx/vHN8MW1Ayx6I
UJ+LPT82OK/ukq6pFiydySYfF00gu9OGhr6e4cDLqIapakbBlkKIsWDSYa8R6o7EHyUQNAG2P93P
miHa1hT6hjXHDcSmIjRc6qgtR1Sx4Vi9qihUXvkai66Gyw6BGi8FHWoKGvgVdN1r0GR2xu2Uok+x
xL1qcrRT8ek76JtSehc6TNq+boMcUNRoEj2IxF0GjvIcVAdpIEF2sUl019LUf5p2DzOEwp7M24z4
owjYxdhneUQgtKky7indxooLfGYMMNTn3ZSEIsZJ56lFnD7mGb2qomNfXNYsx2JicmL2wmgJQIRZ
F9Tlj5rEPN1xOBOqwFuPT1I9lRq6zSMs90449mZU+jOXHRBXp1J0pVG4z/HPZg4FmX8MhMyfQjSa
ctGnJWic+rJytXYZ4VcxzFePGMpdI0jHgQvVBAa9PZceq85EBt3jqxcmCv177tUbH5yQlAOzo7vw
fp7xmZ7t/upEmaNHHFjGHPnAtIweXOI4JqNe1dMKpnq1yiEs6+Lm1BPXi6P6ccXh815EYK5JrNVr
kqJB+bv5l7CERvhYhG2gkb3ooUp1qdNUIoOe47H4jsvaqE+FkTuD7+J5ZK+3kQYzkJrtYQQPpsyT
QHAOJOD/5WDSt6f0l3P9Rpmv/TcsaBpIcCNM+jiUf2j3HSDYsVdEKxh0/NUEXe2/eiwGzRCWSk2I
246+CiALumxCfLxjSOOVlORkVA7AridDIamosuqg/c7puPLmmMVYU1q5YBNyvwgmF4pBKdgr3zVP
8Qzk/KqoLaAi0DFAoZi+QqGpnecXEbCeHZd/9SU7xHLdujAwhWRrot2c7IB1dOKnTEB0lZp7mbNa
1kKuQD7KT/maHYZqIidD94+ELOXvOnHf+qip6QzAvpCqa2ZC50RZjqdTpD645ovL78mGB6rHkxnS
L1vOH8/dBcCaVEy3V6AYNBmuNzBJJFRDPwciKLayIsXzgvLidN9AgsluyEnaAgA0K6TWCc9Xc5Pu
ijyOI+USZ0wTuX0lHA5LRHRjiDZPytzMg1OPX73B3mUn6HzKXIjYz304m7nKm7uuZRMTtkkmRnro
mpTBYyqWtKd8DqFqUB4FXZLX3X85TzqDwkUAK8ZqQhQGRTpDrdw7fODVOKaaQ997JreyH7pz/YJU
6m6lMaFKG8BJyEoiERYmmGkg2sRuxSsq3kR9qN0JfurjMx6UQCAbIofYJacTBzDQ6QkKsk9eZ5hk
UUVEEinXIZD0+f4bAhsQPRaoqlO/8jL94xS0z7tQzA3tUx+1RoKmR1wGNRPoHHVHSC1RsPW7PAbZ
t6ZsI1W6oDn6IRIQ4BdOhwJQRd7PEtnS0WdVh4W5eUAmKRjjsx2GTjpj3c8wgjYDmmAeh0byxcps
jAT08Ryo5Z43HXMEJMUOFVQqqEY+7KTYiaCnOp+SVutHcpLsY0hDLBEu06y8wK9ovvmKKhsbWkpA
ikTQgE54useBrhfjeYhDxFhZzBIeL9MhY3y51AgGRtelIxfTNAcBHCJbxVS8eJZm9ZZj8bCwkrE9
WtceMpFSXwsRyQQl0ulBPGJ2JQMstO/JE1uJroXaYo6WPl3H8e8q3LzG32DSIzLzRwmXNQrPhm6W
nTTN4wXech+Bog/g/uFjENHs2DHVC5vxS/Cp0OUp0er7Ko8IdFg5bGsl1YzRHeoNAK46XRKi4I50
NXRBDZZJXxE5hpfPWGZEOfBikZe/Re7tB+8eEcQKzAL30ZF1zHg/mWEWvUe3yaNjMXR3T8NGQE4R
j1bObgUq04lg9i8RTVWLQQhWDHE9beRjtEZrebwWD2U2cT3JKuAukuPuX+j/f8R3d7NkPWgE1tw7
Ms4mtHhNGx1Ml3Zx+XCVakVp3hk5GxDhDouIBKpG1OKgOSODlYmDMxvKecY7gSIm6AIZU2imY6wF
q+68i7DuI1j0qB1IwQp5cV84fvGAjAbl8r232g0RuXlk9oOpudZSW1K3gGfCFQlAJNUlToVjggbW
9fd3snNrFmR5HzHh/4dMvnTMkaBxaJ9AbrK5z2X1ryAVA0qZvMjAqc+9+BoMbZaAj0RScXYl8UDZ
c+dGWJ/qjkRPFDBqLbJ045wr6OixnOXE1Rt71MQVn3rnMttW6x0O7U6ogYjZjB2UC18zbGfDx8Ko
sarMiWAaTp6HolGDb/vuwBvTs5fEjhanoNi/3b8qizepjVumk1XGG102chYgdTjkm/bri462fmct
KOE9LPDnSIcVUZpPjZsOVcFLnUgfg1NbPx9buzpTcxZXOxRrSkXGewPUaqmGwYhyukkfIfhzVvxf
SQwagZwUU4201GUQF/C6W4RdblzSozOQCciEgqowSr1cGXcMbRONq40Eh3KmCw2JJ+6eAir75I28
LOwueL45/G4s6K8iJ4WU2ZH3yfduEHK1v9CX2G9funMszpiahPKe7FUSmcd9M8Xp+jbVXGaNEoWR
z/qYAWv/dQ+ptj4NAjENCiioglig4UKN96j2+EfS5Mg7ug56GjhRH0bbOZdnbFK8odEPkv8tZ8te
6pWFaWoJao1xTfSi8Tsc+0InGTQ5ZHGwAjKf+bR9ekvQF0azELDUHcG0W4R0tRd6vZcwIL4sqxoA
PJRqK3yhMpYjxNLmLXbS34zWlVVoKOZDoZJ0vEBzzVJLMQuSULlkh6BMiWvPpfBtmpakCzuw/u87
yWSdLjJCVg5wdB+4Z3UtcJtOO6NNeXbt8XhoVGZTTkH82LIea66THwXm8D80zTqwhjjm7u6U219T
Yq/E+zCYLDBwTJdmFeE+bHkjQJqu+4Mb1WcbHoLd82URIIOtUHYrlTL8CUAzLf76yllsEDCsQymc
69YfwfsUt3D81GUzSJj7I9MXsUWQERtNLTfkDxElzcfjM4w9QWoKjCLLIvdornkfjPgJ/evuhqrX
+3Q+rRFfhIRU8E+MHqdZ4jHi3g8IeyWwHusX5mc+r+b2pJ0nIBZGbYAWs/BUUhgixwVdOGxokJbx
GZKyM+kGQr52VgimnPGgvmxO+7rbLNT/B26IysDNuVAxpqi/xJ5PAXCya8oaiNYFZze8YgIupn0z
cjFrlPzSlbpVI1X6mMZ+oyvtx5MVCtMoUW5B2St9+z38d3axfuzov7QQS44T6Da+o1sFe5WTegnY
KbVG4VQl4OK47JidwtcSG94xQSHBXW+mFmD1dTBxwNRXrHTodvkzPzucMyLaIsugRN0RKMotDgV9
0sB5kgJavSAxYYCELSCMGf3S9RdJcsPgQbV6Y9ykdkzZHQyUCbBqwCapBG+e164jwOU+wPSx43Vg
OPky/lWKCo8jrLtXtVikd/f+ApR9OMv01pcObv4pFSENdY71zC6KHl1QsC64jtXezgrqgq7WXQiP
NtxRSXKNKpZ3gcaMfvyN9PNCOg6ZHvkTaanYIetWl6XfU+6HYYMpYvKE/f6EFpwWRJdk/47Xey8t
zrFAmTv7rKWuDS+b+KbQR0QYfftC61ggBnVHxvfxxfDoSfIEZx+4gDQPNdK7uCQi5Cvm9+GPu6q1
S1QJghP8zPtjjdefKvp4VQffd1/M/GVfH7D+AMKHEE886/HMr9dpt4K0WXAPRjuNv1e9T9eRQXrR
y50dT4fjuqGt4Evmss0zwbYBgRC5sS55FJfI6R8NyO8hLbPsI2ZdRnOHIy0E/GF6lU+Q8qGBJGW1
9WCfz7Tkrb/aGtBAanIlnKZPmPPBX4AMyySgPalwbJ524O6aeFOGAN89kdwIQZlTv+oauu7WZ/QC
e4TrHCIGVktVsRZtLBW4w2ebdIOC+MgQJt2o7rjrAWokTL67pt3zLkdLK/B4TivpkHEvUYnY0JiI
dMPxeX9Qis5UsyK9xD/ZHQu9gD0VFxpDI+cg/tRGu+/CXEX41mkz7g/hn2e28Mf5s4zXaJwozKPX
ZoSfuURf1kGkMGyXbA3/y4jIh4IQn6c0VtCnFF2sAr5ipnDSZlig7shXQUzSbCqcLbXj0zV5Daw7
NckfcC3XRh9s8oHzeDin9dWVmEHwroJPvj596aKwgSc3ZnXdLOSql8hDXRfdf5r/MdHqu25Kzvhz
lhXHiV3D0swMd9eXWcuBnpW3H6Orzc5au8PSszCCP/73WyOwuTt1kqpKmp10wlRyvPRSL/idKfzZ
dDe3ra4bYWRE578CkRVph8Oxy1nzEndDpsEMkJAYvL4Gtunx3A1pafwQLIQuMCRsOsLP44qpxZG3
uYxntDCa1JYqkj4FxqzOlntykB/Z73dhzw6GQ3Vd66WGC1ZhwHx8++1W/KHF3AsAdU76H/sfPj+v
ksL/WBUR+N1vBaJJSwPE5BbWglM74Y+t7a/dKd38hhJyOck/kEfLSHVBmsf5aSp9XC1XrxrJ2KQ4
NFxY69xA7yLlh0ez+C4wLn1zGxTSNQ6MpohNOcbN8KZKVVElWQNnOabU7kW7JQ/TYH/K63FLVcf5
ktjp/miY2P2JAvAMAZJZVNFP/XtdD7FpYQpbYUsUxIMzi5DxRL9MBP51wtzWBNSTz0Sd9Q1v3QWX
cimzSwIEo6mDEyV0Ep9nvyeVD6cmhyz2JLk/n8bRRHrGYW3cUR0Z2VXm/blKRb9TC9mx1I539N43
MONMKTALM08NXzqenYeuKQSEHEsjeElmibt0+06RPS/0mHVTA5ad/qWzv+gRbDOa0YSy1sXhcFmt
CFHXlJFxv7YMT8NOVfhU/LsH+1jq9h0WXsz/z3NEIcU6oMSP5VjYiFouFS8lJADzDaNY7g42fneM
JLMfPHd2fWhVIcLtt3ocEfbVxynDSjxcVL7s/uymzA+yoY0EmzEwRJouwqOSCPF0s8eCRRd3mR/m
9mlVt2oG39wPV5ybitofVzryF9oks+yXOIB99hePSsh9LleNKjPRB6Ml0pFbSOCnQ+Xyv9FVyMsH
N7NSnY1UjnysW/EcN4fxGdcjInUUit6k/LFeOIjO4+coe0T6+bavqlCK0sCsWmDBcnmw9cQAn9MS
z6TQ/WjbpLxsdExvD0hIlEegKRvvGXa6Cxdv3gQFbaySHIGQ6hb66Y1WfhIBNwpDZFwcd2ZlmDgP
89V70GYALqrw957SkzlUW5zvJhKs1NlhfTP0NWdZd9IR4vC4H6/+637mq8F4anVqyyuf47W5wfTN
d0JZ7hZKJQuBnBFuV+TE75lfE4+6O43xdbQe+fuqoXtQxeCb7OmfMTeG8JjYZ5WLIZvCFrUXQV3p
eANtASxa5C8nyK4y8xIa3TjqbPjYjRmy5G93fqt1uybJGXk9Y/XfCAbIry+V2DkEWj03gaTHCIIO
Q8sySByvp5rCCEM8iEQ1dFgxBgerj5NBPGNHwUCb1256qr4bWEW3JggtEb8XgI0X+QYl0TUwkxay
QfdOi0qwthEcZCca0tEVoxmKmKGIuUo3IZ1e4+jxRDru2GNeCE0V1rfrfXY/k0Xl/Q+GU0dEd/+Z
8dV/H7GQy3WwaDZ24iAyKOYSqxkSwRb7x8k5vcSbyzhWKrq7KdPTpumNmnHyl2u7IUkzBgdI7qWT
7b73PINFr2XpyhNxjRnXPPlT2cDtOwutTXZAZvjqGRjwISKb6PNEKz30o80hTXdmCRsphR60lQzz
aVpRQDwgd3i940s+7xsOr+QUbFtjEEg7ccIQR1V9N0MWk2aBz+8iiqE9gJo01fuWOUD+aUmPu4UM
WCR1UXtvw5QznTjFF6mb6SiD5AaKC3V6rgRWYFfBYQO43yfc+4qa+DFjbyS1TdNm/f3vYj1+mm0A
dKq5XukBzwhBHwtTgJE8VfsUhP68ikpjaaDUsVCt8RlmFSA31cL9ZCP3NmFO5FIF7ZfxzELODfha
Y0FSlrvq3M0ln9OrpKEm8Ki6p0WVwAfGPX57kRtM8xJMZZg/K3/8LKTMWAeVOOxM7wmdZdwd2Fl7
g7dgUXuqK7lC6aI91qnbIOGKQQDVdBCE3O63aRo3l9C/7EWvjX75TRUcbw5h7J8u5pvDwYJ/tzb5
V9gnBBiB/s4RUfrBQUvg9U0lEOcHF+kfwBF84RY8z5U/cw+QxjUg2B1odOnUS9b7qgYRO0UeeRat
1gpJQPnwoGRr6VhfFu7d8b8JsBQ1vawvh70ouSr2nWcAklYuNulMLAR1OkmYmjkvjDFdNx+yvIHo
1Ey61ZkGVAK2lyUbkZZchz2sun8uRgkMIYyxuTUVaOqMAsO55Q+Ky2xN0miAbT4oLZ0pSz5/2aUZ
ouoY2hm9W8/e6G4sLidsETr2uGW4n/KRIcooFeUVdYYo8cV651/m3BJLczKoQkAgVWyL32SmciA+
qtozg03tSxSTFyNfjqeL1iZLDDX70IZ2QxTfKjkUDxKu+VW/PUdU+0iNWJYHjcPsb2mNonSqMKzH
ABoN9YhobCKxfJGEuKicVmrqjddJO9fAVJ4pGBFvn2YUzVr23jI10MI8N0LPtgm7iUkRDH2TtZQT
baUWqn1LvgLjh/FmB1yjuuHD0ZrgvSz5R2K9+VpqRxydpFj16O9MSENQayBnH1IXrYUtOlwS/RcU
TflKP9cVAR/7XOVFSDtYnr1reYFIfOf0Se4YaSiHQtXQIt9WDyaZnKicr3w7360fqKwE6RbKluM9
hE0C+TIDc8jR2JwwW8mtaL+/b8ZT5bGi7NdIlYtlNUUnObRD9hdXrjtN6fWIqq0iXx5Q3OIY7KPc
wv4yNrr3QjuZW5KKaAQZCFOJu1jIbPzi44kou1iurtSOuC5F/qEoq102tcTR3Y+9b8uu4YtnaASi
keoS5+Zsmi/yiMDBcU29D4v879cG9yC+oiaiwkZ4asgoE6opTlkcGObQIvZKjInhxi/pqdcSB+cm
IiLPosUmK6mjeSaUB1xoftt/FOUExYCQJAJ948DlrSt65a5qcA2n2iAnAaigw6oJNvZC7gmEOw5t
tpZR8R0Zjx5QZHe4+5Sk2n5oB8t7xnhE4YyMYAv5UhhqogUR1xgzbxun2R9txi6M9bA03XekZIvn
v56HyzDnZ5wHgQ1I2HH4Mh34uYA6sYq5gu9qejTGWJlKhSv9JWFRRee587cDEfZXYtyayJ23SuEt
KYYLLZdjO70UOBD0P2oIvhU8sdWg1+eZcB4ZIZNGj5MMZThj76wnpKHmjcR1T/iJlFJeEwfL5NM/
J9a2yF7lZ26C/sXqMKL6WHX7vIjJvZC7EpaEHqhg59PICJhQ3EsEewJAHRuf9dw0iHLfHc8xQI0Z
fWerpsT14lOHSuN+bMzFnrQQFEw5GuBI0REGPAKD40DfpGCWi+PdGc45j/DAiT7mL/PPJKt/XQMw
aePXcQNOyieLpB/q0oq4vlTVwsvRSSjwakEaU+X3P5iplhUILWupww9Zkuw18FHbcBi2VKY/0PCD
wEk34La2MQ7eMmRuhuloeDVtetjxrEeql395SjXOtz9KHm7EF+p+WJrAgEtwnT1Q/UlR63wKjWgc
lbPex2/Y7tKtLHtv48vyVZVfP9Q/Xjql/18qeExko7/DOyW8JxrDqQ0AfbY0Bymh9I/eyw+IgOae
hr2/HzDgcHh8m8egzR2xcs0H76Jra1rf0+BOzZdkYA5ai1vULVZSISz0F7DSdVFuiCUvJbZmU+3p
FsK1d5RQZQNaAzGehXMkYVPETZrDozpmQ+0OxkCV0Hc7YnMi4vT3d/R4rSMWUTIIqya/UqCbPMQh
nSPQ7lIhs9O4sSKsJgd9JZh0UUAq4vBvSnitTudPR7X4UDtgHFjHR8X1KxfZNeVLVyEQpdHO3DQA
fkmhvy6v3JOh8MDv36TGeM1Vzdbog6UrgqwzyO031mMnWHzVrnHD1UNuKgkbCa+ZRp8uz0iM4cjn
UtNfOmZ7W+KsmGIsqsD699J4OwiaXMTtWChIEiFGhg/woaEuQTVXZL3Gq+KVxU1geCq8+W6CQQuO
9xMl5Xs0GUmCKhVIoGn/ZQjxn2KEe7S8vRgGXiDcF8IcuH/SHg967Ow0yJxpRd4PynfdM7Ao5qo9
zqLY6wxiGlwew3ceo3w/wJPankj5ofA6HKOJqelgvueLAUBvi6c0VRGTKjmF7XzpQpxlp01Q395S
heL237MOdZguIphvkX4WDpEZP9gUpSJSVBWE8LyvLw114vx73pC43TmnD+sZd/2h/EV0wn1KeCxp
UYv/G9wQOiN1ehttONQw6uoiYmC7gDQuua4rZGN1fAVSJRoIacVgUCr3Xh+YUr9JZvwFRWSuGFtb
QnnAb84AEpEUtnNXJ2kL/CZm4CG2Ak2JcSLlN4GX+yekTMr2/x74snSJSzAgaU8ZutFXIgNe0vuD
sdED6bupXsxCWhKhrv03ha0d4Xa6lTdbG2zrifEf9k1+1LIdJh1sU4Ghn9SyFONoL3+ZSescgutD
qVDQocWfMp2hQIl+pbzCHgzDtAQeBcZXN+T9uQ7JGCwlyv8JFSqMrLenNMlXbBqfn+OB4PPADm13
n9q1Uo++CL9AywKHN8s2LMsMrOownZSd8JnXB3lkDTLQvfN5v3TNHhbyBB26Knf9lM+9UieZwodB
P/RZdiZUiuL2CDrDtibEGlwTuM4RtucJTKowX1YDZqKOM6i3zAsKz+kR8u6zCIvPD70wYMtsU2hT
peJyBmeajohH4JE6L+SqVgyeJv9wDhxjATIGOyEYOAE723PnUGerl8vaaPJf40BKtpGP/xKky2jw
/HIlOgEk9/xzPrZrggmoDV+a0k2UQq3NzyAK7uqy64uGwKVhRACh2pvC+8y6jjJshyK8tiOJKSUM
wcmEz0noGl8RXQMVwJ58hTNnIgy87Vtl4z2t90te4NOteTMO6TUeX7u9ex/PfxvStmopz86sDLfd
QTOMXWcMCHxK2KVp35fS1u+VZsD4+sOohBb4kEOT0PuxlSkoo8afWmBBvYSfDhqJOAejuFxq5DNO
wm4wKfhcyCZH+qJwNSnD8WklBXk/hAxoJi9xvFUAGP4SGeBs5wRqjf8M+FzSxofnokXmMmTeNQAm
W/8S1s9D1MCeArvLyGWvJyncv3C3NQzYY+ZegALuxlAn2AkDT/oXxxSuIBPG4FvYOi3TiYKwmxD8
F57R7a9x5Ki/LWSHY1uiyukyTo1TAY3DUvb0ZXGEKqdbms1Uno2g1RPmZebz//DW+XKryTPUnV3U
5mImIBepEjEwzE8/BBl3a8/X3oXiEnfsbp+7YJMebq9sLm6yvBBUsH2miYkZkn/Ry0CtzJ8BXjhc
/If92KYh92zTSgzGNul7EBbdJ4wAskL0Sk4kG5einepn8XtfgLHYwxfuiYAMxzoc7yOeN72UWBIP
PdRfjClrl+K+EMJdt+kNsNufeeHSIph4BY1RvGRPcCERiD9KNKgh0GnWap0huWByuzAM7BdtmUS4
Vft5Z3/oJ3SIHfPmV1KI5gTRLLHEvar4X3QfVmBwkHLDzWBHI/UoZ7Ktt51nBFucx85cCuRhNHmo
32EM65hLC99rMvcgeMsUfIgWLTwcbVpOyrl7JcPbc1o5fFJjNxqUTbN4M94/vmp5jae53rSu30eM
w58TRdmDu30irYPHLjPFpjZdFPkvO9Zti5/Cy2pKtoEFTKv7wYj9bi6RUmhX72JT7cDr2irfEEPZ
xtt0ICwmD9ZeFpW1LIw1G01ikggniClMgWJN54762sas0EgCuWJ2CE7kUSxgFGJXddHE4ZiKMxIE
VjYPrwOyNZm8M9cgND54sSyrzrR+Neh6UBqdzX266Ou6/aihqjfAR/yAT8ziaK6A1c0EDv0xXXGS
qdvrB0VvToxzLbUlJypNKrRyi2mPJ7ufRnUdhXtJtkWtXg1Zu+nxkL1U+GjPnnMfubStUaLoS0A7
qiO9JJDvlRV9kS+cw6sd0jeQR7kZP8rd/zXvhaE+1jepg5Xdg1A/0TKh5Nu8ZD0DnGtuQcnSlVi5
6/F/U9sW+WDW/EOIMaiYf6/x0XM4tHzqgKK+QDb4Hp+K3LlFAsjlm5Wn3Zu7P7UKr91/+3SGgDNI
0qdtr7kYgOeP1ur+ePkZtlaiNUiqG3KQnDh7BATVQvcVTzY9xrF/fjjt4kcuzpO+rZ7/6rYf8wV3
rAgTgVRo6f13H3nFuPA1QXccy2+QAQjpDeDukCai2RIMnrAQPaRRG5qsW9FmAv3S8jvB0JXk3Nyx
/c7Ix4i3mo7GW+GkLW4nC1I7XKQE5eW2sbIPqcWxTrxsCvhNAbKhf9yWs35Rt4K5eQw1Zkze3QHN
Cw5uMGs63tWOE9fufrjr3cKlOlMgFEb9ts8w6LRGZ80288sjZyAcj/317UT773boM3be7HvyI98w
8hNX9Z348iYTUbGt8wyW7MjFHHfLpGU/jpAj6vTwl1PwLmRY4w/XY+uduFW5SDVU5zDbsypovqtx
p1YXO0RPG9eVq+VfJMNo7eLZE/zNn/8VLQSwv/drqFg0JoZkiXaMR91Z8+ZpqjmwR5igyDOrF3Uf
ATCOkCDchkype6iAquIHucxm6F0uwv1yImLZ2tuewu3scoEuCnr7LbaEKja67YuCyeNtV8z6ASlm
rgVCbFcO4dfbk+1J7M9Scgk/H5cGg6dzeT/2xc31ehxWQS8gjp0iRvu4ng3p0gjLVL7c/yEKlKj0
+fdd4vGdV/Aq8YbrTQDbM4Uo42Z/OkQzNsiqvm2TuZyxolhmxTHWu1LetURwuVv7DXFJoFSBioHw
uWhu5taNBGBuBlDjP036OEf1ryhKhYb8nZtiyOGYhUSze05im+9hdoZW9d5WChJQ9TCEDkxmGr+Z
6VLN0idn03bXebbihIDAfPE3GsOFmKKZyme8H6FcJ+6geVnjLvVlMKRKP44iIB9Oq+v6GAvdMcc9
3emRy8iAskoOfxvb2lgmzhY7yRDCMApFyylijZWi8jxisluOZXWOvBVNs25oRNkC2CmuSzpPT/Ve
es7L/3kOotMF0nceR7wlrPus1RWn8my5aTTcDcw9BomRNoBvPX+HHO/a7SQqouk5kGYdE50ZS+bi
YuW8cVvfA2cdVnOvnzNJE95fwY30G9gN8kbjFIVSc9q10nbZ2JQGMFPFCAW4GPakM1c8VMRMl6mK
Cw33SnEhZe4G0yi72YF9vg50S1Np8GMY65N0oiRRIlzi0AyRDP7iEDJ0MoLPUkr5nw+A+CGwzkb3
s52vPhLSM9lypSgFsmrAcNVMoe0sye61NuiS/Zgkj4ysf22DA1UrR7vdwweEDNaKOa2ZfkQn8KJA
gNZuUIbFloLyj/zS8N4csS/+1NKs3H5anGLPfN+/YoZca7Y7Gz2G7l60wXVd+KvIQlSpNAxDLLK5
pu53vVjTGXN3LbzGU5L21Pb123N8lQuOKA18YEzOW/345wWwHMgtvd7wixC9T+Cq2VpOxM95vuH3
qAZg1vn8Svlf00VSWvn+zzaoeDytA1opdKpFsV2hSbMmvQTAWuAJubQphySrl2srqO7bivdDrZFj
pq9SYyT2W521MLXsN+6WwJlXqpyVtoZItarV5HQLtlhwtGuIkoslJRJqKFJPp0KmyiyKpdQT0F3l
1O4nVY82kz1c1q/1qRiOqWx1YkK+Uh5ib3SJF9zNtlf/YpOobiM7bAvLkZIbWPIUuFCV+A/2F6R6
eayAg8QWZXjBBIDakU0DBDj+EjPETSHsu5Z9UgqMnp8EO2xSioWF7ZhhfHsJAZgr4OJswc5zzc1/
8dRZL4g52G8sGlEunIWbU7BmDGRJ7JcGPhxQfcJ8nzZPOOff453Je7BlFd1d1W1pCMb8SuCMnz4o
HzLtu5Sj4p93mXp4HnGdA3AwCnDkEmes2o0PqIWUyfQkhpCJMw+PlofppHiAcg4MnoWPcN7Y9u67
RBXqdzQlaN1bljZMmjxUNJsCAVggC43nplzYiXbstdV4tWl82KejJtZxkmC/3aTzBmYcMJQAy7n2
k2S0y9JQp1VMpJCsoBjpwm8QTbcq50Lg0ZymAFTXhBr/jkR1aPEjGVEYV2f2GHto1fxmhjqiea1J
wE9a87Cl/3Uw0uOrtvx702H/US6uhWo9vEP/0o2UU1Qg2xktXYX1zJFcHLAJJ6csgBnkBFB8gWth
bPocc+apiVJ1texMLMNsIlwIaVQjgYknVbBcq1b7/OIWFgzErYk6Z87FqZzb0v32Ki9GLU82Qc9K
43N14w+wxB0FV3x4S8R43Hs0fhR2tZhGC4T8tmdqy4GDmctCxHXBjolWQ8SEC7qU2pjcTfVhaHrI
JUGLTKGYeq1ApZtmAZzr7FWDMzL8y9EgdxD3LsWJe4K4q4ulPmEe0lhBBzxFKxZ+7mMAY7GDC79G
OXDKitUsNvcGuipMHyGXPcz9+dqQ/UHhBzNNCVp8vn9NuvvB1iNZsrMwUK4HwS+piAPHE4gyPdco
SSPLp+oSiaHr73S1zQGTm/5GHV8He9vZA0V3MZEWVqeBDeN8XwW0Oy2E9B/tc4B5jsiyTREz8x8Q
Pr165kzXNk76HlMEAoefr69Qwyn2IhSqIOIih7M6Jmlduq+TKURy79HdcACHcOkyHEJDHimFGH8S
RL9ApThJIu8CvcAZiRik3HLDZZ+8xAwjUHR344ScmGoZGGYlImtvHuRnhQsyzHYMy0VLzUGEZzX+
pTUr0125b9kHR4a9FxA+Hkz/exrw3BMFioimoincfDzd6vCQ5hzw/sCJMx6Em18FjO8JFfb5+2pl
goYvBMht026F9jpIdhnD1Pcz/FwfZbyuPLXpafsM38sdqvnB2sy/1GHL6aFlkMrl2CuarfIhyAN2
4tn8r09nphO07nX19ZHMXJKvGi8s6hH0BH2MWe4KWv8XuOX717ZGBg0AS8Px1LM4Sjm0Xz36q6NY
3UsuZcD4a0kI+DIG997kvnSyrEhM9xfD0LzNBl1SF3qo+x1L7VCCiQnDlSJUkvrGhxiIYyJA8XIy
Q14xrSyJjWfHoMvlnqtlprnzOQr+bGAQJT30hacz4p2sfj+akCnLp8MGbeub6eMVicil1LFAifpg
ek0ntPSRELsm6pKYz+t5m37Kd+mIsAHqeWnjpMqbBmY7a5zb9inzrZmOD/zmW33VO5q4ZX/ZQxHE
6BN6oGNq9SRNXcD0biDv4vhjnGOUvwN+wNAe1mAqxhdI0bpbJCYmVHzCQC8WC1vkgDmZZ8CSh/uy
Gi900gdOk4mXi9/rUgAunenIpbmY3LfVxHUSlj6/nk6GDRrXS/amDcRqyqO29REoikcrHq9j7unM
0iIF5MdyZItBpRmpG9um48D/mqOnd6Zcic3DQ7j3j5EwQJ16ZDLfal/vJe2mWi37/yz8ux3/RYeL
oYPMtt+aQuNLI69eMOiFvP76NoFQvCs92AU57AFlMWg9h+pjzZJKRVViGYqOVnD06Ra7sYoUwCJD
UcBdym0vE1j90Zjxy6PIyjMZecZeTFIFkLFid/0TZvhidg33CeFsOl6D63GiTq/Mky/qOrFjUFni
0LMjOBQMmz4RLPBoNk77/243KF8N6K5PkS6/AbO4cDqRbDCZK4l2w3Sp/cOwMk9O8uDA938/frbR
gx4cQyLdv3Caz1jGmjOYqnKpMse00FF5/OBUvfJ6ltti8pMdAK0IksFfIl756WDSqwvOSpgua+H5
nIfiih3hS/INUXfxGHg+Njt4b8A5J8zo+7ekMFCCOBlu/Pn5nHMxHwVyVqWqs26hN637ITUMgqM4
oGnQCt71YXy7HC3E9A55/fwZRrFWP8Xfm4p/v4Yz1QKm18k44EK2RbYiAAFGSUF9Zg101M4FnlxG
xdLSv32haCfAvd9rOp7n119mWOgpY8gYllr3uvO6ZHePctgBjl0Ulccj210/WpLfYeBVJikTirpX
NXah8ojsKpA0zi+xEghh3x92iUnxgKyx53QF479z2PvlsYGwpF5DLXV6SIntAqikeOfWmVzhV8fi
QsPRr8r++5XV2d2PpGRwjAfOx3HDhvfkce1lFShbuA0t3ZHgX82rYIq1m28dDsvxuaQ8nkioBpdJ
Cp/NX2qEQizdwTU3sgaqJqD2lCUm9vx3U4y2SfRNxEXC0V1Anqv7H+MPGRB+E2LlA9Cw5Oghd2TZ
AJGoAgbXNM/XozPw0MOCTy7RK6Jfsu9OVBIZgs3Xu/aw2JQ/V9r1DP/rgDgv2RX988+Fh0yNM3oA
1xgXcmyp6XhpnYNaOLFfL34tCYfrGTkcoMT27N3cUWaufMHBbaZ8M47JdcASshF++D8hHW1DjyXx
pfkCiHbMvwJmTjZTazMg/5Y2KgvXH7O79O4l2L27Wo/KUu2mJmgDWKV36bF5d9VJcT6PEkQPXz/o
uLLwfYWou19L8OjNVfyRM/Kw00qokW8hsLFh+TWpvf3CFYxX66kkHHuFS8HY3qDohL5AuMijjnO6
2FL6yh1ueFoBkIhtSSdTh3WU8kAuTCAfwKlu/C1lVQcbZOLapZUxRXOWpi9pQNMS2BFQBhkqatSJ
MhAibj6FFtLXFm3dnVODE5rFbD6/iA22k13aKgq68yv/8acWTMIzJaag8dH8kMZXts3dxcbsx8N1
3mEseMEm3/9DrAee//C+HA7MYU7FoGQAcSEd/pGQLBx0Vw6/B/OP9MYC+v6tn7Zf+M/04PC8AtcW
3TmUup6Ix9T9kXwJt8biPh9HxHuLT9maqIBA3JKJghE/9ayXGzaVkK1sHxwxs7TIRT4frdi2UR4l
0NBWQQqUtRjRFgCmVFW7YlNlNiIXJgVk+kBDmp9ETGM2zSpw+3MSyKzUs3jLCqkquinXFSnWB9Wu
l1ehuJHEAeKKga0PXl3a+Zr9D4k8rbjhb6p05j9n/LF9i96iVqPteKj8HXkJdpdo2odKQdQytcs4
qJO86hdk+fX0haVPWYJukVfwrY0AG/iq9LNVovQEF4BJLS/SjWcU7YvWuQHzVkz9VaWiX27qTCsD
qON4my5fRGiX6qMgovwNCbMojajZ2O8d7BJY6xVJGYhuy5nbul4LrAi3JI6l7jCKQPtlSBGx++KK
nrA9yeK7mnuKlv/mRHl4BePlXypfgtG33ZruEACaAhIiSCq68fdBMCr7C517pjgmK5paaTC2dHy4
FHgzDGUUOJZR08VJrqTruDZ9a8aDvnuuwMfHtG2fnqu4pOOESBAUMQyCjMf/QWADFJ2zS7MS7ytz
ht+xv8Xn0ew2h8KnaKbvbIZD340AREtuJpF4G4W6UGLU4Xx5mdMt6Tlvb1aoVZRFbmiEOusmya0S
PO72OVGHcEu9efdKeRePhbN1/VvkXHU+fEq9UFNWezSwmSQ58sD70OSCWkdB6+eenw6RiHR98rQi
nNoezbtrenYh9P0ewLp2HAJEgZ9qdbsNneK6hsebiY2DoAYVlEbZqzua9SkFcNyJPNbAQLxoqEAw
4R3nh1ohCm5R0cugsWn1+ZXB+ZdQgE7M/nxZ4ILL7OHHyaFE5jM67PFiOaKBaya3nONtRSCi5cuS
J6x43iurdZuyXy9JuaclJ8zAQMijNSuySUgXm7i7fkSVunZT/BZdSzi46s3s9AJVr4tfNCVrPaCG
L+DeoLEcfHMjm7HkKsmQ1WHXOCpOoS3B4TwkNfL31fbY8M1iGo0AJQdR3sqjsM4j2TUOPrsVScFP
UvzpFhedoT7P0VHAgmF8JN/lDE7HAdoSuBgluLS9zgY2+ZYeZbXpRhTBepPPJ8P0sfN8fZQULtUg
bB1N2CTefYbS8Am/j+S9LRBPiP3o5PWBPIpwjKR3uhKxYFR3QjCBIjfOqLfWazrfOvXAXPiq13ae
bRtZO7pwRIz+avYPeGMEm1P/bRLmzVaJwYJjsAKNx6EymCcV1Suqw15ZiSIuaN3KLnzV0e3abXMj
/vgM/l0Lpvt6cfo7lhkiY0dMRNCiRLlFNxBtv2+rRVcr3Q2QfQUIjIpwv1iDodq3ps0d5u36QMjW
W4uUFsg6zxdXVu1hzsIAjVl1OuPqRNO30QREtsZIzt5ofbza5nALDklyL8uDTUXzH/evDSUnBfet
mL0CcmCITBenFssLTjvy2dZFy5Km4xXKTD1ue00LiKGR8j+x5BrmGm5fczbniPs8L0Tno7kWAH++
d8HS1P8QxAiw3t1GAyhEg59lrNcYAqdvMkPNmMb0UzlDI04roewfr/FlLasUCTLIBpFtCGo7QBU2
mXs3fLwmWS0m/ZfubhmvGs8d8bKwt9afAGwK+Zh2jPKr1/03ffaBftVfS3tjXkcCoG0KernBnOYL
h2bc0KybW/2v82R5DzGa+fNc2gScleT48rmXzmXjmS4iLwKalQCPIwp9C33ctZRAtvWM7WRdReGU
tEbbA5AcXuy/fCjTfvgGT1vxCpwU56/xYo14sf5fRLSVH6yKCDsuG7T5qlpdykUjq5QioxtdbXiS
hZtcUzjJMdA7HFAI6VMAM8ZJ5GoCq3sE4KfSHPZcngVj8t8nlwFyI2yBscYH1EuyYyfUQ8Aycyek
1hoP4FF1dL5zmlgaJMBFAriPXj8NWTpRanTFRWtUjBcBjlk31deXCD9JJY5/WS2LoRBF14PB6T5E
HvT9N9qSKaPeer+KMFcf9Luf2FKn4hCgFHQNlPt+T/P3Se7Q1M9LqoNUnF2+LVk4g+z0YO3BESv8
NxVGYxAiR9srmrosFL7zqjllAriTo04raBENH1W5hA1KENOG4gN0qSUFuyzMVrAjEQRuFDQboRZW
aDxM7O8LO0NQg/Y0fcwMPtPoJX6WRCk5LkSNSI16SFGufFY8HiLm82gx83rn/4oPGE998VrLvl5T
lX0HumRQKBpxi2Solokwli7Kn7Lwe95tJF1hI1gaDr80G4DjVqFSnSwES1uaCA7yA9k3Egf6g2h6
CRtG42RNfu15PqBvhOSodi1+nb5N4Jd14LneKV0nswoRGuZof++3V29hRGG8zuEavyZV197xyajU
Nz0POs6zbt1VcZx5IZTFIC51AxFfiKrGo8oUNnAMZQFI5S8l0H2EEau3s9V/CHaifwU6kr2lIaG6
up50sHMw6Bj6xTgOisoDe6QJJsxOHY8VcE5g1tVOpwF2FdWcNjL9nU8vBk00Yz4T5UuQeDbKtUZ3
HycRcXqEp21qjB69VLmGZ45rqZ1FcsEvlS+edj9HnVciAaZQwraSnzZ1jlzBtE4suvitpzNhX4zL
lTeJ9CXCQhTeGGuw0VI8hwIy7GlfJl6KcCuFCfA3xG9Dyq0ySfYmgOsem0dEeUqQ3GlUgCf3wKpC
72321zQmSIRNhGvmLdpATIIEIJVlGic3ZqQdruvgOx9m3ziwgzozaKBB5XlJkTJxwFN6bn/+NT8X
WR2RfrEofM0rlibJHQdI98+aYIRZbTxDN0g6tK/DM2X2VBBU7SRIts4Lb0FBiswho7T7Yx76Kf2w
mdalj8OOCUrPVLNQU0Z1l0a2stnxusePYs44SPh5J+QF8jaH3I4ghCHkwI/hvX87pSzpvhge6IFv
KejC0KsKWXGy8kUUJnT/LwXhqq+X4rcY1PmEH17lQO49IcJ6WE8R554FiNiGLfiOstu5k+p0asU0
m7ufVLdKmdQpemGY+iVtJ0nKs+ko3+5Ayt5hgmbsLL4SKn5UtWHUtnlsf4QOKXRsfOuM590A+wwD
Hp01x/zGzyQJ+EpEKZ/GGyCJLpi+hpSfJWRsMJew3LGHRNP8ohHU2Bb3UBXZkldOeSho037R/18f
HKw4uZZDAbBwtbD6ZIZ5/TNsnRHuZUhWaDSTAxITJSp4lT6+xby1qkmurPej2bb4JMp24WOotjw4
GBFHF3UJGjOpj+hV4nKvdktvu6TOtspjD6FDV3kccrge8iEr77NL0Nl3G14Cm+ZMntHwBfABLm/E
ksOpnRXR3lbMkJXieM4exg9td1qHXAbyGYV7dt7BE12JuFXtocKKNr1Rjhf83SsNYMOgHqP/D7Ce
88sL4Y8q1dXUtP/DMADSb2E9CJkPkTGElm1aXaJKMkd1X7KrW/FZGMXu+qLU+dJCuLDwzYic94jA
YMVyzjtErsbqaRaD9xK07Hd7Xpl5r1NB3y8REHfr1Lub0v+IrLtlKKqXMnBRPaJLSr2TDZyvmgR8
7NU8rLicihwEj7yiWVA178CIU+J9Pp/CWRganiit/9iRRRdU895dO35d5CAZIa5zjhBEZhBVX5S7
bO7e2JOrCnHcP5K/484cOV/sVoOXryCuz0ez8wwXl7sHKUB+kHUf9OWs9O/7R42kwputqQrZIQ+f
Z2U2F/RCqe1ywmbF71BrMV4E3m87V9G/csUiBuiw82zPPZZqKwgXiT1RBCqXhBENxe1CwNDnP7A7
llOccZwxoGdJoLYrOlzwCFemFsxmxn+V3+1exC5xilOE5bYOk5eJK00I03njkngeGW1jjOstoTr4
JANzm5Kv9QdpL6R2sXutDIeABKsqtdDt8xphb3QyXb19gQynU4uKRT8TowGp+HzlvKM1PSUU+34w
2xpURrAgKQEB8HrVDXf2KRIdhVgPXHicIsKhyp8CSHct4NgNpRaIaCk8hQACpQqb0eNSMrbQ/mNH
Ugky9ps/qP8bR761uE3tJqmirv4zi467sRsgjB4orj7kc2WDTiL69NLQ2wTnpoxBcMngC0QHL5LC
2/bckMjLHvNJQlZuDuPAmK+uIpnd6ANpBcXUBrU2IzVaFk1GSZh/HtVc42v/GPx1MWGhYkxBDhY5
XK6pipgIcoc0tyRU6GrPKjH7zS1O7O6tZTm2bfkgT4k5mhNlbAaSAILNTpixpw8A4y76GWvMsQhz
Q7h0PKS+ItEGEbnBH63UgmunwwcB9Yei0CWUs403LF6XKRxD1zo2kQ+ElaOcOQx7XvwJGoOeLADc
A1RAuZ9ET+szwJ3MVqqlPsAhPxd5Gx72l61lfan8ec2T5wp2ACiuNy+mCIECuFWIjhJNZvp/VUP3
MEIxKb599zdFAJF7h5aNAQM2AvHJC5Tyd3fp6yUeR08Sg4yATJNJ9rQgDs23oFZw1Ilf3+WPar2h
EGQQQXz4BmkN7N5p54JkaDPoOQ6z1pXuJJu52YGRQXN/0b5ga1cf0s6p1h0LgwuXJ3AftMb1lr7G
JqQtaMNYwVD5ZXU3sp+Aapk3Oh2OsjJGORi8m5A464h7s2x7UAfDtdY5vMXcuq4Z/N1Q72vkc6FQ
zujrj+hketITprNe8MYxlLl0z+ZO61fXF12815I6oKJzVB8JdV4UBH2yJIhVPdkv1FA7wsDOxYdp
oms/7OEQEndM9r1OTcUOkxLjVSqmcYCJZSQaNTeBPyHk6pNTP19hxxsJDUs9fZtNkIgyYmImo/qz
+8Pgk7qAKsn0k5kotPedLj85U+pA81fMEL2Yxcm32GlTBr6ePGR3Ml9IwR+fULIyNBPT1ldCgoZu
HBEeS1gOrpSjKuv3Ul4l7xDdyQLCcPyOHJe93yXdwNomse/jLJAMpxz5Z1x6r2tlhEAq43Jx4OTb
llOQh3jhof35RDHGItw0muatQqJUg+wSo83HBc0x3rbWkvU4ayCu5qHUw8ODExFHJVnDKczN0cFz
R/0GHioklh7cJkM+uQWU6mfY8gyAO1Vt1bMwwo1pDEXvYEg63w1cV56PjqM8bs1xdkMdBmdm4L4N
AlxzNNEW+h6Fvf08ZImTKukxEUpub0V9L1EDAxEiwiioMMzd40DSH2Fub46caWvAIFnwzpMWGRG7
Il6dxbGDB97HoVEhWf0g1md9m4HzjqYU6OhBt13jby0IpeDIyhb0Ce/ISd9sno3ZCVuhS1V9kTfq
eLaVUK1dN2hXYlGRS8IPqXs5HZTTV8yrDsMAMFSBsobbXW5Ja0y+5Z7yVbQvWzsQeY5UIjBZZ8nB
JtiANeYVt7HjQHmpWwErnXRxHDk75Ep/fgDYMEf9lABL9W7lcNjswWN3w6Z/4JACe/zndTr0ZF5r
WZHnECV8Wn0bIddeqWiEpMCxq7HfjDv7S0Nk3JNdQysZDAC1VwjNeDqbW84n/wQWohmMujl5UQgK
h1qZUDKQQvVnSaCKanqYe2LAvHrSQT0KIyRWNhlWdQgMovejD7iwYmg0F/1h5hSWg0DogNSMeObl
pd/0a1CEXxKFMnaZL4BXtWaRWdGPbEBvJ6XLs2y7JWvq/bn31IBmI6d9NEe10vJpx3nlm/prEd4J
0VgMbB7ezy/jIleCsCkOC1xhQ8zxb4cdVayjtF/+gjP8IcFQNXig4AguwutT4pAu2x4bDUCJo/7x
3DHGM45PNW8gays+F8/8m9XsGffMxtw/60tT0HxDC3KrN0dxsDKYMeh6Js2Sw0ZIGp7mR6cDuCNO
hczA7DEzLroaB7k/duy0ITjUs8AndddmARZ6Fu1phqt+2wkpjX/+os6QDUs9Vk+F4fZZ60WgyJKK
sTthRZ2EfEIekcCUJGPJh/r4vnDJQoGGr/tOeYiehMGTmuZ11z8HrrPymUBQE+TJ2brNEm9ystRa
TaX9GDdkg1K+Mm+80CJt+ajV72eAw2w/tV1Inb8mv6JdxwXju0Ho4cm5z6CEP044NCL5gEGn0rEd
hYtAH/vaCTRv2yqmlghM8ztIhLud4FTt3BwBBYp2LLBXvd/MaUrQAo/22f5l5AG6aVJt6GqHB8YR
k43uU2wugbQw8l7gzjIgzE8JUwZxUecgTGimw11IDEbjqMMp9dlESINbwcjk23MbnWdpgQa81IV7
HHGyQbL1+xy+A5ZZ19KgJbEIyd+GHUawlNp24bYRPX4S76t8aNAbdyH3prlb0rxlEETXi/LsStrn
acmhkUaH+ELAmpJcCpTzotTGlTMqsfMbR5NTbGCRjxXqxclWTd7ewQQEwvsKn0pFP71BUC25R4S+
CrL3ezI37MrEBeY5iyVAz9+2IQ9GqbSEfdBDvDyPCaFh43sanc7r0pGH5pBxYhTCtdwKIjhJjSrk
JLZOQXJ+bn6hv9gb4QOYVrP0yQHnIFdEZNkK8ZjO7/anF01ZjSbp84jnQZbch4Sv7dUZV7rgln9h
mNLMHpY4KViqQepRWcaK+YmYK+M901Kp97N86j+4Y5WqJwvTacguNWy2tkIWe0FQTZnseolkT5hM
j8hDaY01TG7aZ/FhZJGUyWDkAo3V45WQQBcr7/6tUgoS5pk2TAW2ZAEO/SWflx+7OzrnBKeHqoZ7
px6jqMKcOY5tt7BUP42bzXYNpIofv8PdO0rK3PlOd6BxlHGT6ADLY97zHVv/QiyjrhygOnLuo4TG
nKSL8V987c4Yerpupu6t6RbjycTvbKa1OzYSXCYJnQ2sf9HtRFXrMt0um9XGbcVeAR8yrluZhWJp
nPF43Iqw6sYhw5aae0fPvZWEi+cXGj0/fMvJNs5lE1e5qhmTN/E59EWGaiqnhZQ9v8z9UmCsuaxi
q49Omk0d50oIQjc86iTF1fcLYMrQtuiUjaFwwObHS/nZT6Fsfu+xdwPuFLfaAaZLvZva6/wuBp4y
0EdYegTWJYlbnOgwXhS07KuMliSiJJXGrTj47lFgSfk/U7HyuyT3WKsXx20M6cDQic2E+PvX+NVv
I4pdo+Gk67L3qHI526dBJxrfRyxvshvA+LwqEUYgdxLAdCAimgiWOrsGjz8XDGPryX7Y/yW+qaj8
0YbHQwgVVQi1gdtAb1jDNJkKbmznx4LDtuDpqSfI3yxh5HwdTjfuYz9ZtpWh2L08psPPCxndEDRL
UdOxkWxfPsf6pVTXwWzux/ZyksNmWfdFFqQ1icjOVLnlxlfLA1aAQSBdgDpC28oFrzoWjs2uYzSn
vSpk778e0jpveWObC3Gzi4lYv5vK8JBQWxc9jvilnVYL7ezVvavGqm5PEnIYLkewinqaGQK5QVu4
AkIuggJRMsbT3Z8fyztFRcH7zIxOsDCNrzk59LlTlA32VdY+GMVE6K2RRibT5CHKPz345DRwhx/3
RvjGSwdRbQ9OiPV50y9YdRinNK8Mf3QK8Lq05oOGr9Py8LKiTj6EtYeIUeTP/OGT1qIrPg6IumHO
OgtJ3GNuPlDCg605CXmMuTdYXAWedF0IdTnSyHJ64JRLudIdc7NCo0bfvBkakXCWenWaKgquu7d3
/uOBAGE3rTo5GrFhNCdLi9U5Cwg6sDCHp6wSZvl4B+LkzgygbENRWckHOAmut01FL1YpytxmXP2c
9bypoz3v5CQOONDJVG9em8MHivRvW2+hOHJstgtg5L48CKQLTN7N0Fb9a/my5M+VtwaW1FE3u6XF
GlplkyZi42O0jnZafvSB7Rs5qT+qzZQtWAK8tharzP2nCYxAgxpsXvX8z91ATzRIV3HrerMlzZVU
ZJmhAKbNx8ZsFQO5DqEbkqviYvN0/BOXje8VcTFMZqHYs0lEIZqLPwg4Fy2Ihulx5CjwBe3Qk30T
6qinQK+WWqYXA7BTuMHzd8aSsiQIvwbnLVHPu5WXk64f+VMMlaa+Gu/A4INnmG4gXsrSNO0670WA
JBu+ATRPtsJgfwP7AXGYJa9iWZBOnSSRjAScP9v4UjePyPnKaqP2AgE6MJghEvbJLxTmJmn43Lyu
ka2NxxCUrBLbgrOGxYW7fL7RNjUOl3GPYwfNCeR+SzIXwHko2DH4y7YLJIFX0CmOR64AVuh293/Z
7NPZx2HFv1wcd8YEeJi3y8G2hD89sN8ou0gH8xXfYkWdO3yE9LUJEjyNtCuSaqKF+ea0gDhhfm6a
1yAyKgD4eamWG+IB4xOy4HRi1exBdrjuN3b+zWPOtlW28b8ss8c+7qnju7ZXUtFeKzNmdplO85fu
XXbIzqbv8+vUBytX8DWaarcpvKv327l8rWhmzY+ZI2rHZ4Bz7YxEHadg2kr46+THd4HVURmrSKWx
DzsrYCNZeYVvIxCt99mJERjDBPLtrKPImUR3te1KPV/hgexURmsvZtYM33jJruTAPO9tYYOz645P
B6MfeSFHehm6E/NsQH7b+OKigwMQ+3002RwV+wLSie1LfEwvAdzPLAeSGKrtvuyTACY4B8QtF46R
UpQl8dxWjmjhzqpnfHzbaTaKCbKQyerKo33FTdYVXB+vhfR6EO2MCnRLc4+pOk+zrX1vrlYpEkts
66lpyVk88C3V4cIhdOV+4EL1WcVdfPrT4ncVVYXl7jdWEblN5YiQ+jDau/9wAEOut8wZd4RSHyP/
bRw1IQIdggXUlD7KnyVq9wq1TPU32vrbBPZQ8PGUbzubdY0vJbhAi6k5YKHjLVI9bKYYhf4EFqxR
/LyPQr9EUgpRXdnjVefI9ytsHZIX+j/nzeI8810lD9XkWElEwOb6/wS/EYsVov7okbk+m0kKl2Pe
cfVRmlmpW/TtwfLwirr6jEN1ynZ/Cr0RPcJDIQakd2NcueeH6oCkgwZL4WvnHn0HiWeH5GRrK+JH
TWEN9cWPfQWXE/CB/RT4T16eQEk8LXb2oNJf4XsDAmAUwGG0EeXNlcM5JHnfcP+lm7IyZLOGaCkg
87o4hrX5EHlHner9gpRfYS86bBspAa7TSZWb6allTKJCIk6BV+jQ6oFxG3VCX1tggqRlJPxKb0z8
4YBWkpz4PVEFandk2b2VKJYReiAaoUEiMUvz/5Q6bmLu37rC92bNxrDWdmDP26vdl2syMp3cSm2w
GQjvkbeode9mib0DI/e2Grf5BnpTnEn8sfwgKPLlbG2PDxFmWCdrMy9dBN7tOtJrtSrXyfxN26Z+
/SgGx20JI7mwRQrD6rNkAdkvnHTRoXRcECJqQcTMEr2VTSfy3m6c9wjuVhkRATUJ2rg8HdiYpSuz
s8fI33LOpuLrZ32+Y/qu5HyRAEPgEgmYgFpogzSLcws4ca5tii77TzkIb61eTgBMtasQuPgqIQiD
FzfG4fLSxUIaehxzkjbrBztJddLtlRLHWWde1bEC3D4Bnrx4/qY+tzVZUq1y4Zw6CyijOPJ69/rR
IQzQ1ziWb+qbg70TU2rZeILfKMpzhX56cO9ByPKmtbf0ULQec893klF2FzAFtC4IhjFYdQTh6ziZ
ebo4akoNLWuUJnfNQU5AjddHALeC26jocL9Lv3T4s0qknVbjjw7pLswQXjcypdcn1ji4vUw/T7ff
RjuP87w0RA2HXCAEXRv4CL4T8Gr0Y4nLru6NaKOcwLzPEV1G8UdLT7SMiD8IAA4sptFNBsT63/rj
J8ddk+oO3mZU2B2Tl/hOveowB4niEDjl6byTakDkbNuDULtUQC0G5zoFQ1R3nkmrnqlwRjwHp4Pp
VCseGj9h9Dzkk3R7DTVX25e89DghS2+JBXXMAWXJ0aTnEou71oiq5k8LCNZ0hfDe7juVxKpDMMYQ
9p9evSAC5yAJXD5/xrcFv8izSce4vOJTO8kLrZiC4w9+FxI8kOy+9dJTQqDC7TPiGu3sU7D7s3MV
zGsXj76F5hpSrQtXCuk3IPZyinmS+d1zUDDAbiHDAQmde1VARry540l/kjFkQba387U6enhU5X07
x4gCFOineqrjsmloMDtkwJhy67KZMy2inxZdphQVyzviHykgqSwf7vP6kJtuOF1juF8reVZ0gpy9
bDAowLA9LkqWcRxhrzfV0rDuxZ8h+I5HpC8WEq2YhCvrWyI1efqoljFr/HKrG0DZ67Mucdbx+0/Z
aPdbzFEfxL52VtzJNf9INN4dkUYZ/rBgwetclyXLbmGQmYZGcaX+856o7sikq9QCFr7j/kWhfW00
KvD7Ixv+0IMYTXV5cogTElQRJ/PtxyhAe4qjgaUmQPW4GZBBRAtGBjl4CJ1xRNsZHU0wKjmO5bR9
x5o1gRQOOb+wACEL9+SRaAEcSC/aMyOKYzO41K+s0t7tOgoGrMelFpX7lfDxVnFigEG4RZwJe4GR
/pXxqJZWEMxT4Ua0X4vk5O7H6Rn7teAdHBfKZqmEmwJV+eew9LYJpjyBNIc32TXjUCh+RrlP2jQm
ff+fi84wUrhPh6NaPibcGa6b/vA98jK7Svz8liHCorLlzddabuZMfXN7n48ga/aBH/KNMDFolhQC
RIdVDU8UhmkuadUms8cP7ifpwTY8ZKrJn20KnaACjTFBhU6CwpzJMfVSq/SDD8LqxZM8t8ChTRsn
ooCw+10CSkkWIPfj5H+LhY05+yKW6BrUbamT1HjjneT//ao4e6WuWWtliJfuL4VlGHhV+Tw0F7dt
Llt2kn1ZM0PjE01N6nXxPwWSegOW+CKSWcP+3s1AXesRkmTD+qfncrQ5p4jCVfE7pKaZIagwWHi1
HzZ5F62DVzzrVCeopXJOwojQQ0YMVrLggusDv6P30NkaBW/tulBDP+cHK+s+GU5se9z7RgqA870F
mTZkuRhpRWnACrZvi77hey4DFaPgBsvDlD3iUJD6GCMY/1S2UADIAhhbm6mmmEewTmCQbmSsFpLe
aWMt7mxenvMYQxJOaUVxVY9Thq7ZoABt94Rl25CL4wEHJXrbvn4GUZMIK9JSNFTRJwpBHQINnwur
/neEakASmxL1WoPLy7Z1UN9g/j69esxxIDsG2XC+YZBSVzg9FPYzk9YcBtusJhL6jOiV2uKvurQ6
vYBHMqF3vE+QyoBVlFd8qGmYnF+8iJdolVklam2wTJToDHwVrja11W3xuqTspWsOW9n80xawym2m
XMcxAzVkYlzAbm2VtUwyEnjApMY/d1oIrlaNSehoGlIZeoS5ghWiVDBvkix6xWQaw2wEUhROelW5
BRZ8c11M3IjYRrlUt/3KObSUUCEfqNMtVOK90T8oeTTHoDNn73qIEpoLC/mU23Juo1vaoMahj6+Y
1vG3nSXQ50wgaUVTc4veIjeDgkBPCsiNFMN6Qiqs0ECkpJlcrIBEV4xK/BCuoeyUOQFxmI7zNbJd
VUj/Xli9dSJ5eNu04SybJnsOcs5dsOt2YiuIhHf+6z7ARoYs623Ve0PTeNPAYYxxjPMyrFOq25ST
Og5tuONjhVadahMkhzdySGqWaMWX3igW7F2fXbjbtpr9n7l5MnvNemhh61JTXg/eYkAkxPb2INat
jfwvk4vD+frJjDJk2SHOqbD3tBLox0djRjnS/7opLWah3nm6a0buUiCmxF8+ELxeOsdEaTkjYaru
uF2Vh4JE882FYWZE2EjDu3WmkapWIbj7DstThubYLUGcefvFyCyqhV/YIDHEHTC6S4Zhj2Mqm9yH
lqR7YXKf6iHW2kr7fhwk/sT3N6tKd36zUKv7H9PtOXMXRoGrHyQQiZDPFGryDmYD1MZWfX736RGX
3A06B/ewI1tTXxxu8/cm1xtoo27RpbfpgY2LY7a/JEWqHKlk1bKT038hlWQPT1pTTiuED95/g/lt
MUwd3J2FitjDtMgtga7/MwOPnBlejjfqLUZZQLjnuJqDoRduI8uJWube3CWFMM4cGtoDpJSSMIGz
b/BPI8RGBDiIZ6mX6eUVbcFtlsBnEEuh7GBAdmkQW125NR0x8WSWSts9VxCV17bhBUeDdXrvjOSd
Bs/+s77F6YbYok7e0My5JFRqkbW4iFZH2nfh6UnnLb94mhPNQwgGwVZaRmyPrY2V5BnRU/Ta/i8i
rojZ9DFaqSoxSJpk2LzxcdfCzNJhRhT4ZmUM9ZMj0XTOQX3qyDUfLUuFJtKiRqPvYVslvby2IrMG
lK9jJ+A3HNls4/RFpz4GaT6FhtRm+dUcIZXdyN72dljcYYbtAvc4Uyjs0a8fJbqt5GeN2LBg5VH0
yfcQAXqY93aVCHQ/J0Qk87PbrF5SPoHAy54mNQ+SaF23f4gs73Al8JFSDRVFl7fe9B6GTTsErADI
JmycaOh2jQpV+jTkL8LgRw2F5SAj7lve4xFfLnMBuQdSGOGgk7HLF2kZZsn6Vryxmdh9doCBzqdS
Y1eiEbkgd4fMzKuzuN/aBtf24Rv6/IqD+bhKS5a++WWf2Sb+OII7LbUYfTtyrD4sr5m/QOt3xIxO
GfmPtuRuq5sNK7jNouBrCCJB3N5akQoS/0Ah85D92BSFQI3HrW/AbjtEaV8hcCPsM0rL3R7ClDcR
Rs6N5syWLbkbCli3bcTZ3/sAyDsVCXlmRhRwLr3y8syNNNsDJILLIj8J8nKLxCkFGiAUAK+do5D3
zulK3D/ftAeFMeH9goUDuHfvC35Pd3c5KLgFfRFU3KNkRzJaBW+n48RbuO9gjnY590EKGoxOVD/v
FbbYXvYd9wRf1dDBmiAzMDCNyL7VZbnHOR3ZHMDZTkIEcFK0oq2sCu5qzCUpPfUltZXVZH/SPkMG
g2SyC3XiVroVWYGgux0rBO2C1ATrSgNxIgUOX0Tq/kFk+wrL2skYMEQ1tm5dMM+v+/MWX67mc0f8
i00ginlaT4zM4+OTeivJdptV+0Q2qMYZHCAf/HO2a0i05d2lf5DgU0jIddS8EUZhOl8/DMOd1iTK
eGnV5FF2bynufiMcPEW19Fmg4EnEzXK9aR/2Cg1TsCQqrPCunCeB3pNWHnvjb2KXNRhC1Fq+xTTA
+U4jnUgKpMm1Yg8G9lcwsde+pqggAIa0h4mEzoXRfGk9kI/sn3FQhAa9+OwLaMfEC1tOYSIXNktz
MxOinsICIHXZIahvWAIYvd99FhDWoSfJAVCSOVY4Omp4DWsNJ3CGDIb+OIz55J0evfhm+EVWIXtC
uGEeK3LyHMdEsYGyQrzvzJHlajFx3M6kxtS7GY73XlRceJ0sdGMa9U7o2TaSUtmqRCMtwARacZEN
j/VOviqtki+Kz8QjHli5PRT712RuPGVa5XeN4F9JRSf2Nk2eJq93pHQpJlT0tH4dm5et/fMb4lry
rwHJ3cRZC/rqGPfcaxonWTK1ZkqkNtYWC4H1AZ03gU4begur5weAzGg61ipMtJkKoMODRSCNxjeV
/ODha41+M3Vt1op6Mh/eHssSJvWCmbHLM0/HL3+E9Rn9U9U36mcw/JYaMIqlWPkFkkxpCwrZCDuV
5ap6Xyh/4gif0M2onRtfC7tTGdvke6MGwQjfHRDbxKg0aPErZFj3GaL8dT9WcubwXlMlWlLXfiYN
Kb31yAr6ST8ImO0yfoAEDGCQGHP6RF01DwCo7ftOilvIqA0IeKpvToKdVy/ZpdyO4ouwycUQuXTH
GnEQw3MO7Rb6yFX1rwk9zdCVAifcqovFrq528PaunPHba02eN8cmqxzxuRKlOidxUQL+jPWs8yaV
uoo8THnG+sLx6IuVtUaZNIL9XUoqkvqBCarAcpI1o9oUthtfH10zWrh/PDk/nuMDHbzZsglrdJno
K2h23qt6sMvQps4k2kyY4GfWE4Xec5Wi7169rjLn+11pcF6H/sn9BX6d4datWXQfP7SoPHDuKdVN
jogzYF/fU7xizR7EcHUwu/4XXRcH8WFUTn6Gb3KMlhjwWdLwFTeysYO1o6gB2JRcm+OhgQgX2YSP
9T51PYgXDE0/8BRqNjMOm3cOhkCH5RSJUXOlHDcHBQyLmvrjXzXTt4oXIHjzK02HrQMCfkns8YXA
L3WIeQ/iIuBgi4OUv87tcCF04fNY4QfC0z8S3j07pt+WhKio2s74vi3NnKxonaTACcPCU/uirblR
+nBahzObuYJN9xOPCl/D+th5rxkiw3yoFjRi16uM8UKbpCZI8uCMexl7LdUM67l6VMnsvI+278CT
2EUqL5uO8sBocERTgFjXqa99UFaiWaOkebVszL4uIDHckyKRvUgtRSiXyfQGmdg/ipsAr1QvwFvB
Lq/w7XEzeBZNDLjKFELTw9LNI8hJDOLXEwdMpTFeP7E27ah3KHwH+JvE+v7lPvWtsp1X+gydG4fr
hJ+1b6hRAinsk6jFHsoCwRMpoLZioyBEK5Zn8/Kr4jbFW0qtHn4LTLZXHI8io2CYkdl9ByfYjSUN
u0iKYUkeuqRKPVQypQp0fFiEsOEd06jHQoT2S31/fs6byt2AWx6nzj2qJB2ABdpZQjdEMu3p+SzE
JLdszRUg0ns0Ggcbgkmh3zqTlLzcsGxQxPQCEvJtPJZDy6ftSphf7RM6p3/yPUNlIQ6zvQjRxAPH
Cw7YjqkqhfFtDgGZ7EozLjsloQYGYqosILfW9AC+C7ewumu9JUc7sByxPiKisDeujq8I8KnrThnp
FZ0NPlliEI8FS/RQOPt6uLVQs7D39kBSQYSv2KvNJfSNhK/vHdLA+rAZhoG9QYrctMWBQO8Ndv1r
IdnrsK9zMQJm4HEcYnwZ/svMvTPsXS+YtKUOWrdu7L+L2om1NQGC4rHqi9+TROwO/1gdf52wVQm/
4q7oIEh1NA7tzA78Qo2XCIEv4VFodBFYDOUSYqtwzJ9rkwLfgaVQFnPf7efJkp33+FwoNpZ88OJ7
pfLP/qzjjLEKA2B6+kuSrnDAOYlIDKC9oFujvbyuYfWEm4cB1I5WhnzGeyw7N1Rn8GaIviqpMesO
iQO/iUTlxCa2r9IuVM+NwbrAzU3h2akba3o5Mafh9nvhl6JRfHUWIGRuWTM+EjsPexXIzsPnYP6N
7a9uxlDw26hQl7fX5BFR6tIPH5LqkQEyGI5LeD4QSj6HofNWvQo6mrcRNrGLU8b0CqLWFgLCJu2M
65sIjaWzEdo3qG5dCYhAl2R2K+U+fTL23lE00MHZiEkKZRpNULIEXIk/PKeRMbmb1W7NILAFYAjN
EZqECWJbpGCWHO2u8za5hM2ARmgVgWpqKv0d6cIYwLz2Jab/0DFsu5IzmtaiwSL5Tz7QmTQJY/cD
V/J3TXfsmlRdJXTULNoaFhZ2Xol9lCtP96PD0CCuVPgUEv5FPu8mvRlDPifoSk/uym6PrVs/+Oe1
S9uZj2rAy9b/PPEtkeO99wwTzyT+AVtIC3jFkIyEZdpeMS2cqBTdTWtb4T2TUkuKvkh6x70TjEoD
md55DJy0vb+ZSrxnRGLaNQ5Of3A1ktCLs8qh6BAx8rgXICI+sIELuMWzZ9liPDbgG3y8tSB7YfZh
7lLpmZgkGYxA9QgtKCTt1z1mMapliccnPizSZVbXZDOdR+r209PVAyAMzIkIDm7x+57Rp3HZonm5
J4blJdHy+NDYfJbz4lCHIXnOS532VWmUCuanIXyVNggB6VMSVUyQ7y4BSQx1HMERRZFwe6CtvZBT
G06XCxlyzQz1UYNomKUMCW34vDvmysMjOcUZ7HCdv7Gg0rJ6BoofDggIpDb6GvglUgf5heuWXqP9
T8GyvWZczKhOlc2Q6rhFA4u9ourEjNPswFsWtrez57q26ch7JIOKSk7E+/QJHN/UtR7EZtJq+jL0
dXHFOjLk4FM3wkvHMfWfPwXK3+SqZsWzcuKkV0+KlNS97QmmQufm9OFfPjKKkKHF/sRdQq3YbJuV
GcTt6Z2UdgQQvHrt5pV8eJ4aFYYrMr817h8Zv8Ek0kcw+68R9mWwTQa6zKCHLyxmLQPikRIcClc2
Zx4egdQLv82/QIw/cmOcLGkRUqyLmzFL7mbjMFW0ofQpwhZu8Z5YKJ3c0t7qKgrIO9pUASSrHEv2
LgUVWA7POXcqSCeIXeSeXIxayHT2dWmuxlXgKPbvE/ScuEp3CaUGRt4SuJwsAF/bm9bTCSUBX5GM
CW2eQIkOa1ll/xcOiQy2/b3a5Mcapn74ZbAIK0F/EE+DbVnINI2tDh4Hpa71VMEFinbrUOaqcHfw
FpKZ0b7qmFzQsltpMod9m+HxBBpZG32Bw4C4rvHivrw6tlMdf42WSxI7ruYDD2+UDpJebz5jpoLe
bOqfb1VBttc5Y1vNTnypE32TdWtzxBeh2R41nyQHyqBvbcMre4fj1wNL9Hs3DYKlZjpRCzZeYb1Z
0gVsl+3gHNIj8MIZau0c85CQDJvsvS4h5+Fhk6zgou48aT1n2t2yUmkAR+p/yeagO3mPZNnA1JLo
SGL16hICHLYarRV1f3qa4a8QGHLvjIfS44bN0CuyzIWy3oUPKpj7SBJj3b7pSUoHZUzAD+24j9pj
+bBbz+Nal3cddMVZAKnOFaCje2Ne17hnWIkbVY4c5McCJUUoTQZTEDapSX/HsOUWjDbgrEeLVqYD
eZ+QIeI0YLvqNRsLgGgbPAZ1Cx2DjA2iF+P/qoyHfYV7pFEyewP3E1qMq8v8dJU2F15nyA5r3CNU
O8mwKPzYpSaEkWpSrXhLaLWS6LgUPdLFIzjPWamMcMR3+8fyKfqQN6viv6rvGyYQA+r+fknsHi95
ELnDK+ZPyjtn0saqDa35XvjH+cP06Zg4/o4VKmv/evGksl0RE6jEMBaMAelFtmfM53W7l6R8EZA9
7/fREwTOEpT84PmiCY7kc24kaZYbICe+cDVCBlzpM4XIA6AD+v8K+09fz9Txn2hQGzpCrUtfqj+i
ExhYmzosRRBkDlMOpgYvO4fPQMZ+NPSRyW1WHmQDdFrWzpikf7QRNglUwHfQkFPmvWQpIerhV3qK
qcr1xf6yG4HX+PjmQ8jhFPrxXAUD5bXzFP2YBsf23kbcWmfQyYvJ1AEI51CdoJEA9zsMHE2dutiT
nsf4GIRj56rGAq171b60xjFrUZVi0+mbQnCAgNjvDhU+3BRay0PNCzUrivRLId59xjF5m62n0qgP
lSOpp/wPfvgjEsWujoYR6m4SFS1zuq6XOYK+aGvRKB4FDYPcUBZDE75f5jANGmKfnEWtvIkHQmSx
BuWLSHejkpgTXwBAkw+SwkH5yu7Lk58jIWd6jc3noqOuRtQR+tJY6sxWBi2EUQD7D2c+LwDUCeuI
3PNGYxUL7pN3BQBbeJitgFfyQmWIF1XtWDKNzk9nKJr22unHiWLCTx0dPIzhWAiqfUER7yev5/cd
Ybq0pTdztAiyYwL/BpFXQ/zbRXgd5RlwPYagFkqUJFYKJv26I0Eq+V9FdxMnPk+MATBG5ojGYphg
l44jywrZd31tPHfbSb+EFpYj5pfFIhndA5nYZjdCQwNNZVu4G71CwrIMI+6JHMMbco8yUY3zLP2/
rZdSGrI5X4yIT1U0bPwTirwzXXNrepey3KMzfb6CyZqg2AKGdq5WZM7gj54VvWAPFcx98Yt/FxQ8
CkMETB2E7ZnxZtiA7ymP4RcvYVNVqnyj1hmULcgcoL6Ig4l9OIKDBxs2gBuAvvSlfGO/PfvURdX+
7NZReNwbsGGXcLbhj0obmzM09N78nw68oiG/J6bm+XNBvvUsTPw7mHrOZ/B2CgdS6jbUclUPOwcX
PYKxgTtQFh84rHWpXKe9hYRXqqguHRKy7K1mZhC8vQxDuFVv+0MOraonaFpcCm7NhNjGTa25jXP6
ErykqDC79IgH5JqsgTP1nxWcvv2C0NMdKwuxsXWRh4ZbXZ498g3d9zu1Nd/CTruACHUY+KaIA3We
nIDvc6+VbqmvC3py69yZPaSYm4TAGqY/gES3Tq1Cu1xNOkN0y/rCt8Tw24F2V9xgp7Si1uDrOnI4
lDDB7bjYHyICOtmJ9dzBu0fbJjLJY8ch4H/cuvlEF+H797Li/celSJlC7pZfEPmLo1Mbdddd8Wsc
loNYOU+KyNOE9pAWVKf3AxHtsgHR7DGxSIc2d8Yb9Jqj33a8gNxNEsWyEmjn6tHBywRxHm7fIOnX
QTmXU0fSWEUAdJx3aWfa2ld4Iy5466l0/RUD3fsbG4xNcLHv2zSFErTJzO+d6Z9b9GrtjM/RiE25
2/t7yMZatWcc/Wyui7IsRx+Fzz/kEBc2zoEbXIsV6fdp+5ZBHZjntnsnVZUtO2/MIY84OBrsYtG3
R6DypFG5RbNKNXnbZmEDlEOUsa1qneHIeMGsTWnFJHkDjFkrTYPE86jrHXzcCScobN8MY5YTbD2a
ksFU/BmyIkOZo7jDhTRnFMpd113+5DS6ECVCmEZlzGXwz3NlLJEa8pgdHhtvRTJPFCBDoJVQyMEe
YQZwBx65mRME6sFeQix8KdpY6nGSK0dtyeigDaGSGKwUbkAhBd8k5b+ZLniEIvUgBu15tfvAKh4M
yOYp60GkBQ+tpsXcYf6ggZxtK3GEisc6BgW/5gTFpGhHGREIrrKCKHjebb7LDXEFTAsPpqsVRTBz
JPbDKIE96CeYjcHph250FsStpeUjENhlHk8oIeQ5B0eEEsLZIV99eG1sJVH2r/QdOXCMAxKg2rBR
EH1Gq+at1QscRp7r3bzutnuCMl+Gzf8WG8pd3Cixlb1nnVIOCFKPyQrIA9iXgl3+ilsV+EDXkQ80
A4fW1wpMkyHmVsiR+m+uw3wgKmckHm4BlMCRU4Ve+nyU8i+NCaGzsxJw0iy+rzUdqRO7BW4csG57
K7pbV1yx6iLhYCOczAd0hIUtQX4t8t7G6kg0NxGjvpC9bejMuVAWj8W/BZ2Bqn9t7ornKmSK6AZr
IOQo3W1GQt2mXgxk5OLW2TMWCKiMLzYhCQASdr7pco7sUdddUJHItXaNrP/LpjnoBTk8BVEIuuH/
CTS8tM0pSSXEQPfMX+Twd8dhZEE1Wj9eK0WGJIhVqI8nGUqxkQBk1AV9ggd6dDdM0giWw2LnDaaY
TBUcN3tcQhrqUtB9hXxqkoQyEBHw5HjvgP/bFtXP/aGYf+xsQ4Tcw1vwuHsU3fVRodP0MbGOi9TB
mL7iJ5yPgOlCDlsm2ivL9xpl+O95SStpXt3iy8tXEY5vPsnAoMzNWXTO01R6SQgvHMTZoYi1Xjec
zFKyEbmttEoVB/iUMRBYHeM+lWemUHnxnOz83gHM+rAF9DZct1up6JZYVOoLq239naobnVXfdZv8
keuGrPbhPopzUnYmdHFfgKhh0V19atmtBpTBBvqsEFAhfkNsZ8xjf3jOWEDq0YzxY14CBb3PSC1T
zZtJDmlrW+cpAxCDrZbYxBJeeR0eMMEL/dI4tl9RSfUl8zrH0UkBYqSyI+Qy7X5uQyb7qHjAehh5
rXYqubLbWAsxeywg98ffb7cOok1quP1ULlhQ9MNSMHJcpf3uWV4ZfA8d++bfMeesbOBnDU3sB6ma
syAB2C69vsGI7OfLu09NErCsSd/hJDwVD1oZ0Hp8noiOfDKnlcC52ia1Iv09jvXhRj0v7mtd7V6K
VyivubGpIy3pBTrThHC/Nmwg6IxNyfwnDIRWvlkqjgXAIjgOjQNB+UFFFSuPyLVDLa6A5kay6NeL
Q3e8Gv7GtZ8t0JoQJKoez5H1wfYfnqFyQuas7f6rgYLYZZsNm+k1t1x9cOKuQZ7hEFaKMXh7tZCg
iCKwkwK1K2efqVDi1WGLQHG5kon0cy4hQkOJSdgA6c6ltnu4SCYoQkPLfT3/Pa+vSWpj0L7u2Jyl
MO0YVirY8rZW1dhIPrVxkdRmm6eskhpmbNxlFeWY1ksLgA5l1BpUEx0fhERMbDwNUlsSn1oNatCg
C+XpVv53JUtNyJc5XAK5A0DVfXmTY1A3j65/TUtkryBMH6g1kMbwWbkY5A0iVdC4Xel0pcnehjHF
6de2Da07WwobrKNnq8bWyKXksxeyfy/ImJ/hSeupJ3ftv3t3o3dvf00E90KatSmlEVaiBOnKWyYK
3Bsot/OV6q2NmcU4qDxk51Ami5451n2VN4RIv1fvAMoWTlA2DfjCT3fzmo4JuPgw1m0jXZDOD/I0
0Kla7bQTWuUQ8SIkGVJzfUsw9etRxFY/s0H6uCDC81SmqIWWvc5VA66vqbpaVlpS0sD7ZTLC8rVz
gKLrsdnNjz73FAXxA4wuVp/KdUj6IBR4JjsIrlcU83HPCu5iDKCoJ8nPWoKwma9B+L66hVfpZyWm
bC2FHflo628Kdu1m9Ov807eXTxRQvFQ1fhQAza3Yn6JXqR+pyWHy3jcLOodhyJl7oNohBg6aw6XA
D3I/FZcNUJrsQzVEQG/nqnKBLQxWqAAyWRW+NlAznCRZMG0XzBzfcLExRysiZq3mhxJq87WxkWeP
30jM24JXckbFIFDC3HcfFL1Bp6ktrxC0DWGImjT+C8D+w9QQjnG5cMSWOWMdYg2fKwYQ0BRD3kjE
7XtKoOAg22nv5zZQT6Gku+xX4kTUv42y02StASvjhAJHvgw5nGYIYq2KvPmBkKeWhJv/YodAhx+m
XFGOV3ZlNPyiBQ+iExT7VzjuGa8zkcw/19ZbpH/0YcrmCj8/DNjhrHo2rnjLFzD6Q7UnZYyGc2Er
gs4lOFbvXuJOvFz4bqeEExDpUPUAaJymtlRwUnS7oGiS9kKAq5PsFAkJxu2m52nchhxO9H3p3TnM
spazgiQDcikhpG/91B8TamDXfLk8MfUjVN0pHYXlOTk4eTcDDXW2+jxHtKXst3uXTBJE1/EWSoRw
43CqWI3cASts3dAoPkr+WnSkEV21/0qlUjwRcnLs9V04AbGrfMrVEJZFDln8/XVWujR6OHWcCZMj
vfoKSrVzjFcPPRCdNxqtbWA3yA/Rh6UgR6txmP+IwggYLOQeQZO7eFqorr+QDWd9AjM4RYvPILOi
cAVC+fr7u4QX/LCQk/9igLAQBXS/QlP8kN2H+m+RShXKAIohiVsWlrq5of5fcVDnJ74x5mFZ2ZKe
butkGZEsqZ6idfF1CClzBueZ6fRo0UjI3NqKIimP193DroRBmADTUrjFtGy1bN4uTPoXByaZsc0g
kHfy1A0XYrBDa1j8qGt01XBa7hnnH6/zknaZdrpqXKBZL/R6tyHw93aaS3RKB27vfr2XK2TAEfXA
ri5jx+XruayBAOiS5D5wTbc58OFQPH+tMAkQfBBORnfTlmDXD2VeN/nRSgtXFXWA7L1HKhTjN5+Y
79UAUBjLZE9DB7R8Z5dmolYVUM2BZcLEDwHH6bHTR/rkH0Ll6/vTJo4Yqzt8GVzSuHtbFVqFpky4
2NNM2+50eMpflLCRDIqsBvuoUISq2PT3avtLg0KnsuYhlK0VRU07RXXyYJxG8xo7V9kV50prBDDW
/klo26G8gYVFgTGZ5ad3rqvybmEJGGQdRxd0gEMFQetq3qhs2ionnwDHKh9PwRumc1yzUHiICV9O
rUp1fyA+5StpRVQbcgkm5v029Z9xiC+eOMHXtyWU0QUXncZ7KhW670BkLOHWWN2bcuamm2MSoJoC
ypdwdvi47m1qB+ub/BkATNL37xSr76eCayIxoAyQXks/5dcvJu2ImsWb3MLgqm2VEyxPN+Lzk78v
JF2hzTwpTV64tj0z7RgJk5CuZMueH5gQBxwqKeBctcNyDng4cgIgWelFq/+pSNd9UgEXB/przn66
pOyK56bCnd8209SOXFw7npNnNtKT8qZohbbHH5uez63+uA/MqRahsugkMbRg/bIf9LX4oHnxFyUS
gRtiFSP/WUAWRG0BSB09xVJVkuTxAo9Zot0Pu0v4bSk+D2d6F88ofbm+1VxlU/7edURaw+Ewll03
XvEwTnez4j+KWkLQsSpSD7Fskx8yPsBXD0wwbKmBqaCjEBMIaWJ8PBPuLALLd2gpdqCB+Vee0VYu
aGOj1Hc30bIEQBcqp0khI9so9mzL+ckxOei5s0hwH1R4PTSBBhB1ox8M1N9MIKVCczeFXsgoVkxj
Qm/L3mk8OUeRmiSEtoC/MjH4CITGW1W8OVBOJfwcEJie7ttAUUopJSvqSzNnYVDkatoLvRp4GEWy
WNQWZbneTptKZrzgip14t7fIDeYnYVCw9r14htb1oCXVAImgoi6SNTIk+fKjF32/j7gxbzb4UUNt
f6YqLjroAwD/AE7AOIRNpNMns7QgK8CUWu/bUWeFuFGyvU7jpNx2C7sY77oCm+WQxrQSQHwL5gRM
vF/mn72alE7wAQDk8WBws45accZKTIWjd7HDQfOB2CUTzGmH5zESK6QwW/vsAwN/b2ioUqm4CQoD
GgP3TcYzjrfiOJ9IU+/t/lpe+l0oUtdZ0XRac2uJyC8sPghRorJf+Pd3AhdotsmfHsBv67TgkqC1
txUbDHNzKBUePpZccmxCv8zbkOxB+OVH7KiyWjhKzNa4xCw1PjYZC+VQMj2Mz47SnM4kfSMxIAmG
rFXOqLMf7ohqc56vmQz9fDi5/ydH1gFLAapjHb7CB+t4TJfLYS/503DHcKj9isV3u8YJH659X4ub
iNJBwKxJRSjmMtWgjeFy1tw++RGkf2fbeYfH1b7cqvGd1gK62EZK9bmys27ZWSXltvdSwmaTvF+3
yKUenkW+6rkNU+3CIcgz3+cPPTCisZ/fWdBu+Df8lRstd/OgXuuSAmD+p8iGytWESB6nq2idrEwo
vA1vLEhEzKRdxvfqwZYW3MSthe6hh2GipZv+uk0yCaXssVfS2SccdrsHfAnJvs1i1xHMzoKDvMrT
4k1FSevx50vwvtOOb5Xayo7L30vOkautwjI25oBbm7dyxXgntWBe/go8E7dCX3dhHef6yhwxjmti
zGAb8kW3cgQcvTRKaXiSQ7wbLe3aWCIo6lJNpVPa8hfwTvcIGND00yT63ZzuhDIzZdaIN63dAO88
5hKa9upAZ5sSpBBlz8rZB8sItVqHXSyaKQVBqT7FpargdMV7E1nnQWGWyJHjEx22xSXRFXLjPE7+
GPC7Fe8CHlifo4xyB+taZvqZBh0SOP6sCpfzQPQ1eE6r52jQV+Bvon6b4//MXgcnbKh8yKeUZ/KU
Jx9dTN8FGTBFULfnWwst9SoeuCeYr0/1fIhB0MUlsOj1tjH9omKRamvwPZy0rMCQw6K+uVWhCpe0
bG9v0aleIWsAPXTjFL7rYpCjWhytajG0F1n/TCKV6I6Tt1ffLy+YTk7OuM0fVRPe/jtG6ee/vPj5
ip8aYWkOWOBH4nSQ52TkPikmoVImkhAPTyZHmkHapSTt+5qqzw3wuMTeK6kTEJ+/wr5xVKX9MhrT
B0PMUEV3XVsvmZ5CirQ+FWRsw9aV3pB0wosErkfyeuK4dfDozjjn1qqyBfv4MHySIdA2S6XNJEnE
3WeNr3vu+Cdg7xE/9X93bzFGX12+WlTZOqFBWu4GjzgFAtK8mcR4OnbP2jtKGhv84qlIS5ppCkC9
mTpIIYuaYFAUQh/Z6eBwWtodmTpgUxDpe3FzEt99yRaBlOMy6sIBQaOusT/9yRj4n0DGUoSTtzOV
aN7rryobAtV1YunrPkHe8nYCZ65rFg+7XE0Mws1i1HNulfmWm4ph0cetgIFVEn5hxAfgtTtkbjgI
2HmMs/bkMtwkXwPbin+iskG7haMjQbAMo3FUJNstVNLNFy+UkeJVjcs0NoSQOaaYK34LYIF7Gmup
p2GA5ELzQ7DK9h87LOg4WkryOBfDsqQjkMwMHdNcd0poWtagBSOf9TN6hL49KGpHs3al1KYlIe8k
7d/+Sn9k/HurJydQ8nBAtUPnbmgxa8om07G+RmUzdynBbowd0MHXR5YqIcnKa6bdPGa/om1plRvf
83Xkq5mCLyK9oKZDJHjupWOZOZpW5hLGd+DCQq/GPJ+HiggG/IT9o/7Bhn2jgQzAfkTCi7jKWJ5o
eGr9pnRHEqRLocbwwX2YTN6gWDtx1LAgmUIEK7FtAD+/Vb1uv9EMxPSFhWDWb3BKknjkl+/bNsZF
iW1orLlX0usAywNQP7wd6Vgzpq7P9O8dM382aF9d6ytnjmblvG+zgGZN0Fu7KXbzyvJhpjCMKS+r
3+wsZ1s4tN5eYAtY10nsFEdwpQV1c2mn09ILdw/Yc1wHJOahJ1mkSPPtLLDN1HRC1a+pAYZwqIAU
2JD7aRw0YwOQn2aXPc+8zJufNqGMgPfvnqjm+lFdzZJK/GRUB0cAiWx6k3OOsG9kx33d/ti8sP9N
W2XKXGVQ5S+OOGR2+nmkdLKE3TkdqB9CkhLnEyw5q9t3JuQD+Sw2bUxVxXi5uMyhwK16ySwbJG0V
qK9/Z/fZqE4rLM1hh2uGcB3elXku9zFOd1CzhSRX5bHgmGCiaq/b4yjQ3J6+HCm/C5r9MGuVojUo
vDIDXBw3KZLD6s5PnDgJtL+wltiNGUHD9eqwZuKce3nQ2DyDJwaScDfAD5uAyBR/VTwPQueTEgdu
czdodPr6C6X69BsLsQzkYcV+bQtGCVEdT/J4x8jOEGXlbxpp+D4/GddHXXSeuLeZGANa2eW9iUnb
x1cRlrFikg1khMqCe5J+YCvZmfCtPdP9wP8scl7uCwlN6oPvDY1nBuW8kSLv1QMX1vrGdvO0+54C
tl7PrAZ119lhdt/LT2twvp0biYdmFKqDvdsFABBsn4jw5mc6gUjAyj64eTIwdEI0L6wwkPtwajIN
qk1IN7+LoU1FrAcof8/WWbcIIMXN7DuVYXCP1VX0xcH9YjDvFQO6vCnRq6+k0emYbcpxCqZtL9QX
9xB2p3ixNOTPk8BkxPtbLWKmXsjf5nj6AUrDvM1bR/P3y0Q/9DRdeH68+qiZTn+VP6vya6H6O2g+
oNjG2ZMCE9drprBjaYlZC3mvAoeb6UVqIrsfOXdTV9wt20dTrQlBgHDbCe5vhhLISzYVEBIkwJHA
/hXtZjRJFwoTl1lvzGHY5zsSv9/3FFM6oMoip1i8maTSI+1TpIkrNcTN7EB1+poU2N38UC/rdtgk
e4D0Pb1g0wOLYbKiO63O0xcW1u7ukgAATuynht7vLUv/6rvWn8eurDXJWY5McSeexslJ4osEikuX
ZgJrod2GBBGPBaoeNBdnHU1SBXXHnslo+yzNXN7Bn5DyAcbKYBKPA6J15M9uikpMmilYN/iM9FV0
D3vaeo/ORi3pQRJcY6CFZRldzd3udwME7MPW05crEyIa9joBF1iIOzxCkVVnog1WeV7tBmIO/YK5
F/4r66p2aYsXw+1fX1gZDQJb1cqlgG8GdO2qXHTpFedczU0e3nd2NRTvWj+kOdKup5Vp9fNFXVav
EzbsT9pGlMnwMBG4lNq2Ptcs2n7teUOxAYTrHrHAqKUSQzMXsyw54v0VyhYCP+ZXGNaVmaDRYwaM
coaH3z02TdnFzwNoyBOyFRnQMiJJwvpjnqEVN+Lku1fnI1ejFHy8EOGaQ7LQf8i4A44H1hyoXkY8
8/SksG0mmJRaA1K+n+M6eAtLaJvleZ5wHDa1LgJnI+ltd1vR4gqZx/0W6/rjApeNYFaIVYWJlX5T
j+nJC+6AU9V8s+O3d3EmL/XE1fm/LJfuGMmgplOb66hzwQjj/2LlUUNchMojHD6U8BTwOeeOyGB9
or60efe0SWtXVqpf3ZJxcVNy+ql9U/YY8NgjKOAYqZFldsFotaiFZo7UZd1O3DkKNfenh6mRqWOg
vmJADkqXhxzrWW0iF7DkCfBaZuy7PTYzvYDsnh6DvPKpRjOsxaHwSdULLL8s/098tbFgnQLdJ/aL
lfoJlfaQSGqTldDfwdO2ADTlfmrzHWdsUqJE2YNUQV6r9eU/dt7PnaTAdC6zGkPiFVExmlzsuRT0
MQIto3XMRYMeGD0nVQQqo5QQyQSxV03ZKwU7sAppA0X/+LB4XjlJjouLNK00ySDi55I9P++DU3v2
bma3OaVhzqsL3UXY7E/1KOnHfNPWhWs/mfKLrwD5hgycGTTE0eAgs0m9vE9emEX2Isd90jxgmlRC
yALSFUO9ArFxaG/4FPY0dhsEX6EG4tacEnRCTTv8eIfg9+pUgaFoVQpRg26OvKRChi7UQ+pSb6Mk
frW1nvkkv0nZKMlJ+oQQ6LYSvRMXXckwdXiuBNEcgcAl3mt2nU81wlzDKpWeKSGE096DibtnoEUV
UFJ+k3wfzVWxhflhSfjPlwmRKvL3VfDnGDVsoTqiwbKVXfLwgHSFiny5WOsHAjvjQvftVkO0iu6y
wkCJsCklJQT0XN59rXRvygh4U6W1nrcZme2Q7UcHccF00iN3oSG4KkDINObntghVE1P+xHaP/JHH
KXefUfEQwjsprGphVzqsUdJ6K/wao1X0FDSU/qtvKYQshvakrLqVde2ic251a/mcX7ojnqzYmBba
momm8HiUYGCaQ8ek4rvoAlu9QKUDUq19iXt5MtxTDRyoAKFvw7on0fC5RVtZsrWJ00gQ0z0+ukGI
ZvE/ZS8M7OqVe6r4oNDMq+6UloeuX4k5zaJXDZUmKlMwAEZkWJPs0uk5OlIe1oVPOCYpwx9IuGwf
inztWSy4MJREpb8fwgA8yJ0vCGJAURof3Cc8N8Y2hXxj4xajilIyi/R5zCMw24nEPFA0aWq7hTyu
zwBck57OqTAQQRRvtZR2kujXWDjCELoWMao74ERBuCuUmcn7jQ08ZCthKb4AV797ObxNuBt0Px6W
OlYkDjGdw4YVJBaXq4O6fiyO9przUcYW1pRJg/4pnME6wQP9IUEvst1J6i/nluxpHrxqFF4CXiAo
pna011QDJo6x/GKTS/qtwOgg8J6YJUtxRmNbM9F8/cZQVAw3ZDtleshXSlygyIkgYR5su3JcMK+I
auBJvxIYVM9fuLF84goZ8SufaMOLFoo2QTFf0jWpnQ672kI4Ph6vE0CVc7NJihbHWB4yz9QIpnH5
cWweeqLVztoJGBnParFrKn/O742rxdByFPwDtfOVM9XFpF2NmoxZW2UKzwOW21lL8Sg5aHCiAh8H
BU8KKMLBYbbJ8BRj9MQ72zoEOV7r8SFmIxVhOnOI4fdDuko5FOISgF+1X5SlysAZVBf4JS5d1HjT
NHX/kUflbRDNhBpkPwr96ZRjKWCiE0GjdN0MpizgmKq3xw0Utv29kchlmwCVpIU4Wm/s++KlmRlU
qNxAhs3L9umykIuauuZ7ZN/1wzwJqQZ9XOKSiN6ewtt0qw3h2YKRjwlQNcFAYd+gw16kT1MAtm4e
Yl9l685R8OWWa134qGaSt6IIQFLKnMmJH2Gy3TGPshX6rh6CKz70SsBIYF51w0fo4RsZiSr2+5zF
lnPHwlpt1vM2yitxgt3kYSwoCx+NJTC6PC1w2uTpYgZ2Mk70NOeAvjHY0ISBQEypsOZjjrMjXHSP
WMEZcPHhQZX3fOGWg+1F1LKNYhzK0EIgop2Fe/8nlSD6dc9guX0FiJkpWZuHvVEgJireiOswGr3V
cQO5RqME4pPUeCcPVk4cMZ5YNqcPfqjhGYIjeB8yO6HdmjC/fSuBB5qbDbpLYIGZCv4oRlTffqaF
2X/nzIf6DcZN5t9KIfuF43KaOt6tAoMz5b0AI/z1avqRH7tv62AjWJj/mmU4dOFmSz/QI9mNEwMv
6TWlDWI/dybicOH9rXrYO/c3X4cJGIynG1DO/a4IJ2BzsXB4veXTFh7dMfy9JfX/QLWQzx1TqZYs
NgFcYPcu4NQI7YxJ8pvmzjZ7cEBs3mbRKorZb81TQ2poGzt4e2hskL/645x6jy+pyEmAKUnqxaoZ
Ls8hlhdSLGAg7zq8S2O2U71Kzn1PcZ9QpyZPjV3SN2AulQaXJUX4ZWrom9WIIHvRJl/MGqDWLka/
wnKYpJKrW3g9sphRCM3cdexy2kR2q+KYx0TiZ/dZbmV41GtUCop6jPFhTgmoYVL/WjJOTon++gA7
sTIjq6rnDBaRMHPx8XT2KeflP/klRNDSaUXd2BUz2Py7GaFJDaIVuuLQP2IQFMXl/8ygO1HdmdGI
G7n4X+7rY5IAvdRJcM1QkVQGrno4jpobSKzL6dYCXmtBqyK0OQTxX3iqtvWURfUDk87Y+bJgVMMy
8YrFFet1Yg2DuLvozIiK3uLd+jptcZBU+VGxUEmhFHPM3qgTcHnsOqf5RrxVVr7Jk/agzdTG9BT+
T2HIU23JrvcaPAagRjj4Ze2h1mSXlGxOfZi4KNpWRVb/+/cfH+mQadnbfmEeIFn9oMgqdlwaWhwg
DBPpxGFuNnk7R+0ReJAjSSWp1XmUsydVTc06FjFMSz5lVjbP+DBiNxILm0pCKnY1vvE9QGwezflD
hwrTyuJDmhpZJdaK4taPKm22R25gnFtoc8RyGDeWz4hrY9xHhmwVK/mOg4aCR11B0fVFQG++duYT
rT+4KeVdzRMimxh0hxRaj1Qbr7bwqQsdZUPq8mfvaKSko5jqkDgj+QHqwpTs1iM8EFZXgcyRaeoS
xLto6w4caChTG3lBN4UNbY8eFPW/LMtS/p/3Ze9sL3MFLmVZ7K/qXfyfYgrdi3dcj1CKrO4YObCp
acbhluhy1ANrsonnRQSQBk7Rm2sF9tplh6BFcwQDhn1WHWWtWrqjfiZEWwC5yXA8/LX6kq2gW5Nc
ZfjvuGRkWrNU4mnZfc46T53+8Lwe9QJhleJg61oBkC7ybUoMjrtoLDrKhRAAjR0DS9rggh6ZcxA8
n3mNzYmx90PlaTqzRJPXbhH3AZK7vN+zNs33xP3MXv5ue+mBNiXKAN7oSlvt5ZcPycGsyV/nDKn7
v86PhWh3ITWnEIHJh0kQ2AQZMZUkOShH/PE5xcYQJhPsheFspck5V0Oh/6jsY/ouPP++8i04Q+BX
wl9Do3O/sSDzVlCik5vJDozSm2eX2Bn4yBLZMXHWx3TFLT8yE6Prqef9SB56FbSEVlApFs+3KabE
SsvAm4QKlqTFRvM0BnlKxz58NrKJ1cppWrXrJronCl/p/K6sfSDeLei1pk1qn/TsWQRNJAwwYW8i
qJuEXPsqnxlRdNtLQlOYH2T4rFmE8E55zYB+CEBQIMpRIEql4f5GbFHA5vRePhcxYtMozbVcP4CC
p5zrw9fLANpK8thn58KmiD2Q0snxxHNVx6swj6I/phaPwu5D+d9SA0Hhoqk6fvL6Kws4/JzSFIeb
sEtstDjbSkaWyWERYPG39Aqajv4Tg1oZCligangytO/yYM7ztIdBIB8PUjB2TCUhjUcI9GVL2p+a
1jvHUSAZnpKvDQbOv3eqtulZdvxgTQ3l83pZVxHiyY+jXY1yFZranal3ZSOyWmqVkA4NzVLVZXME
kEWojTOzDlhquGuxcRQ/+0r8zXfgQWAz3o4uEV7D8LVmsvX5pQNhXPc8tN/5q3RedBHzUj8R6zBP
Iz6AO4JaVkHhErJcmA/LAic3ML6/gnDvccaGfpvwJRPxHUxMpcNUwKHD7/1/HmnLSj1Lnysqiwxj
MoVu2n6lLBzHHU7L+SxdE7kqI77oMQoQVGhwSMUKYXO65hpTr1bTOniI8X2tOfUSVGrnD7IPaoGz
t5ppmjIimtWumRkQhI9SqbE1shWrSwW057AOTNIUNjryqvmrqraKQWam8apK0xXt50yBbIpUeqRA
SK0jSHs3la1veLG2WHEJNn+i7jBDFGyHehY2idx/L0STXa+bMbo9bp0mhsza0P8fnn/lY1r0M+jB
yujbdj5OaAJXqa4tQelv5c78vM4CDybHaQ/N7M1VWwQi80AXT4C8EBEQASAGcdO3xfnLR2ABgDZj
jVaOUstFHWl5gSLOerXSVOge61QfKUtfpalHGu9GKZ3/v1rGYI9HCwLM0A53g0rbamJ1waQ6G3VV
7b8wNNb9Nv/nxMMsAiiT7q24USgGIobvqxhj2LBnUcmBHdQsyYTVRjEOI+l4A+MBJRjT9Ppi/9mD
q+oXgP85lZ4uzH21vzHp8DnBOr5Cyc4mjFIfhQaJF5Dwaf3JThVY2JokCO6D81XrF2ACZdMf/CFi
CFHI0GT6YeNoUqpzEenjdCC2p7dJ9JDvHmykAHuWVzpshDTjot8kLT3c1oeaPNqbZLvJessWWr3c
gJ5K6/ydQSHKMQYkPNpvUwZMnvdxa1l7nbVCDSCoXihCGwe8G0EV9u16h3d7ZX+N2nkeOjPKQY3k
B5AM3fVSHuO0wAmraue3c+IMtJmoXuZkaLIJaQz0zyKku3W8gDnnc7Ny6+nyKHJ6+YOHFi9niAeT
NqKRwZf3F0HlsK6V48UGuuuU8qqh4uq77OBlbrhdcndMrqXu0LxCnuEZb98bj0/vTPW1U/p+mooa
dOkBFJKmDAOmx5u9MxcKCHqqRHuVHpDo15eb/AFxYCQYRckW6t++n1MunGmTSnFl0ap0omcMuuDX
X2tstOzspJJtU5kc/4RfloAXxltIgy1C7Yas+cxn5X4/nqkSJeDaqNtkwr6a3TwZ36lfQF5uY0g/
19Eh0K6GfKZOE53ZzykrDhS5ndIbwXEy7PI2Pk+BepPUpracV5AUHgYhSoAPDqBAdpiR8yRsEbMs
lpkplfxkt9YykNqIRy5VsM3q61nhXaQX7twnKDhbcUdS90SOlhevk9w6Jn6NueO97QJSELj33j4y
7/SHOa0C22vodBb4D3MAyK8zEh4Jytzpf6i8RIQOKoR8hRzKClT6EyB9RPlz1Hwqe/gjOcxGg6qF
fyHPVmf5MW37n4wEt15vcJQYwLILEaOMHKjwb2JcZgxWi2+LE6wnrYEX1zqVwaLOKs7MvzzfRD5r
kuUHS6DKpUGJY0wRRhnS0LdlxnX4hpC3bn4V2nWzktaq4V48DW4TwK4rpHY1SRr1y5dq903Fen5r
pea5qaG0hHuf9mioG6TIhAuC+bLZUHx2Z4CCbN68q15//fVLWecNWOFIFNpFpV2IAS6Pg3/+3PSg
43QNEOW4w7TCKGIqZW92MlmkIqHajiQdOb3B8yoMUXcrjcxujYZzfSEnMQZSp/erKl6N3Tg08CZA
HNB9X5dqJPd0/7+5aN2nmEiO3lv5i91ziEmIWE4vl4TjtNkjafITewrkhXtgc2nyf1M8jGLgiWpY
k6+CL8ameNBRSx0RxchPzsCaEJYayi1U59zdhW74L3jclaC48ActC+SExZGiZEQNXHeCkDBprU0J
SeIsn9Tha2iWsuPgBj5+4fiNypiCiCsV+htYCiNqte1R/yT9xdfAYhn/JWclGKInjSaDcmjdu8+C
X0eJS1jYml8kzj9oXA/kU01YVtgAipmj0nV/lr+uZQ3evxdc7UZiC2nDq6H38hstfIx92H8/VeNe
jlr8KP1E2N296DUNlzRbBp9WgRk8DHVBcvPVOxf/285vQ5PeOO5CKlxwqW7vMq2oW0Auv2S/FQZl
4lVEznc+d9fLNQCSLoj0OcWqktLBcuNl+eHc/pa/mP+MdFm7bkECEoNiZRQscOzn3p9xfBUxKEtJ
mWM1/8gN+diiaLx3L2QlS+35vDsUw88rmF9T7uy60Xuk4f0CzFMPDqIlDQqMnPVAdn4HMB2uJ+Qe
sF2PbiU5NLMilt9JglKDJm3kYX4wb6fXNVWIejs4vPD/uOJSqhFTOoT0Mze0/WdNsJAI72f+XcVG
JZ79Yd58vcvccKd9stqWRYgsNMHcof8hC8c1UOm44q/cWcDFw/uzYRBG6VrQoOvHEfgr/Y8Wngg+
s4ROdQzqZYzV1s6XVSh7gJoT3cDCK/bIR+8zdinW38pwRPi5pZQE9g1fO9/p/2yqctUZ/wKpiCy2
Kj9gic6bn7pjPDIhS0VAufX//8mNzuQ4XRmgpr/A6t1UmoKhNvoR1AlVXKF/ww4dQd5XHPBu0ZGI
PqltQH80FqXQa67+Qj+s/NukSrrSX6Jlh90bYHAwSSNAWP899Om/XRHUyxxAbE9Nq6/QdPO4lxWh
x4AEaKXQkNICDDgMecqi2NXeMWrbl3mdL68/4XxoZK/4NWRrwvVx+XyFASwy8vb4j4XZv3vLIYr4
TL53FNSMRfRyB/WfSkpE9i/Ie5nCdEVXXvJzlD+Xzt/l2r7RyOI7jiD32+jOHlryAwtcQIw4AU64
vFV6nIOiCVaurAUF5pA3pb0GFRhqolewuqP4wX+oMibBx9N31DH2nRIOkRUufWWsgcMR3IWnF5za
pmKeKNfbfqSFzrDJg0M2J15tmGLGhMw9hgp7elhx3ThWXmr/oUCURZSvfDp3lf7w41T+gad+b8qU
b7bRphynDVvKps5EXbwbYiePKJ2tRI6iNcZ7gl5OKWRimGqilqImx6RTFppkqsoR5qEuryya3bir
leyFEnqwgYim8XgAJ6y/B3/q3sTbR5dwYr/gX6cF9+pu8XWc8qAWlBJ4oEbm4q/iPDOwDJf4BqR3
P1M9vXa2mODCl2V260Wp0QfrwqJyOC3zsY9OGaM5SV13ArRNkRXMotiYrkR1o2KUaxl3GEqNgKbD
WFgoAlHybf7SYsm1r95kwgKpm0HJBjAeJEbnDtl9/o9sDFAIdaLlb0m9799aqONhFm6CEnnpmVDE
qPc83NmbIsOwUCH6ln+woPnZJjq+K2DBnSFV9fwcxZ5NsoNa8L8PbecFEdH5URTlnnp+sJL5HuV0
BLceUhLhEAYYhxWlHcKkmOJ3JLxMsgX6V2MnnOPn0cCbIeI7/oBMPoRVvvVxDtj9ZmPBXCEmRtyU
dLE31fMSfBoZglm6BxL0uMzzRuB440fDUOsbkoIxxRbWh8XJGlQl4xveCvXy136fDkTfwQ8i4RaE
QkgGYG3FWjVgUQ/QfrsatRTqD0VZsHXqQVYV1b1drU4bT338a5nPTRsK2rBJL5u6IFR/v5ByEnCF
rvIZtJDWj5vnhHySVlEelmEoPQwTZjnyswTFMZls4d0+EQTJIjnXg151AYzaoYv0cHGgkCu6ehfl
2U5T/kUzhwdxsVRxRhyibRnnLBCQlF7YP8MYWHjN2FMvhV8GcJUx4ZZEBq2+movJsId1tgmv86ew
84vQtIPJAOCTrIoaScZwY2OWFJAfS4+AB/Bxk7EhP2m59gGxsXMoIZepcNqfjnVj7l2ZVj9aHIJV
O3DBh8dN1Z3sYXsCANIR+bNyu54FzLAJozDdQVv9YKWjN/RS+r6QXAkEQ78+MN62CG9DsrBXxx26
3S9ZWNK+b+f3gWKmEUTS9C4UxrjCGCbFTy4uOAiWo3/3VAEudHQ8O95QHay886jDuxzdUimMK35f
H1UZ8x7lLVyFi8DJ6BimZ1zyZLjoudxSipve0WWNQzGV5uNXJhTo7y8hCIL/78JBdgFpHs2P2K0E
LqDLJmiebK7hhqG0s9tGUXHVx6QjN1STXO/GssuX985KuOZVkhnhnVB+9h9mpVhRQN4TZ6HkVKlu
UFJ5kFjYMyDH2rpfmbJd/nDQm4mJ1uygIBZF0ITRaYxx2hhjgU3KPr+stn0teZDlMrB544xLJOmy
j3/1RF1ehGgqit4RpTf+ZkMXkTi4ogOrrUJwNqt9aU5KQknagpXy98eYkxSCruz3ZgNIBgmnjM4P
MUwfaEkhZyaTfgwX3wMZ1svp5eDsA0SgaPwTO4msb8SyT5PvVA84IXiDfcjA/it4S5Azg7+1DEJy
6lNMj4tH1VM6TucW5eZdSzn585+dQ7E8M4ac10ogtpqrs8lLF57kmF5mIE8k37hE2YObNWLvVZay
gxed+PpDDLIawen70sjGP3SUvnVlbbYpOP+D5hQnp5Z0rbHDNYDT+lWNRWkOQ3i2vrpf3RbBf1Ay
L0rIE7T4o8h9EnrDoDq1mvx9TFNP76k2I3HptiunAoj8tV86pgvH0fEyeRbv+K9vwvBITsfZisKx
GZCTywCkur5mQqWurdl20bV15Kwa9jh6kEy/8gkVYGfhVvOs2hGyahAO25oknV0DefkWbradJkAv
rZWWK6PDY6ltxjvzqTaQe8lqDXInWhNZk+D54YPpHLVfJ8MFnTr0Dy8j6igV4Ev2HyIDtcIG7Ava
60mbl5dDi5nIO7rXNItKn9B2CzY2D/tO31fvNpdkMsog1Ozj41DW0BJ5AqIEVmbGcucAYLtg6xMb
l9lwhtfyCI6IaedltLQ9AC4qdnOUPk6ZR1HdWuKdlbC0REePKMKwmI9Hjg6qMpLmstxUgCGaQI0U
z9zPG+ZpUcqLpU0RjfKmBjCN+KHB1PWh2MoVu6UdNvXnnkEk6SnSh9NhieG1t1unbUtUn/8lI9tH
jwI6E/WYeKUU9NlGTDY7aQPRBAxv4OdNxCht9RjsO1YSCH55wKcr8No+hQlwFk52yCLiAY/L+WAz
xAxmEDLKalBHJ4ybSgEqSZj0PznMxlBbpff+dJMrSF5S/PAe+x77E/1e3gSjtCiOPoxEA7quXHuX
VYgm8H3RI1Cs5dTdtG4wDV5O9msiAXMnVYlhJ34NwIXepyc7dowsq8yy89JSddAPXDHD570qGeAp
MVRWmnNGH6as+617IRn3dS7UnOah84cO/FG6yGFAGHJx77q9m/0t33EzfCeR1rqC5zkg0Jq+4TBS
tvIMtd8zRELbejd3HAyGfjpr1/s6PHKaiDzR5ZKCHgGB4LsR1ZYWqR0PCB5j/Q8vRyKFUJtE1EqK
kv+nak9DAedCmZTFrO8uCEGP98ad+CO6TgDDDUpGCuvznlyKCXaZ72nco/EOe8UL/zrJgurY2dgR
IXdAqDkaQY6zcQKaOKiDZj1BkE961WOAJASiWjM+bsUU5nyyZ5KN3DX08JsG7YEfdaRt2XfjiO0x
TSXi43AtqfOrYHhKkuMROEavGbBfwMjhBnvMW4KdF4kvYuOsoq8wg/3OvvzntIIlpIT42Nouy3Je
usCET48xsdG5HTUej0XZ/BBQGThgYlq6ZbSMej+kgKzejkUl3gTiHJ03vFwsvoZk7JY4rgS5Ayrx
enC34HfusYujo08MnEkkSJK+HbuxTctaaqZ6LJZaI/ut0ASapevsp4427D0d1OuJh5N9LmbThzKq
g89lgtu9FQUNvt6fjJ13YJtBHkcUC1OuPwML4zDDrlxYWZke/OFFMoc9dAi36tz4W5hVnGMtOugW
PZUZNz6Es9WE2cF4DY2fa77Z4JSgkvZiZymN70aGoF83vR6DdLBSNDy7LfQhFXkIoqCl80Pqqx/K
00IyVL1sDYCX3EJUGF6b0TTHuugICMrB5NOeqbZNz/IzBUc1x5LHKqk1plSJpMjtOzP0vz1qJ5Rp
A59Rl+ENR3lbe9VY1ot0dzsuK81LuZ9tB4to02HD38KXtBF/hHK8YuJRP5zyH3B3ag+mt/XbkxkL
qGaUnaVhcHExHk7qconkwk5F6dRbgxtg9dsxCmlsIRBVcxh+crzDIeHEO6HorBZZaCo9LZCfoUnb
XG90SceAMVLlKseptC8Fdo+4+EJH6a46UCNxRyIw9YJJ1zDrCId2mwAyWyv6aKdGYA4ITrduNOxu
gK835gWS6FSnEQ99Bvzst/m61nTWRDGSEv1GNMgNE1hxbqQkwjUXEIPe+6oS91zNcpyqxdoxu1hD
pJTKT6DG3QinLtqNDcGwL86jZSoWLVCGjYYk1riaDTWBU+L/wBYnQiuMh6l0KGNUk/jWKR6Cd0DI
cSeqbRlzYLPeBFS0ygAE82sWTjZtlT3ur9wbir0lnA4RVmKuqlEJHqbcmIp6TtRLOs3B/mmjTWZ+
JTKgvD+HegSe8EeXFd5Af1ndrMK/H5E6PCdP0uS5Qi18kJreXMwGXtcJlAt3VFudCRARWNnJYArW
N0aNCi1PisH1AvsJW+ZCGu4SvF1rz5YEdavBxVwxCCnXH+hXCwTJQROwNuvATWOqAAVrMFwC+fU3
nFoj/aPn29sO+DbgzkQ9MNjIwdxufhwHVObMCX0r66tpml63UlDVil3nKMka+m2BANI5n/BDY4Pv
OTgmPabAZEqdzbxXiSRBq1c/Ks4LEFkzBVCEhih0DRTW0zOJbLhhpciSh/NHXpjUcMUP/OPj6dcS
tJAi93r2ZUhCLRUMfLnjH0bPt2nY1vmuJsqvmTFX/gT32/Uq1sKH6MUKpBPINlSfyHshHyKktBYo
dIdkT0b4X9qIUbZTjY9SGNc+ijtS21JwcFVnlkLQaGn6/sxySLQngFt+jy8lKG1F5rHOmp9xjTl4
9fGrnoUyB81kRHav0ihHq31vlDEsZZCC1PONrLYUHOn6gwQsaZQv7xE+AYzfa2F+96l/L/roB/Ls
hQgOfhG+8Yha6xiMz5Z1ylYXx8U+00SbtwY2KPAEJhevyC/t2RKBOHsavKJofVc/YJplwBe41L/V
wOlcU77lgt2yG1Uq1bBZRbIbacC0gS0V58oSSmwqb+SlsuMwmozGRzH5v5oXWKOYdwVZ2/ASnuKg
ignFflXkNtykquCcCS0CH4IDT+6xz095iVpnNKF686jop1A6Z9iM8m5HJy01NjkDgk9KZ5ZowjMj
DhFb7LXyJzIc13Uz+zNFJ8rQWVg1oXluUXv7Guh6oF0fi5KLM86kCOQwUXag6S1uMRX4mMWTTCF5
6+Bq+ZRZmpt4W1MNm8tn8Rdq1inL+MLq/n07gzNfp2snM4/1rJ5SqVGZT0iqtuBx2dpKPSU6W1qQ
CWE+g8Zz7DDHjDZIp2rhrBfNZh7cUz1flPV0E1z4lp54bB3VAvC4OntS/hF0mK3cmtXet7ge7d//
sDd4ch7xFEHtgn5x+Iz/4KuIYUzVxSm0Q11bnaXiY5y/BchhyD7MC1U/95556Z3DbV0Ku9UQQtVV
u0lAj6ZuPLO7ayvRvPRgme+teddj4SvVz7pIAtNuF35z265Nfg3CwQFb7mBC5aORU8JAXqDjhyss
eqfygn28o+xAFg/62NVlmHm3wA9kQXNaaSQbHwIMYpTnlVviSyxusoW/UuxxdeoNcJlcW30sCllg
DhWL4Y1mtFV9juLoYcuHLPRkATXj5ASwPMhJc6IKRQ4hDY8E34XfaOLD9+V6h04Pkco17Sh2KjL3
llO+Brc6l5qo6oh0+e6rNQq+XXs7h2b+pK720fqYbBRIVfC6jTZuhE0Cwxx/gXpfd3AcKb6P2yq4
9GiDEjhYLhQibWo5VaLo25N160RvtMG7XRu+438sSGne4IFiIRaUkkXN7y+nLPY+j0oZKYJ/7KJi
hKoxWfmnwQvFSXJFLUBRe/wT4e6npRvizr5NlhkPWOVHRgnzG/gtLXh4fPavgyeC7nID0H3CFYYb
WvFrtESW7eytHYVgH00K/J0RxhuQ1cQUGl13bVeYjugfDFnf64iNVfv1g3sXLrBhdFGx6/hwsqha
3lkdkFQKTGhMRSXtnMhLQTWxZZ0Ok1ZEneusqP6+rMKo34A7DcLbVA5haZ37iA/fTtWjaPGJgzXf
OGGXgdQtjACLabYnSlHURC2yrFYnED5EP47yqOC7Pu1OKo7YL3LAxgj2W5iyTyMhYA52/3XWnHa2
ls+oQU4pl3IuMn9Mb7jEh8XH1jPBYLBMhd3bUPQE+acQHL8qrFcaoABk4dVPH5hFLrWaqi1HhUSj
68EUm7drEDQKxWLHJOwLvI7FLvEjAu0mkGJCkJOa/Ch2zQ2iRptU6m19da1ulV67AG+lqvDxkum/
4If/dm8P+QNQEkSOJNZPdpqlO4oZQvpA3QXSPOLvFS3XKBxPRbLdVAUzVRtRQSZHyTeGyo4W6UIS
ThhJghaA2fc+ywDMREk7gmIF5B4+Dy/vECkDpK7IIEoTIqpL0LuDH0kGDlLqF3v357/5GFmUQ2I6
7CTtDfPu1t/AmzAlw2x3Mly/UmjR/y1jvuBPy/UaHKlS+qK0mrX4X/hsVioemC3INT34hSizZ9pl
L9vChSawl4H26bgehhhROWhLzNVPK/rt85WsljgTqtEKmnibahBkp6JxUgHvokpt7twKDqfRP+s8
7+JPd4cv4Mfgb6bP07QKjf3Enz3VpLFz71wltzicxfL5rRJNVcRHtiosoUCKe8ZVtc3bxw7v+GCE
twbvH9B25AgYnwqiEPb+nFIr39QIz/SfRnspB/LgzaLZrwTRXFrAUhV9JdM53L7O/FwtJf0pjZ3Q
EsX9dpemEj5uzvbEUK2WIitjuinu5D1s7lhr6Y5EaEQ0j45xIngIBgYYmlWONnu94Gng8nJ8eRO0
eGNnp7RTe4Y3ffWZvfkwLVRcANMviQVxA4Xl1wY5ECKocyD4kYV47ZzR8gkp89PQxBjOe3fA45io
+Bf9JsX+KamKfSqa7gwmgfjinthbaKdP2hPu6F53hVb1zpl1Qc9Pv+ZkbGRWjIHC4Ribei/CBFE+
W4HKSh8rHHLL8oVTd1vw5c8v8alhvBCp5eUm61QRgeTix/WWdEukxwt6d5wA+bBO219m5aq0kyzM
b1YOIu2A2GlIYctzkd16AWW5ZDYJUbwPFbuubQwxpz7Xz6OTCHuHhXkdjttIqyoDQg4LViBs+aK3
Qvtiwi0F5qDfAGkHeCNvfh3R1+6QtDDYPRKJ5Q0yECu/Bt23WORV3vAYElO3QXgjO1zZ7nstm8X2
9cMYHXBUGef9UdDfwNzBbOEgv7Px7PZvP2NRfzuZsYdyQy3nUztkgulnwoUrAJXadahZRwivsGEu
eyb+XVpEqwbEMDu4MFMXow0QfGk6/YWX9iQlSTFUUXZajSNYNN4sfkRgwW30IvrA0fZvAaSNdne8
hgJnQjZ0h89ZtoBDPqbefC2pJde+LFk6swp8paJ6jmQMQKfnR4AfkLczQWPiqkvfN+H+p3BPOQCR
hiP1lOSopOp1cgl28KDlsrzY/iK8gzUGdULCYEuMu/aQMYEdH48h9UxjtYKBO7mY6VyXg9xNorLb
r+1OvJEICN1Caix+Og1BI3bYy5vwRUSaCTDdA1HrobD+uTaZRSxH44BzcJ1rC325w9Kn6PHyqmY+
hubuG1Wfr22x8+BlePcarr77GFPR93RGQymBYnC7FlGgmWK6AmTQZQgBBGBO1LWbX4B3Vmn8+ZQj
28LI971MvqI6v+hAW76Uw4GD8XnxQsfgz2qhFfUCZcR+N55cWW8YCOxLkeCs6Z6o29D6G5DWWcNj
nCJk+xRvT2KM+xLLZZ9nkuzXLxN/+LZwcIP993Q01nKccof1PV0TjFIRFta36bIcJcJTiklHREpf
XDw7g7VaiRUKBbdstUr6xSyF9crZNok7ErilTjcr8bbpuqm/1ThQTquHeiEF8ClKMuOrgRZTGuSC
Bi29ejTeT7zKUXCuRlm+Z0DuMdW1a+fu73RkKLhw2OwRS7LBjQmzHE1sn80uan+0l/OybMrsy4hm
JCZjvKD0pBqKEKFSHY9FSsjxF5EGbdKh6CRotNypvUjBOXgl1mcskxaFXmODkxpdc7AZJA2Qj/My
p4z0LTZLZb0kUMGSma57ziD9iyD74vTvxaJcEZbgFO6X5tOL5i+t8e/60qXXOVSFmDP+SXI9BjNG
RQ8XPI4484El+0Ms4rkFX1lwLku9HMEeui47l92fM/ejILkAT/9+4LdEpnvSUtcEbRVrPC+YisvC
wNAaKu6Vdg2Ud0ADuLFEPMjpfr6nUORlGLuI6nTzi14isGSO45WlY+2OodNRqSP0y4+Zt0SbYEwr
pTXwZZz5DAK/Afbq3uDGnSZSLEKLpPWuDGASprCfq6O13MdAvcIzdgn51TeHDT2eo4EYPs2x1Vvm
ZqsrxG2RDLchcIG7I44RW5oLUafZjx9TRlOpWiCLSpZtiTgoy9PF0AeB3tKCa0A8yaAEfr1h21Pu
ZuxBX+uHMwrpIh/MzTWl41yZOuoJBJJhDNnxQn3BckQd/QHWtn+IAC3q/ljwE8Zwm4ewXCa+s3FX
f05HInPDCpTCdvXRBQrVTzw4g+FDKxK7dsa5OIqz3lauPrrT9lcg+pEkKaiUMrQh96rvz7Z26BWY
81J/JFYMlxbHMzqhAQyTtdybjhERLZAmc5rDU/AjBlJDyA9qFgD7Cms5Jg6bSjy+TJ2EP4NaXGYV
eAdoyNuKpL5g5WjmUxUxNpvDk8BKz0fFijA3qIvKes5npifxVwQGC0abj3xn3N07SBOCx2HtuisH
qSN0nv1rOTNkLX5FIS/dy+CcOGBGwlyxeQDjFAOZK/p/Yqtn4FUjiowJuwwm20JnOkGmKNKjMeSo
wqjCYEJMAUMqjvCC7WMZCiY01jQwdGz933wSy6ryby1X5R18Qi2tyj8NdNfsCCkFUWslTgjJkI11
0KWX+LTmWT7Jv+A6nRBsdwZsMMLNqJsH7UFgSwFVElQX2bpOBYc79pHbU/eJzFdeJ+6lo2yk3MTH
dPtXEu7ojbuolWd0Ysibd4zZEyPOiQYkCuiS3R74+46aKKC//vN2R6Mn+0CHxMl2flSXrVhmfPpu
lxsRA6u0A9Ylx0CyvVtsPx5wN6SC6vb4w9lso1lwamj2io8FgJg+7dlbaHyoQ0tMssWb/buzyU+t
lrB5RTTiaCcaRkuuQ1VusgDPjV78T9ysgB+EcujMW+ZguSRXvlWYs2dUdYI15MpXr6XdiFy1yOs1
0m53KlydxuHRsS9kGG1jCSQSJseedUMlxKtUCcLrG0d76nI6UEnazVv1bgKMplPKd0Xf6eeVDYfV
SA5cvcU77jNUfzUZhkP1qJmPwoEs5fPc6E8W4Z+uX4KnkTVFxuyvWMAPz8z+xI/JufCobUcefp48
+iCZVv61hlDl4fp0NCQhO1TwjdpDFhWhnErH8hVJJCW+7l4usu+e2szwzFftzUIy7w2ZcvVzJwgw
urK2P/8SxNjDPkNtS6FyqNuirx21mOOQ4nKEwWpHHuWeAyxIV0FG9JIaBDcw7cduuKybVrakufgJ
0+woPQyXMhBfspdnk1BG1IYmJ6atBAyCSMfCfursjS+q2x7mm6LSjMlbxuxS5uiSMIKxJJQh/202
qGU6CzWeKUu7W/vlVpvCWJ/F5H8evATjt3YFyY56v1pqc6SOeNgTOV+t1Q+c9HPQBVanmtpI8llW
xX400P4OQJtU7sXxQ12tozJrY7MD+wQSSoa598XXeRAusBmT4P3faPQC5sXzPP1pQcKnoVX0Y5H3
0Xf0pYbYHKybKoXXP+Jf9ed36/zjvilnjWrf0TcmpqepTX4XbGuR0Gi18876SgBs2kvhKaIOJKb2
pNtWr/0qkaBmokQ2L1cPoy0yjlZRy4q74WfjzdWxxmf0H+unZl59xkPysQKDSYt9ZSSbl8Q/E3u8
xdBhbCIQZzEaM48ybSum8GUQC17tDRXiiLdm13MuPQUh4UIVj4IVb9ybTYSmB389vPrgSQ3usmTV
ZmGWMaYfEBp24+Arwdc8+bCEx6MPHM9cMPFznUe+67bM3YI6TMJBeTMRDMbuqiXSqJ6JU25Rt5Rr
IiMnrNZ/RWjhsIyAzapr7kY4k9nZp/EniYXqpwTKk05u244uW0d3BkfFqwwV3Ee5r2Hp6Jc5MYBB
xGhoRbQnxK/P9WQKre9HXJ0ZuzoWlJF+RxKKL0ipdyXDfopMe0OrppUMbk7NK5qQzX+zGCJS0kgX
AH+8ursZHCoVqfYHJfd0zM7+Zq8dv6gKUdfI1wppG09glcF1KzNJnhU5eW5STGqoaYThEQ/Y7J9t
/9fn4U0KnKZ9+0yqmN9QCr8NpdWEEKhn6bDiTa7uo4YIPVa117AiiVHkEkD+k//xDEcPtcHI/w6Q
jJX2FdBMPA5bRiChb2IRLJZzV3Lp+/LnukXlsC2pgy9ToEz1WNcNI2loMg6h9jYwr/5LKXprKX35
C9Qw3ONyowP0CpQWU9v37cjofHCFAmIodkb8ZCWpNye4mouZoq4+K0boiMMHPuktKhDzPjJak9Pi
Q6FbRJ+NCYKgowZbbhkwaeQ6hzT/J/IHWR2cZ5IzFvoIwVkdmMJ8qxhd5+ek2v94IXu/i/OBjrVv
35rivangBEBH01k+B96b0Br4md9Xw9i0AmNKXFY44DAzVd7+8vd+Co2MFu9gTU7bmb39Z4nZ+y+P
iMw3MprEYU39natH3ewGenemAIdenLJ4uJSeygEYOK27mKCdwLdJb0hbNMFtT64Lgv1UeF6vZWnQ
QjZhTJwl9cC5obEMnqGI/K7bZ02dRoWbALllvjO37KbnFciAz2KKhkHi7vPZgh66T4qQWWJd4SJJ
DnOdtndGRjNfQoDVwiwzmRjR8bfUROg3lreC6CCuxmlJvyK+zALR/ELBGCS4un2MpwoSxWWI3NbG
5YK0XIKd9qb3fiwGE3q8IJ8OJ33EL4KYkQvplWXFxMiesKYZbbLPZZroblOW4G2bQ4gugSVOedtN
9bFbkdgCCSd+kyMbmRSQuvUOPm7lCa7vXkyCbLw0RkNUmbDrCZbRouM3pQylq0sGQ2r2/4t+zIAJ
Oti9ojSUBvvyrTHssXtlluqsaijgLoU8roy0ck2Lfj6Xzi1H1v1K8sCmWSojY80Dz4ldV3go8HqA
aviR3px13HeF0ZbSiMMmP621g2/ZMtTTaAFeC3+4cMQcZf/AEovJNxf/8bUFl/apzhqe33/sNOma
1L2iPuFFL1/fpA5f5ITRIbQV9a68AosqwPlGeNDbDqmYuBIJFUDho7PSOaNmtvMb+//aoOOJBBam
2m6wvMycgGyZq2wlfbRopDGPwp6YJTSQ9cPGwwgBKb+NZvgx/LewXLy7TNAc8fDulRUgTR9rmA1J
/BQn/3bu9NiQAj6L3BveTLkUyBGG5+TpyKlnX3JQlT7OtXiaGkXMZFqTkS8arruq0Fq1WIj8q6wU
WjLWV59AxMhmChIAeP6JQQBY4XlY0l18T8f1zV+KnAa2ovQF3bFCVBj6b7e0W3R7/rCGrz/sMt+o
9gzrwd1SIS6za0gCVpi1deOvbDDIT5Y7FRqKEuuoczF980yyCM06SIk9vy5ZURSHqtfIeMwYMonG
5PYj2q32KY9ppyElEA/gKENQDCWuYMMZtch2orAgSC8KCLcUmq2t6Nabqv3ySETnHv15UT+KVDiW
I2Ptoq1XZoFNlitlJumDi1Pn9Cetmb0kTSRUMQuZEFbRLxsOsnFKvYnkkouYq0a3O32La/2ZprR0
eHgz+msfZELgjx7qjQQQX4kD5zPe826iuOgTNbJxWg9Q8tb5ZEP/rTydB6MC1jIdt0EUmK06Dwex
3Br9iIHXswGrAhFYBxKMPjNwpte2pHF7DNeUYfMnYOifztvBupSjDLPxtoWw+a31+ardXJGHTzVe
greO1AUFB08QvvU+UpKiC56jdiGVelZ4ULRb3yEiNM+rAYKxbOsLpIxxEEGhcH+veTzPuwqQThO6
57Ka+qUxD/rpkuiaSlFL1EajryJvz5jugQeKw2dxMmEOlslB74lHPpeGiOm4CjK74VD55lq9LURT
qH95Qnydre/JoRaU9s0cp4eGq8Mq3oV9ZNnbi7RizG8xLtRymOp0Ihetvyp4Fiaq0Gs5bOHBxaKZ
AQthDDgHjAFb1RVpZxn43aHcKyjQdrHT3Qy+sp4rNSg2dYE7WXEshm4K+M2e9jFnCTKiYxfVPEPL
k8JL5vgJqlVTp04jMXsE6y9jE4nAjbzpP/xX8hLVo1LW5RDetb3Vvbb3c7QKdbslhNDZr1q+I8IA
cPaHkUeUBq+mFzo5D48b054bLyJ4ybI72UAGDuBgt+WsHtZt0lM3o28os9dxeALiDdXl/347bHVx
PGxJ9WAZMQIY3OEMcmhtjdyYfg5BecYND3zws8r7A8vXv0iuupCy3/na8bKhBuKh+1Yx96qkMM/7
jwvtSxsuxWp4KwtC2zqkp6MUO6fJbEcTYTXvqwN5ViHym3Wp9mGYU3F658WqxU0lvY/2tpwJoEBN
gcqY8thkvAXsu5kTyes8kDJ7IqymaC0rdc96iHLrVwP6GmyNB4UKQMv3ky2CU9NnhkK+79Uqpc6J
B48hU1ZsIm6Sj3rRfCkoIdRZuYG+43yRG13wGtQMvYTbrl3x7ie3K1ArWUik8zeljIRY1R0iLWis
i+LvW+AP1tJaBi8DxInLieoBQve+Iezay3hiIZ2vuzQQYxbJo+uo6PfccgkjxQIBNDjilDgsauEt
Uf3K+z0CTsbh/Jm2EQ0KdLP7NlC0nTV9rxCUlpD1lskW75td6+cagjhSLdpTG/qlWuVlwYROkeMY
1mr3QdIMEjvErk44yhkVpBq/cYSmK0hpS0KQeGWO8w02YVOB+cJedog/Y9sfcltFBMgRfL3we21U
otb0M5x6HGczhqsJ0giPuSWmTwAvHA0uC2D7q2gTyPkCzN5QnR7pByBCsPli4w0sdfvAdnbBfcMv
WtBxTTbPwtr7UuLY/hmzIg9TGe0t2Zao84Xq67wgayu6OdyDOVsYME5TfZ3loxuGGvoadEEKevTD
vy0KVLPkYL94I2DLxnQ80Iub+mag8caGU7OCg3WCm+DW3tc1mor83Z+604ooC94tBm6Nr/X9V1cE
+97EJr7UdrE9eDXGC4C1drqG59jCQtgt4cDlA3OlOk5SX3jERxFBpGXVXLvmMAs7a0EAmdgpHqfW
7bWyzM2jfwyguC+RieM2aB18uZoGUo1JOQeSG2UDYCDQAEeGUm23bxUvd9gzgpekxLuex31ik+QV
ZfFRNno4nqjDGW05Ej/hm83g/JyrdE4mrPvgQkdhJPncxldkkJxOolV7C/3iJBKhGl+U+L5zHFsa
4A2VPVijPbuDbBLDkRKiCUY/yBGhGqgsvaBGgwWBHXieNnTQI+vLoI9NHhNNycDaQHKA8IueZr17
/bZ9Ux3+ZQCSCJqKRRgTIScqhuU7b7KELGaqPIXaqtTUlesTSdqb3/Bqe8v85YYtGQpLWUp7fFF+
UBrhJd7Ha1hiGcW/RBHmXXv1cJ12ZNInwYLP/wIHPtNimsvyZuliyKBqbLE6toAxIIJf4Pw7bP+h
Xu5cziZdQykprkYYCVEpCQsPaXO1FNVTqhkhZcaIcLSxOx/IVehKLW+Ej/2vXmtPioZ6h24v96VN
HymPMJ+mj7ovepLHrRGUicHA7+O9vh+tiMx9YlnK9cw0nZKPfzSItHS4+6HC3R7SAydRjfr640JU
D8qT/IAEgnW0kkaazzUBE1XkqFYyAN8ObfMV+LuQDGhL6MlbPCRb9yqCUdi4JHwrjFH988xkb43P
G518HsJO7CWHzv3f24R5+6i8qpBlTBS5iRfZgYC58BlvtxPxKWVlVWe51UC+c1DAw2U1DMue2u3T
OcOdI6Xu54qJ2kXxPpRhaLxHFn9Qurlpj8G0N1VEpdv69IQhEGLICwaXDQsVih/AuqWmBnNQ+dSU
r8cAhF52v8dMpL1d6OIzIOXnd5+Vebl5L21tSewNia9K11V51IC1sVLv6dxi9mv0Kf0aaILRuhi8
X3Rsb1IxrmYcEyQRWJ/8uLXQu57f0376XQ5mNuZeoZuZr/MEAfDQ90/gqIhm6khIdkClDsy3aWIB
cqTzrTywWvA59fNi1ODKbpO1hdSoIXG7om2DroF54Rgd3e0Pqj81OycVkS0Ku8p408kK+EZJKkAM
kM3PHh5Mhzti0oE+vA+8E4MhsPlwDPj9gl7pSd3QPDinMYQw3BiEBzZUQ4gqn6oJmMgDoQ8fapNF
a/pToy2OnXkehRSNVlxtC3pHmXfyUNGwwgfvO7CDW33AojED+dBZDoVYDn22Ehf2XpA3Al12XjNm
+aQ/XIRyP4XObTxmuVTUcqeLn82L3U+KmJzVNFhuGD1kbKr9Ui9TuCXw2v+iAw2HnmJjhBvJLcI/
IJtU+EY4MJa+amBcmNzxfjXJi38c4D0Uew9xSELm5J0dDHWgEBgbl+L5FTjkFUyIV4xv3ydeCBrl
mA+Ib22AXH4bbLgUJP6wMClUsLp9nqjuAowGZOnxoV/DSWG10kPOhvPHoX80bFXNkeGjL+zfMSf7
fOG1sQRr9iLAr9HPotvphg33SrfV/tCO4XjazYI89cgaNiIieoqYBlyLKd2IOzOyLNq7IHo2mr39
WOYBeO/4jbIyuNiDuCKTT5eAR1n+7iUfgMpSzPT/PjM8hPhWU4SCNNZhXcNZoXBjGXchkscTGLZY
JRl+aKLHn4gZOlTZINQFEWCeg64Hct8ijRLbMagM9smzXuvD/SmBNdG9T7/cKaglgObjvGGHbX+d
1XB/wW2xbN/6+mSsKBdPI+YeYb7a03K/mvKJSgt4UimHcDfMq7Vb1rZTjURIkONHHClvC3Cd5bVh
d3MT/rhgi1Zu8J0J7QbNva4XPfpkkKYlkCXx0EVeGu92kMfI0FzzwU38yeORH5phQk3QB1M1Kkz0
oZapLC5LOktDxC8bjuVHrPX8doxpf49rPHh2zsC/HNhXDaZGQhBR8WmLBevosluE52KfsapoUhno
i9mBxIbP11C+c0Urpha/uHO782GPRjwbNGB4D4vuXseJln2DBe4tJwgT/m98YDj1PsiEpyO27mYw
LiFs8aaVP09ad1hKZDtcUQYK18pCSwX5lQ2zgJnRoSouIF7loKKY18sE8PBu4gzCDT0xryaZyxmv
KoSWWQ1uTiJMJtbSVJrtVLPzk1zxyiDSOduX4yD0aH+gJ7Z/GeZhPH7kSsGoGRqumLlmcnhdFSZ3
NegFbyo22NvLMRT7TI65renWf4PsneoxzchxQVJPOo+XYfsvr54Es2GqwLnIH19V39ietH5Bjq3b
bPGnwXRaifjUeCn/lYsFKHtUbwVE0ybI9gwqrBERgcsZRo1d5rgGinT+y716VhC9jQ7zYd86bIUK
NgBRsUGaEbrKHcqPxdxqxdxSrMpkQbzXUPf4h21/Xw3HRHw9h3PH1+ZdxmDCfJjdjc3suJDBp+B4
+A5fvNfl8ExhG2+loC0aT0PTuu20ywZDm1koyL1g9ae8v7PDPmE9wc4WrkhLKeudkeHSF9hsjGG6
yvIsevrmTo7f4JkrOGwOm7r1AO2ImACV7ANtqOsXrr/z4obAoVCHkgZY1LrDzNT7cQDc4mrmJNCZ
pKNtJ4346Chj0WazYRVymAJqxK4RpaQkdKF7iO/JCPjFctAMRxjbYksZhdbFg60a1Psk0Ry5lqfT
v2as9IPvdnxP37Cvi+7N39yyBP8FU7iCQ1mhdh4tazfnYYuv0peOVWC5/vd95Jj/kD/rEExYMD/f
BKWWv9lsio+cG+4SGX+8jqpPv9jSKhBo/dbCTrsLdw49B9BwiX5mO0rUq1pmk3N9AlaFL059QL6F
C88naTwtxvKJHpnoJsIZWnliB6e7IiNQ+S2hHFllWYTzn+n5+ANQ7c+5adEvlKo13W4ZRa1ClCWP
y+iv/q/MQoVUYh1gR+Hs6tA6jeaWijJoNu2glNF1nJuOL9x1kNHOcItSvnq2elbueey2+NpXIXRb
9cCVmAPEc9y2V0om1VueaACLqGQUvcHDTPmxaQT+63kc7xlEXDGjdQWvawO2XXG5zWIjYNhNeMys
DtVaZPN/DdU5/b2nyWKJQgW5Z1IwNriO6j6J9HKfnaaAZmS6gllVEb6Phcnzq8Wz/77lSuEDSZAZ
ipQkvvvwbaDs6BNl84nxR7KrMU6vA3m9AHHeP8HJEFwXPmx5+1Js8biANRs8AH5MBFppz3i5BRZ1
NUwFpMuub/xVLcDiXJTwNDpZAtP9wTANoASniTHxJln910QnNNW6cnbKcSSrC7sPpNcLwqKstGwS
HX7vOIlFxforGouwifQDQqhgjEZx0CWNiUKpyjEpvaqKgOhc9lTCEAhRyxaEf8VVh2Y0pqEZXL01
RIWxLj8jibRJwVr2RAEphZzSuThXE5egrMI2Rr0wJnYwa/OIH31QWtK0RUiBJZmvpIkwRawvYMm8
j0V61Ytsaw6o2+l9E8X5NaSCDvC6ktPpAOVqb0kLU7w8V5Wk40hBmW6Qhbz/HN2P1aaOTHYxb3mh
aVWQfkBlbXS0iOqB9YALcC+9LwmcHCBe+CVYmPyRKMJnPOu/aXFShifa32eupIq635a6nIrdXdVf
iKY1svmdtKOmYN6JQT08b/sTvfFuepAXvqYga08pIdb0unyU/nqh9ldrhD1Ro233z23XvW0HZFZu
Nm54vh3YP5SCV23QPlh1CvuY47Z+kfvMPou5mGn3ZLIby84Cl5qsj+uu9LBcygPZWvW78UZFRZBS
Cg98BrKUjon+xhkSPICmGFrVPZp8lqWctwQRsY5PgC+6Zwlr4Or12gMAEGLaJRGqXgrQHu1421PY
g9W1PR2yyaO9JuojRwwzp1k0oiNctFK1h4pbaz4WneDDUIy9xbeemHs3w/a8RRVAo/EFVtxFoE1p
sIBCAWsGyDgVUSrTxQiA+jLGc3RlBkk+mO95KA5AgJyuDoTXnz1CWR/FZlrYhrMTs2EkHUow29yp
lDKv5lsFAhNKNZ8w70QqvmIO539OxYA9X/4AYk7Fs9lVxRfAK4+H/Gry8hR2ihXMkDRsW46o14z9
ddeitnjSjNw4F6zLMX9oSFXKKBCd73n3KD5I13eKgWvzARJ4wY+5HWgYncIHdeWoY17JtnAe72xS
bXFB39WK9USoHMCFik2aQivrnK3KfleVdkhS9F3+EA1BIbdJ+S0kCUPAajJAnYU8dhOwTVXtGCul
t7ddudD49C9nqVuQfzBDsRGGzO3z1FLVeXGCjwW/B9YgZzoXWMgeCski8nfkLhiw1NYz9/5Z0zeO
6l/z7XHdiU1WgZ+HFaX8elkr4P1nSdquh+ujTFyqcjGwyFa6vTAz0qSa554hdqtWB/OZZS/YYppY
ovDFELrzjocA4aGqMhYNxnKPyZ4c+5DCSslOWcmEjBzR8v/70YRWMerE3GgF+aXR5OT9bobahbdf
CRKd+qVreIE/uQn5IRtaXin095wEpsJKVFqdKNh0xhpazdq+wHznHqFNprrtm9pTBC/j5DkmaEqh
Oi5fSW4F3cLi6GL99b4cwRFhgr1OF0V+FiBd402RfIjeIEGgbzBKLN+aAoUnCsIcQ/r7P5vKU/Gm
CM+f9fESui/oqBAsLGNXy+ZwFdJwGTMtbjrckZHiB2Q4/Fuc/N9OWsmDNk2QlKrhMlIXL/2PZLAI
oUZoidzL04zQfggwjX9HydB1vWcum8AKvq0qkHjG4F8oEfxXpx5zHyblIoFfwvLhFU+FBtkemGCZ
F9TB3UBvlkuTADjiVCEjWh2IWiCZODVMG6jnxekg5UDziBpglqjgCjDbMZI/jW0jBeYbQPR4xfA/
8jCTqoMuWpmSbubeXCbKvSVh082XZVLVltZkgHC1JmXIyo7eLdMd4PhhGHHTzbUutRosgzah2WIB
lGHAaTSi1w9I94xXbnXptq42z3r1ssvcbQZqAxKDkY6D2a8RqIVhbKTkVjjlBFt84S7qmdzvoeCE
DC71Y4juWmn2wUmIfkxz/dZ+NJKMlu/Y1oTo9ngzIIlPIFnIcaSBKd4ikzBKja6VU4Xou1OPRQn8
t5v83Ni11VMryEtyHCn6h9xyzddWfN39HUx1VrpZxNr6JoYBxB0dAxyt5OHCQWpJIOs6JSG9yn07
5KU0Izf0nC2DI/U44lSpTB+thyoKxOwdudDvnXSA64INTGdnGfUT+aBll6DhTLwt6igbO/MRzMRZ
ERSRltIJmSILg19wvkwOe0NvmsESXK7EVMPsWS6GZGzAl3NmqK6teHT1wd3tO2cmsFiuXKOlOUor
JGp0B+ZJr5cqtCOmkwvSEatQqqCgqz79fkCUPz3ARTt243EHdajECLfcrrnATmmKhFFbrqiLHLnl
APWd5eNuaG2b18bQUZ2DqgIyigLysmKBDPF+Wn1fj30ckjtKa7lGaPl8n9xAXBTR0rc5sdN9SXGI
Fk8uUJIhwcVBqhybz0Dt99cpZOCpA7CiPeTzCWQlbjuOu9zVIF/DSMaZR9Y2QU4z/wpcV6NFO8z9
dEmJkeUxM01Om3/x3TJlSddHkdgfuhTF+VTlP6L5SH8JnwVh7Gmzi4IhwXT/kwbnGsozXAjJ739d
ULrhThXQZ3Dx4z3IxlKQxjqgT5mTt35DrtPAVILrXH7Ymf+I/1yGk09wp79ZOVV9YfxYrMiChoXL
8kwi8bsysxrqBfeZup4U4/+Tw41ZQ+e5Lyg3/8imIkb+CVDx4GsIC9OYEBvCoBBBSSZlBkfMM6Wj
GxdAYsaCxuq61IaLeBsmp3hN+Z3gXusE+c294sV5343OXlff7sKb82YFQkv5/kkNokQiyxrblPIc
em0tQeLuOGGQ9xyZRGtnbROr4Ek/NJqLjgE1yEbXxNyjSVzxua6p5THjA83IMJN2meAHFSCHrSzk
D1FxpFpivZVlcLbOu0hw1KILyUW+7zC0QEMVcplZZOCASple1nt6W5rlQ1oFTYO9AtGtBMb11Q3j
1Bx8Dv3AFFNVSd0CohGMjL0e3pZohlmvXPLGqcVQJCWsiGJQbJ4fRkt5UtTKlTVqpEQ7eJtXvSMj
wikb+uS1ggIohnaiLEv7RYqNdGZaLg62FUnXkY7LZ3Kr7/IWzHPq/bHx2oX3hljPwK+VOgv5HeXW
rsIajr48f1rZq7qHBIKckmk1HsD8Rj0ofWqIwe6DMQ0IRGAnUzRfQaJ7J6a04HSzw30w2MwZ+P0T
KZMn3yM0A6LDfsjmtuSNE3BdDDBFmwcURWnvdBwQSaiaxekA8sOAkXJ3FBzhUxdqHqVELrIqyFly
CNwzMxO0/uKDyEg8h9dTHLjSNIMA8S22NYSFNzHrLniKw9fK5M8AwJgcjcujVfC239o89Fl7JrMu
nsIVpTvoDq1TEvTLcoA/OoKjbv4n8pAy+cUSE7i3hqp7YXc8B/QywBIQWvf4FcrRIuKonqIErcIH
Gpd0HHgCI0Hg+iCCYF8WgAJb88DnUxkEg6aqaxr+P9eSynafPWj2jPNoKLDbFWGzGhfUaB2mLhqx
4nc00ovP2sSoQuwmcO2IL91zde46yXmJdJJZucvD+80ZjhoIJ/Kn9t9hMzLkYm+t7mZ1mYOyl87Z
wlGCVTCBqDMzA7V4bvVF1/gkM1ker7zgjs6Ay+6AuNxZpUTLiGEtHoAzgO8HRJM6Th3+149lmBjf
ayRPqTkzIahb3aiFMxN6EefTaGbGPntMPjmjpTym8UaB0ERxi3fPYkgrCXsWYxsMP8vOyBrVXO/v
AK4de4WLLrmtH2rSZYTi2mDEiaivE0zmaaId2OBciprfqQ0nDVPabIIfPzgsXWPQRZW0NCjYyZaB
SuQnKVeRM7eRyvK8gOuVE1rTds54s8FLBAE9lFB/gTchtPs7XemvE6uYFnjzHeijtzojafSSJPB6
JAcfeNPGkV3wYsZqfbEFFm078lGlcwq7/sdAkTTU0m+W2e6C5LSjdNkET0LILFAHsGSXGOmgFrJW
ZinLrVrrahw/s5juj1McKYvX5FXsj00XlilcJK0YXBPxHwwHhOmVH1OH6OTchivJqc91lWn9tIvL
3WC/i/d+CWXfzwCcMX1w/Xn5NTmU4ZId1R7gvOYz+4gb4zMCr9WvZI+ScO8IynboapKXODmK40JR
nhBRiEQfkdx4iwBLpLfUjD7pBuT19XqjWrzeaNYDo9dCPf/4cy4F9dFoRHdCUw3DvEpJlckLso5a
KI3DMqklVLLPdMy0rCkut9Ej0OCHfeoLlpsVt4cucdED+EKzGn4zR26YBWoDP9aMUtUY+qnTzv2B
ciR/jEdxJMU7OccljgGFVe0lErod0bVkd9ek4mUEktN/kJ6LU2ISY+L/ON3cUCFKa3w/hifCm17l
+0wpt05oEnHlbjhxxpGE1X5rK0blE3nXPJrPtRIsMrjDK4kG151tR9nRrdcK04T78BSA1/NweiF5
t2XKOEvdAnk3ci7JS/rNQi4kSKcAc2k5zLmcQlSHkjG/JEnpKo4IQwaeSHegkjxX8pcy3mCB+jKG
w+hwMaW7YO+n2Aysy8uRgeRnWh5C/IzVZ1r1gQoFmfpTwrQXtjmCjuIWTc5tp6gkO0EPupivQvqn
vQOVpklIo3CnHo3kYxJE72X5TC4/ZfPQ6GuZGIG9NvRz7fpzOOs+yO5zPqjt/8kXXiZB9SWBtIAT
DOhO60u9vDq+M+scjWMu2STPAmsckEDd8KpuSthSSVBZKg3RaD5I20EqOlQmhriC8g1gOx8Pt/5w
vBBQYVrCOtIel/njyjGUI3A6SU1LG8kZsLMBWEUBYxs84/0liTuObxd+tF6xzvQgOC0DQpDEBWBG
u9w6fzIeYXrpvzubWRbL7UVKK117Ok2Z+dRDCujfNd1e6fGtRlERj+UqrtVOzQoCRxBQ2jG+Dgki
g7FPIa9HvcWlKqJg6r8Niket0TvWRQiHLSe66Fkot7Eb9DZi3MTaJIrmj6MAph9v3YcDwNRnoVyN
6j012vdyTe8T7ixmkWwChfJ3EW/aEcOLVudAAAjQ07ew+z2FRxsd2fSXVpN6uvGNjpnKMRoNxkaq
bD0bu97sEDrhJBhZNArhYNJZH8o5mwX+cn138GiG4CrJdU7H7++ZIU7ziU1AGgRXRg5upIwSsi+S
gybcjd/pBzM2K0L/2IcU7qlndSW+++fcG/PrsMH/JR6t5vmidBgMnG1tVOPizvVQAbzW0P0dEsxV
2SQWBpmyNybTH3qPNhepr9HBGnsRPwxEyDmJaFOPWXh9ZaFuNjB34dwZfqxX4FhAzxbZQB5gMBqD
zsierntRzZspEKJhys30sNlha+eKRtU7j+F/AOscOFBPQIJjmY9sPf89BSjwYEte/Rw3TRowFBT/
jiaJqBvTNwYirRFkKLMIHWrd4p5Uf1zCsSYFiibiobQI7xJwQ/8MFUBmbiXQmocVQ+CwI41sP8Ka
cBB2jEHPEERJ8BI2Uf6Tv9bPtvLoZjpUaeCJ6Pejg6UNhkoGmSRAq0kb8lIXxZg+3UrkwEahKODV
W37NvWn95kVIZPIGT1gALp2hyXRPz+9h39Q1XS7xO03qJj33rHK9zTs0myreQpJm483iy4hQ7hV7
+vBQWf2E4X4XhC6FrOlw8qpEJR9Xf/63N2/WKyRsW9HS3W8LVY1S9E3r5bstIQtcflCdsQ80idcL
9o6Yl9QBBh5DdeAHpM9yp6JFQ9ySxF+Ir5Vxdl2IXBgMk2iCbXb0tnRPSZVwSOB9ow4mIOWm7Sn6
lOJTsIu+4jHPSPstG1KxGkpBnt6ULP7lzxdQAlHMPvreavP4BtYZz6Dw+VZcPtczymzEh3zdGY0Q
GMZiwO+0Lr9S7992y9VMWbWxEL38d4eQ4c/Wse7ZxF9PrZwo1+MxP65lgHTp7Sax0wUp5m/OAYJ2
YNV3W9WxymyUdJqcak5iM+GBo9GKI0cn9nJAkutf1hVSuQX9NbaaTUO9vmTEPqXsfEYR3z/72mhD
mmkuXv5Ho0/LTFqRV8EwjpIuTzuZ9D4PcYAZS2m+V/+i7F4wm0K7Y0nJ69F0ukukYj+VHn7UKZwt
CuMmEnx/yk3hJF+yET5O3T5XxVR11ed52X43g2X/QkSp/v/MXQkv9FHc3/l9uYZl22qeC0dztgCw
aaWZoW92eXFJj2xC+RCpcN79pYVKTizUcijNI8h7WPG7ZcDPufXH3Y/zwTn28A17dbYQoAEMIwrd
RkzrXv9D/oZ3ZauPjHWSEdOaUNes+lO8q36dn89103oWaMkWc8hkotAspz1rKNaVhjL3V5/BzTRy
/ReTMUApRxu6GkXCZXBMQi5PoFxm2k1jp6VfW8FGCZmGABfSfUtMpqKCYtWiC6bJ/xTC7eo04THO
LSHzaF8E3jnLKmp2tIlx2JHQo50+ylQXZmtWP10yv40mvwfYRFqDXt6NlkWuV+S4MYeUNSDNDTkO
MQkIlzR/QdICONH9gO38J89I+glNEct1SRKkjoH3W3O2G00wVpBa0/4NQmpf+RqQRypjONM+WvuT
KLgEG4YlGSUvFBILSiBEQQW1+nEP0B+1l0NCe/hLUCyTWmjkp0dVnCac4m/eNTArMnW1mYjdIbLz
fekxWIQUzZ09zT6F0jPRvR17ZeKtHjNLQSYMyFVa1yeyRpX80YXCG5OPV0fdAp4N6uvQ4vbxU6Z7
vbSzQsHRVHgcifcLJDJUKJSeXSamRVoZHfmYs1Bq76QuNS7DQXRRH/rFAkwgMKbFT2A/dF3XoFGB
Ac9euby0m2VrnMod6UglxHjzVrfB4NSwAWxQTCNu/LBtu87Q8cXvNriqYHCjx/7u+53cggpbdk83
Gt+Hn/I2t5Gn3upJtdpqBA8uXeqNyo1twCxAsgxlVi4jg3Z+1zDr6FK9RoNCMysdp0dPc4W+xXe7
kboOHgpT1wmyITEeUeugRgFmbcD/TtuxBsB66+OTRtWZu4NgURGFfoSCRTT9A5lXLcI37Xo701zN
hhy6R29enpk1dTiAqSCxpCbjzkgu881/LmU+SbLI2v5SUuJ6z4tCi+y1eSM2yEBAqvtD2iDHZpxw
wj66tT9qNcVG2cxA/Q2xf8I/PB+RcD3Wq6ta/eBsfNzXimzrKyv72pxipt7Qj/0slBxnFdUNBevB
ZspNHF+oOofoOKMxzelu5JpzaNyA1dm2mefSxEd+n37nu03esric/5bf4g1VB/C6D/qfEHXHqEp4
76VMu+nWeennWYQN9cNJGspBfA5ISFLbeyeago2NS2OKBMkuuCYm3P51lyB6LS4AYr4A/iz9vh5f
aJSoWFsXy9RAP9kIenopLX5MEURJFgJRrupP++jIC4MImmKzg/auYfvsy+oEUG56CR2Bf5VjujFD
djlWiaEQJ90qmpmlvEkozmejBWehxihHjeJclzqO0OVFGPIVarNx7H5oaoc24xIn96WPfaYUVeyw
aB+hbaq4PFt+DJKhMV7tnASjjA+6RFpM9Onh4HrPB2Fvpaeaqyp3299qATqY0shLkmiCtvmzaEqB
y7gHYLsAaWjoktyhQwF1t/mkdt4dDX5aUfe/CPqqtNyzUOxm63IL5NAMBfNIfOsO4Zydck8GO5J/
NuCmThG/6YYTkmAIMU5Z/KtiLwxNXrNVv9VU5HwCGjsAEnZzDRM4Vvq/bew3VikLkBeUk1yKi1/W
QzXeAcGFHa4HZ630uRxtXzn44xTSwLoRtTuZtQ1ce8+vgnC1BmYMQbIxxJlDAz7v7P/ZYefLb+Hx
vLL3lSEey1Fwg+3zc+dzWluB/aNDEFMkR7Ks3SdbBE8YlaK5zEBtOhT9LAhRAUUMdBeT/jt/8f2w
puXhV8GXoE1vzSHsjmItBU2rkDEMrhJxRKckkwJ7bDW7wViOxYbOF/UThYewT32wm6mB1YsRaSsd
n2t7y4PVVOHQvXXol4k+NRpLcA9pwlxNKfKOAWsA4W389BLaPQlSoRc5fBqTTJzituc1A+gD4zOa
S0QUfb4DJ56AWE6buFp/ZzCkXI5Gg3ODg0/8fwwanEb2Rx+/c8Y3uADNgtoTMALGIdVefa6voG18
aT9xlVayGZd52lYpNw9lzUliW8LXEaRQgJoIKylp8vGRZ602Yv/ggCGzPDa08tfsxxyewdnJq6cd
l6h5HU7tWazpF9vt2yLt7lC/3P8XEYi1S0yQHQuZ8xCzOIL7DlMwb1bGpL1S2rJ86wGiIdOpSoX2
mXltX8XL9Rz37Xf2k4Db94aiWpQyViCmNsTrKTd0uhfPHxHp5HepT8n2Hp5vTpsham5GY53ip+wk
jCNQ6WkyYT6L9w6rFhdNp/+6SbzJ7sbY/JVn2oMj4V3oDrE7nXTPho6rMMF4ta52wI3fPGTlhU5c
CjIXTKLA8TnQ/0yXaLmPDR8tZTy6nijU7wKId3svfwmx6l2j5QvyjbUDSW1KXGlmOSxjTr04Kun0
ffCiJrWVQXUG8ZHY7/YyT8MBwPSMiqYwYFZ2WD8MbOiBLN0Uc6p6JTEYEzS3yu+s4YT2nwwXxWlb
WktwYinX9nedgkn0fQBFJ4nLEoBbUY+LTRPOoubw3b6yb6FC1RugTSIZs41s/UFLl1mYB7WsrrrY
NJu+c9AZO9ZaF6QdYih61Xe3XR2P3CP/V9H2IOlPuKaW0uoljaItoZbkBk4kRmIeReiobShfdbkk
LC4hJrP+tkKpHVtxataBugozXDcKUdOgzBr7eIDhlgv69DXgOPbVUFqE2ktUrjPbARMWEwrfcGX0
cLCNAGrmYamsLAgyZtiEPZbC9JhHG7C6274yUs16IoBCf79FgHr8pH7bJurP6+5qCzM3DYqnxjAn
pEjmbFz/DENQB93lPcPjSfZhluaNKhUIbr8zk6wsepUfE2XodF9nEI5dM7al48k1yvMZ3unbcHUu
u7VD91cmK7IwXIpt6z10689udEg6ZE7lQ3iZznHjtiEkxfaEjWDueLBPjit+prq+Q1Yga7GUAOLC
of7AK0HIcV0qoHJda3Tla1UXyrNcTZUS1WXYTlu4ybdbENsWkqLnpivrqm+ELhnMSeNvuDnFq/Zr
ATb9uRh7ksDW7elgr8EEoaSNHyR4J1mwv6s4CwJ54ZzkzPaBP2nnHVBsXEuGRnPJgeGOK4YQerRg
ihykooRfAbKri7Pg5mmvxZ4v4xQyEGdH8xwXH+MNdmNzS3cPK4C7aCi6lEr/Smb3bAktaYNF2WsV
+vHv2fwoonsWtfoH5t6M6/xLTqu0PT7ioc7adP4xf0Nl+4rBA0MrhRXFr/4rXs+Dqpqb0fa718vo
ZCFfLqpGuMPHpvc821uF+T04TAr2Sc0RMRseGtawrzJshsNsobmCgcCFbFBcVd0i+Wbczch6reNc
q1X9S0w8JL0CIfnpT0pI5k314VrI8KrbdtztmrAoTtr/F6i8OyF0s5Utxy+pZTj2E+GuKuNq+geJ
m3HRCsuejw6xEZ4bJX0s5SKCrAM8tDr077VTYptosZRYG6TcyW5dwRASTVNeQFhBCufSR8z54NHc
WApbVXQJb8BSkCaIw6n4C0IuHMbII8tDtJOj/q4Z1KarWSWRZv8bFymHlYH7s6G2o/WCMbGIoSlm
mMqvicil8Z62iVJ3HWDcGOsRsH/6YNBFNdjhFKZ4iVDUe3IVWS001iRE6tZHfM/bbjK3wCxnUp53
n2/JqQBj05QVsl1dn7T7RKTc16yDSQAmBwCtAHLfaR42IY9ABKW/eYwrIttKEcQaTSlg8yp+RBby
bRw01x5sQyMjieGnLmbouSVybd6kznDqT08TRabXD2CbVFp368Xco03vrXc1Y7yNgNeKoKNOLwlt
903DlrOjOoMtou5foNCpm94C1bvdzHPMR8SiBer0x70CGtRHBBK4i4ZySZHm6wlde8Gqq9Zf5Vwu
QBgQG/6cY1HRWKA6HWIZECy5YWCQSLk6fowVx7pw5FOYZtJxoYKg3M+ooQxEsrtL9B43VVp9KVeQ
7PoOXPsry2UqIsIYdgXRr+2djOdUQniWEFNqecdYNxdlOGcnNy8NuvX86ptNpwWg+J+46wtdaslr
z0ZkfUx/UvdfJ85rAnrI+UOw1jPZaRyr9bschIHP8eObJnHV3txKiEvGEaa+YhCCKuk/+lFO4gYJ
okT8SzVXebFKxEHaav06+vVEr50lLjyk603PiVjrgTgRUz3rg5oCbxP2RJ6s+Bp3lMtonSfXD6wG
yKuJbHHIqumYbE4trz8gR8xV5l5nl6ys0Ig5ea1KGeaNNQjRz3BxeCD+znNCjeYpolUEsEY5nkTu
8bFJNTTKAtRaWeOao5RQJWagfG69Be5++j8EtbdZnOigZMRkgyeECQfCkz9CvyzkJBITfxjYP2Py
KzS6I+5276wa4iE+oYRj98H22tibKbOKIWCZrlXShy/pPh1UOhPiY16DSwpgekmYfLV8CYE7yQyB
tpKo9dqn60ZDTim1mrsDOMWOlPmIWvd0GHnRw0cHi2m/6ZgnbiqhvPS27cu1CtBv43Zq49uaBe7Q
wtiLz4f4PPQ/rZ0tYv+rvNqkquKJEiTdYo1sVmztlJRDC+LglbAQRrfh+uO/ZINSs7bTDQf2BMPn
Zb/h5AL0j5VlDnGLgtm9JQTS0CLXebSCoYWvqnCKbjMaRxSRbentXJ7skKn7AYsa0/kWUAVfwlxX
faHJC3ftfaKBqfnOYIhGhwF1ENRL/9IM10jQ9Vw69H6FL8BTWv8MVwvTUL1VH8ONvDCJKsjCAtP8
zzndZQliRGUtahN2FlezObQK83wwHffZXyu2gB4vEcHM7dq3SGErzC4UDgHhmv1hzCFDjShJmbWX
sMFIsOV+dAmYNQaCzCyr3c9ygghiaBQpByzw6DqSyc2g7R1kgOcNn0QRRJ3zYni8aHx7QBNHuhRW
xqwGoa6RdW5yLPqmjGzpcaYBI9WeJkMcptUxamMvRMA/zWE7jDqy1g/k2YZbiBP6rInMxmWT60xT
wqkLDK1lhiIOy2pLpkSa48pBBDv/zcPvHRnA4vfSk40aVuEjDYDWezimO8zBatxpqkYzHcMY2Ukk
bjXpXzbpy/TxX0hNRWgKU/SVETbwsONhAhod3nrh2bdEqmcaiY0dgtKTUSoR0ajsrdVRLKRU2jhn
TZfN0MLG46yEjqUb2CuUj3UVN89CRU8lyN3ZnIFGG5fBfscqpV5hg32Wm+lZ/Jt49iNsLCebVFxi
9Ubw4v3RT73LufkRHciDHyikbgC3zyREZiBx+PzGErojYcNcO4fKpJao4CaKOpYcENlFpS4uYtZu
sCD3/6UHh374IkD+Ba5bgnJCETzYk/2OGyccxQwwv1RxoLTkVpJGXlwJzmvl3rm4bBXGg8zC7L7O
EsoGLvD57SNMY5KxzUqWwOZkUNM1ZJdOEIxZ4ibFy2a28E6MMJOZ2jXXa9VGTOWxxWh3bv1HaILT
8qU2Z6YD33IoZBJEN7R+iWHdR6XjaK0H/BQ16sz/NEoK7x8/XHWuhfRnQhsbIEocCbAr1MkuNuUl
Rq4A8+8fRIwVGEJiRHYg3E3zrZdsf+/O9VIrWAzZjDIpyc6IA1TbbL2v5mLmmGRsrmdZf5ds5tSf
V8M+Oqza+5A18V1RZsjqtJMPSywyM2NTPFRx65N5gEqIuPjnevU9HF/c+Ds+5Ca4mBSZDuB03AJl
eD9hSQw/HFtmbq3ycio9lyqfFxrY79p4wtQfIM06RHnlCG2ibsoGrwX1Gv0iZVPWy0syfrH99DWw
ry9/Vvw4RNtueFRPffFUQienXvuAVemDD0DX8wcDYEHMEA7MkbMqxELwDefbeFKwjamkIqHWt7Pz
S5rr64+o1ip8b4WksEWtyiVNo6ZOcqCB3kIgkE2gsvFiQzIeQ7c8BUzXmE0zPBv1TGYQHJF6DrV3
GPdpSnagYUtDy8LcH3+aB4Z+vf64SqXu7qWt0mb+clStTXqd8RCD4+/fbu+vSs9isuo+Yw5yg3ID
2EDGfgS1aJphLIfiNab9l16WjQMgV++7u09+tvKUQsuHt4FK49U7SwtpocFYttAwLCGZaS6RxmXZ
fu7rzmiPN85m6XRQ6FSjmJHK9BkjafuFg4nzVKqkzc3zYhtW8KKqR42q+YgBI3f/RPOhulumPoL6
dEq/Pt5BQd9TR6VOYx6Xi/in/USZK7vnm//DSkwU2idnV7elIig4u57EQCqOg+IJHAwqRN1bVgfU
BKQWSwkWQwvAVwuOwzTOvNv87MHCzyaM/4+QFzQ/nod2D5p1oCHPh3XtLMGjLPS6vwUrV82e1nIS
NE64LZv3dIUGX3FFSnHNALfqILenBo2Zm41F/YBHuXL9dXUIuBZXypTpQ2EQ71DdU1M6Oum6H/MB
EsoaQBzt2ZROJTfv9ODpcQlwmd6dWwpQSaUtwbhGBGea4x8LYR5L27l6avekuCi5vHM9pZI3yST3
Q1YMSlGhrKo68/2vPQORwid6Vm3dp96FJcoBQ4n1/8z5AQ5BJRuOt5gJFakRUiJVxHcGKwhciHhI
9dBG9PTkIteAMABllAaCpkEXZyGIp7DOE98ZSABaVoPJoNkk9TTszqPU9fP0v5iwPsSWCnu90gkt
7Ueci9it7+JB7x7XsmlM6DgeuInZub226cmpvtreOqm3hzb0j1NRKo3uG+C2kDHFUIqhbH1LXweH
2InYR3PADwCPEG5BmH9Xoqfx4u+gXYuNEhIiuz4uT6xytl5Dn5wwpHM15Mchu2EfEhOqHf5aXH31
0vUIkBZyRhgXQ5c7FWUqGIxGtaUqzyXtKiGFH1MhhYvnlLFgenCv7UDgFFH6HUPwLFyxaaGckace
r7wJLee86qcxmYuwbIsZJ/X/v484mYV6fITW9f39XSNuzhSWjbOrKnxP4x5aZVbji609u1j6NBi7
vJbibphTbPIcV/xocXqCm1QD4jrqX5pyZcQWHVtZ7xfDR6OW7CPsqCq1LGC97i+V3mRF1Gc4r/v+
kuVt938b789WaTPFzfVLf7dtc99CCUPmPIJ3x5t++fqabRsx0ysNBENhD57Q6NAuTLcb9cndA3y0
SUS8ZEq3zgqqoQwvHTdoYx44EnBw2R41IMwFOjEQ8loP72nqg6n3PfveSbkwlkNLTlgxGr0YtvvM
sHhRHG2KFyRjnv8IpcnpXlv6CJcAN6F7YbA939FoKp7t+lH4z0ik0s2xtfecuY2oFO+3uQ9K5cW2
/c/PpSdG2yCS+CbSLPkoQBifjujugKI6wvXJFmY5dbiXTBAokCbYbNlO2KN/p0aoVMMXzW57Gxc5
O5hlLvJXrCAKhlVfe8JZcMc8Y9zKVjHBeEcIqX+G7zvH06ruZtTTg6r4KJ0xg+JuBbzUZunXG9/Y
glf3hw3KZC/38IZblQu+41WFsu/yG9FFaj6kS/vKrxkLqZl5JcMSOMc70SyhnJJspy4sqFpP658a
6U6HR15w/QOT8mDDNq4fQDXT/nXPLFCRanxDApnJIK9xSS7xzlgfjdHbapn/m8icRCq+nuPVuGPR
AIR26yJnLPDcMafUcbSRNac0fdkyVIiZPRQwgbXiOcn4jkaH4I7FlbpA+YBfMn/rajdlXst5vZrP
kdWQSRiED2eIULbSlQmFVkU322wPNpchDMxCfVyJsX++AWErOfH249lFjIhETmeL52hLeSkI8y88
+CWsnbntl+5jZY9ukCWr0krjz60FgcCZ2zuWoZtZW3+dQ+3HhYK/JCz8rT/Hmi1gcI7a/Vvz0Re0
3YXQu/PZPYVs3y5TRqCPoz+jYFkSiTkNvKH9aothwxtRoYcsM41NBOVXMK1zkWAXFLaTDIHtiIkK
BR5jIZLzdqhsC85BUQR6BHuJqSRCYH71HUU1XIrBOtHjGxwjmOfPDmTzy9VIkrOgaV/HMOXpRpBv
Kaf1ZSXyFfqu49gr17k6Wq2lkiXDh9tFYWbcc0F1WE6KAKyniKN3zSD+oQCBGgufd6D7U6CGX8Ov
hkjvRbfhfP55FtPk6awfnF/gIwCd1kSGp/0aMWDABLn1L90VYVVZMVL+wIfbA2anGEEXwGVcGID1
wrMBbg9IeW801qlkh805obdxkKxnut/fm9s09y1IikBHV4YmOXw1tos6Q4KIxC2dUyeTKyzOObHv
AJsmnKs9BBVF5vjoN2WOSgnYgMybkW+MouNQcK4BLpUKpWnaVDnxrrqhQgoBUDaYWz929U2ZiWRX
NYFBiGROMEAh9OXSU+vB9chKW12RnedU656vYAuWgYEE+xlESECBkeNubi+5g+E7yYLaumMoSRA1
BAZyha09JkoPL8vhIkMA+uoC1xsl9si5JoASCGUiAZYKyOe9ysFhWInx27hC4Jp6CzjTvHfdDFF7
AXNAQ3AJg7zVmD1mTuaB3/K0G3vVjufaH2jj/riMOpHVBkkW7rRpi8+lAn8oPD/h5vHn21krmdQI
5oY018uWIAwXkIoxeThJlkM+OtPSKHaHiVJzwCEfQoin3xR5C2cituha3ryjSPcV/1Tug/t2q+C7
MgIa7FlJF7f+JmUM6dNwlv/LK1Wzc0lIIf3IBRiV0YGar1WmdaB0HMoP5sPuyW9QXnysmCnl3bS0
bbUTLYwE5n6mvQPxl/qvq4oOI4ajI5r/hj6Ad5A5zQ9CQUlEHaRkk4peDKUo2qJmPNYfiyjH8uz0
V5gDWXqyhg5Z+Mu8xVWPh8m7eMJzr6M1mCjM6IjRGkfheCwDU8mGc8CKQrd8e3miqacZg1XTewhv
RD8LVMinhvRg0t3bAr21wex/AVb93jady3awPUUQN5Y1e0H0ijlIjfFSo8xGK8tKNHB3JNMlepHc
LLS0bzKo2wjJtaLsuwHbWyqQd+GqUEPK5FK2Xdpc0RPnakj9QiYid0DHfckGrT9ANjf0IIBZ1J2w
gZuHuSwSCxo0Xqqqgvn+e3Kp0ciEZygSoo3eAgfbVy9PUGEBRkg4mZGrakliAOIZIsKOnBPseoWE
GHxhsStcPZxncoaoIr23bIdomHu2BEm0avQwwDVoLAmhjRXfqJS0lVDh3TLGx3Lnw73QZ97FGvve
vkMnIoCsVDV7Z/7gR+dRZ65jLTbbYnhd0pP9teRwRrr0vWkn/9DrRu/meHko7mHovxDe8YPhh9kB
iiObVHsygJL9twDTQC2x1sXfomu/98DZ3PxBxE5UvmrZtEOWPYkTMhup2Vd6MXc9rwxFNRVj6BUa
cP2bkhfobF7+gn6mVS188mky/H4x3kd7+F5cLhahgwXAt1vKIskh15O0CwTKPoMvJSUrvuL2c91g
toGEkW0ZoxR+PqJelmsUqiXIDL3LDtfvNg1FZjd9Dg3x9UfZOmVHo6hFxeVxQtWoPvceqRwD27OT
SG8QXbs/GJoDgVlCRCYG1RDGe+QOuXUa6CMqDsRu/2FAyvrtbl8zMtXZTEcKOADmTMPI3LK9+sMB
0QhCpn90zRMBPAbtoI72HZ9NBMT1WhrhB8WiJcgB+z6IMBAwKvT+22ZTnYGMaSVgL1fV73wBEkk6
dq0xRbN54ALRH/El6wTrxwPO4KbUJSJpPBm0F1giCDkCmRZ319U3dR6cGqm8/npE1MyOJuLA5NKj
XI56tSITDbJw8yy8k9C/mAVXuQfLB0kkfB2F/H16ZQl2vSUrEd0LfDpEY5z+1figNFKumuIU6cWF
sT017vvPdbre16eL5BobnpnQDf3HFooA/qKdBwQjZ02VS88WA9I+K5QNPVZZE9vz6U4G/DGg1jvm
39nbEILLweUMAYPV4wr8sYr3X2LntbUOjNfFQggh6UcE74xM5QwnfLRD6txEztC34RSgiyHup+dh
2IFqiL6FmlXcwhYJQwYWQg98cOg4kfK9DDnsu6IkH1WM7LslEL9OTopBMHXzOPUJVkdeOEc/Q+d3
hcQB9H+JexS6odwxcXum3rzFvZ45FzA9gaaWLEJt2u3njTe+ileJ10xClFLz0fz7qKIA69aJ78Mg
P6mv0+OYZYcVk8qZ7ixkivSzYHhbtAm1Yh552ZZl9vxfA9QQS5+4F9ZXhCHkwpgSfFka9vrG+IxF
kpQZ/mxCWfCLCeEg2Jp4rI1Psb0zsyB2XaTJVwCnxAMbsGFVbs0T+TpCJKfdZaDw3tYbJnv7HOuk
lxj4CTX4TkZtEIB/ObEpYRHFHsPTG21Q8ZCQRWSiom17x/EprI1fFHBBPhUJ41AenR9hHWLIw48D
mIcbBovRlNLRWfDQmhzh7009VWK8HI6jYAsSY0z9K5+x5oxY9G+gQPSZ4fXdBt3JOaL1pzKfB5Y/
9Por6EqOFHOhJd3A108WqGjPJkwv2953UvNDdhQVbYy2itNbSBJS9lXdGJrFKwxMUlAB7WeHhsRL
DIyGuvOqyqgKU0w7TpjqCMZhD4zCl+nPdZ5W21eHFBya0Hi6TAnLvQVX3gCKPDeJu8Bnhmka6L63
fQ+gD+WNuMNjfo6igKzLemF21iSXzWnyZjXzYpZS2d+pQsk4zP38ahl/ONzqX2798I0K6dWDuzym
eXWmOnlqZjA3S6ng1lZ8UJPR2+f3g1QlmljL/H7PGjL21wtUXIqSNZS4hF1mAa39S8i7I4gmtIDk
xjjKZ1ZXUgVGtRQvDU/0mDddUoK8VjFadTXBPn0YMO1kNmo1z0gPPoFLWCtgUBhx87FcXOBa9zu6
o/flbGpvRXH4VBQia9aDGpCsxE+UCUFlveoirQa6NdSDf3Eu/3uEautXeRAWg6kyDLlfN9ws9ktz
cfB0MwjQxHebKTll2zvUaPpUIWBVav93YUZZl/fdrlyaR4t3SzkkxOjFpZ9RHhnn27YQ2uy7vcPU
F8TX3QhP7vSMTPyYCIFyK5Lvrln1y5A2YonmXlCDH0Bh6CQq5MvmN+rLjIKSbNi8u7tyKPNmRL4P
YQ9L9L7BKTSyfSBq7P1tp67AvRKxdmQPujVaU0BolEl55vy6mhizSioz7CldBb2FYEE4UiGS0qnE
TDUMSVn217lcA+0TNGSb++9snrxETi/nymnvZxNlouH5WNQe7HMbVHM3k7emRH+T7AdCPaXVVFBJ
qQIXD8Sa6RRiLgGiU+tVlaZ9mbwmshw6Su9PRmQLQg/b6W5OqdWAFnS27vxfSPRly2yeKjnx+z9t
Iu0+MUlHe1agIJBHOHRulYS+Y7MaVpDwkLFPRZMVo6dh/XGtuS8q9bpdIsjnrosh/sKm2KwIjNzR
pGEdVl4VKhhQyX+JEFHkeFYAa+j4+gdyB7ALo20Ax4W72Huy1oW1e3un9KeWEUoGYxzvbWC9JYeF
emJnMn19fuLSTP1r45NqUSbTxDZLaWa+KNTKf1sTe1Yu2tvsA0FLVPifjEYViTJdv5FQbE5zF/PG
IAN8kHosv6SQduFDV0uSpkiDmnNR8Uv2HwZkfS6qTO2TErK+ywpCaVZ6ZRJbQAQag5k4tJTsb/6b
mogdnNKtIRiS3tPaO2Rj8oTMaluqV/hAUqGG3sCL8iUUG0FzJjaw4F0x21kpawSVdQ1kbnrSI3d1
SJnmb72X+nBN+a9wRfiPgp2ZaJZVprKQXhdvfdYnwnHrtf4S3hw75vDSQt4BIPMR0i85pWxWbkrO
ZXG5Yf58xj9we8lU1c9W3xYEikPYp9Q/gOK1bi9WiRj29QH51XDJ62XxuOpIoQFIRknBOhPQee4s
QqvDweihHuKvQ11XSeAR/HAIsLPfh8cNce/c8qNpIpA7n6IqWuhYZiOfX+/fMjIY8FrB8KtC6l5/
QrHnQGZlrEO7jPtLD1iL1Maq7zK3OZVddW/xO2ZF2RCZbqICdt1Pf1j2Zh24lwB0Gfr1cGxZF2yQ
JwgEfUqYPElF3+I+5V6CsvihShrMEANqQGXImoQEh/LmMqKVoNSBejpua6BxowsawYJ/ZnQ9dkg+
zIKWFkKZEK/XmnyVmurZU63R2uGCLlSehVpmj9o9wXKeAnhZcPJ2o5nsgRs6RELkVF7iu5uVF+7e
eC810oHAXm7pbct4ke7yOM5Q+cQlzvUvjK2BDP/TKfq5ztYqu9IHITp3w7XTgVhPvMSCAvLYu1Hb
Cci6kX852IoqPq6EYWNX6mCDUMD2IBel2oYX0Xbb7KlPdfpKaukeJjjcefOy+ydLjf7B9jMa24y6
6F+GSB0b6IJCwcHViR0L8kC7x8x8eQRZ5QSJJrFx09gSSGJNu0CLKY/gKJ0XWEsjUDCHsXj2yRd3
FMijsebwmuazNcFscAy2O3XpgeJp5cEaakYyep165dYXjpT0i9l2Z90SczKuIyG4mvI3PtnBVsUa
b/sOsl0zPBuLbG/r6C930ERqVAAh3uQ2MFV1zSbVRdjodxJ5dOYB0nco0ar1bszy6nr5CXaYnjPE
qX5c6grGwmnwR0fLN7Lu9jEJoLPXs/SI+R5VL7iXasSY0s7LcLwRX6GDwPHFPbDTduo8RcMsm6Pw
ywTJUdv9ts9D/suceoOQpV9d/DRKmqGjTikqH/gkaSM5O0Ek94Zfvmit/msGl5Nt1OpFiRycS0If
f4B4jPgZ51mHc3Wsy+MSFHyGaa6ilIv+EyfA9RZ2kH3/fP6qHP+OTVBe/sqCvf2NkNolo/SinzDz
slLkWIKgAk2NdBNCZAyHGIoaJKzY+NbYV+AmEOr8TitcEzKLMyabc2so8MAWL3Ud1mLRJl25KdC+
Lf7zVAlJ3rhzwuRWN7pvKzqtv58Bqd6WfyDM+R/YBg7a40pZXA7M420hLWZey7uNa/jEO5RFYE4l
In8H8o5VDVQWY8NqeV62/vtl4rc7Z/QwbA3WQY9DzzzAWcNfuunfBJs6/rSZrId8q4IQMdQvISn9
HWb6GYVcfmoxBb8CkWb0hctHMLv+ovrPMg02o2w9wjgJW3D0w/sN0gw8UHtuG2WfLvgXcmOgzAOn
uphM3ZFQxrwjLlLg4b3TVIEwpgOvyD24GYzJnYyPeC1FvpcwtDb+zPNaxJaRUGKjboMFxyWcrel5
SNSoULSrG4z9GDH1KLV+R4a6UJG5XNgSe5PJDi7OqryNxVKuTNPDYZWFp7MoLGIYcsox8317XK52
kbNlEUvrIRo0CrEo/p8bUMa4VQgQiZSNtl7HbT4vH3C2p8iK1LZD8zYk+3hzTsoXV9vDOmfcdVXv
UE3wMnEWJxU2/wDBMAppWBx9gEQOJWLV7Vqie2IvM+WVOdxeqH8+ehWORw7hl4nJ9INIDmj4tjtl
GnEdybAkIkGl0x+YS/vWd5pgkCiuAnzDV03SSmI7eIvXOkPTblYOAU3rDdr9e4UCa40ipJUc219I
8hkEv3YYg6ORDP1sRH32bXvllHBjqvLyEZa7/K1v1D6N3G1XPKsOj6+KC12c6Q/3FycLg/qaGUa5
asT3sBufo8EyVg/uIxCuVggk3TstHFiVZEgyLeaMzwwvYLbvjCllg9nSnSGzYQIKiuqBLqOgGkDW
LP9lhn/OHhyD5FPnmqcfjpX1g2BEK7kkcuy/AUJV4jImSVy/Z1HZzFawP7lVnS96FILZcjo5EkZN
5HWdWujZ73geuwICHxzzZN9flni+8zkM1diGn7bCRycuxDMqcU5ZP1zJ29pL2uJY363dCYhuXsaa
3CmmnhYPubd+y9/aodOrBQJw85DDitMgh3FCZqmIqIlPDtNFAauE5aOSQYov7P2I3LUCSGhJ5XTz
Pc34a7/lFjor6mdm47/t90YzOWNEgLx8qXhfCE/4CK70zUVRqZjrr6D3yANnVkTMBzxA2Q1LkV91
bW/QPVCtdkblA0qXzgUJwMyc2uGuvNeMI7a5J3LbIXTRySYcorWmYs5wrkvIT0JLnCopg6iU7kma
lGTvE0bbLfzF4qQOrLBv6yGXVyn3sORnvdoribF3VFF3C6U3h2GxtF8m+6832D3QceY+9UIa5c1k
H25GsQeVtcuvhTlYyaz7VCm075wD4dAqPRr07kjSa2NLaUouhjdqLKdn39quRKegXpwTxgPIMQA8
NfWAPx5p5frACPgGr0b3v6QUrJX3o7ewKfgl7D+ZD+Lz526TMWXXyrKZofvwMOm2TSFyxBOTgUyj
FdRqI9nfxUpRkOVdpyZN+uHpw3xi/j3F/qq0BWKhy+YypdtDXOuUhnYUqUAh6MjoIcY9a7bJxh/7
R+PzehYWVHVbdblp9yT+ZPWVZhirGP8e7a/EOfH9H68K4XBLnn7d23OWdzVpn7TrMT4IzutyX7em
r5sefAXx5U3zpIyhUg6RrZEXXT9yICNC3i1tdIMAyMiEcSVVIReyhss/87lDhai2fjox6y/rv/dS
0NHF/wlDXMQI54OCJ1t0j36odapwTZCkHbj5r7DTeQAGuXDu5E/GLyq03Wxlq5wHOQ9y+p5vg+oa
cLJ2/8BsBD5YKWwRzB/em+I7mM2RUWEvLOwkEpSBc5iaYvjzkFueoxVuY2GdKkpWdBGvlwXWKITr
HT1fWQQ1+TNt4dd1TACgC+tcPRVUsxcHKRoFi5Ly737kJzR/bRc1VCij1KBqlDjhEjNJPGNKnD3o
4K7PrEOG4E+5+o3KY0dYq26vQotd5gfM6DIrTbqs1A1h3G4j+I5DcTq2aLu69wk1vghEifUqZYVC
sihauI08n2WnA/Dz3VPR7sZVuyHUaS+GYZwh+f9ZCbOkQBL55bWJ6fxIgXpOI8NTQXy5w3jv1Ew3
oKcrHQDVJMsncN/mDoZhsD33p7Dr4lC9Zr5GYxifGrbSjprl3ilYBOITmAUyxcqq5EM0+Enu72r+
TOBDkvUMhJp72juM3kEHZH6A6lGzwmAfcfQNkQGMx4MPuMdBYqPpOUEpOPXLxIuzUIWRpm54lFVG
oNeXgCJ863pB6t03VGtB76Xy8uf3XuLkS6AmeGj00MlwkNcTEqfYuz8oBS8Lh1SVly7ymk1pECPf
YK/Gb33zO0i2Xzeg9/rpRt5DmwoC3uNQNSUrzDJjxffTzrVqXcum5RRUfnAH6eMyPBsaJHtPwaKh
8yBY8rQWuGAzRFNxsbslEschhHlrbEyF+YLAhApAKVy1TsYQiYH3s1qV9vNMyMt5Rc1xSBgtYQRa
tWZqAcJo7mu7OJHl15rYMsvdiNtLrK7/fwTcQp2n765z2DCtE3F9YHkPPRA9i7IBHd1fQWqRRMt1
g8NCC3bIwCC217TKu3w6Zg3f2MXbWJChXA9XLHpp0rKnVIKoE1fe9OxxJqIcMKIehmM7WAvZhMJK
2vfUv/zVlAmcc/gaulqiORyVbyhR99uWBSNIpJuyVnr56AhHyGqnM2sv6DnJHAJW0n0s3DB8xeOf
7mPU3OFj23V4YcWQ/Yt6nSa/9u68R95p3fb41ImOiS1jy2YdigQy3TXRi1IcP3qridZZyD3bSOq4
SCvA0w7pK82HxnYCb5I2iC8kCNe4kcBOPonLWCXHiTaPRzFcZkLWiS2fu8k4/pSNmlybqWWiB9H8
7Sbn/j/zeaxq2p8+Xg4ByQ1/NxetjEtLPORR+zxTqUEjGtreWv/1UsUbdS3oGHj5bWtLnf50qhHL
sQrIs0o1A3kRzQZxNd31dfUwX0zHX8HyJncKGndY0fRvWJYg5hktTmgcRi1LrbaWqo8P+T2Nqjxm
00fMlGMDbO/+VgZrW1Xp3zy/kagweXWYieN8IbYwuWowilNCcv6JX6zo9oayNamig4COV3X5Tqq8
8EGUJCtkdryQk7oOhSVTJDsl0hKYeplZrvMFadc96j2wZkUIZKJwTa49PqcBQFEgwI+LQYsYnSk1
YbY2Zdg0nbh7yxSPTKdgfIWh6a4SZoXBp/zXSKZT/siNuXnvRM6pNdGoeylxc1vwRsist3ekDUOA
gs8dwyaMorqDrl6eLJfcC97I6v83qlfQ5m3zmyXPEdz/W04HpqM2k1a/nep7N3O9yxGtCJpZ/oni
MibdS1ZkTUHiN8HW+l2SfcxQpwZHpQt5Z0zjQaE7RV+1yTN3d5mlqAvEAbos8eQ6NlKbKnqOgQsP
ax0zLrJR550V6Z1FyZ+4Z/LSfcbZPy3SRSP19IEiqYHePiz0oq1JDHYk7/KSesCLhFrTlaP9mB8g
vOhbkiMH463Vn/VB2nJ/2QeRUwSzjz1akDuTDXwKbcEYeqJp+xLRAYvFgd0cOnmYUd/nynOTJXr3
o9zRBcoTFtIbjYNrko8oMPkG4FnqqXBu+yYdf09vamznJC4272atTKNBIhSN27CHuGpg5ZYakwq1
ChGAStDnlElkI62TA2S8AigS88OLO9yQwhW9nGXIZ9qjgAuP0kNygfrLLuH8a9Y9NX6wG6ZVvzlo
Bjg12D3yKFa7L3aGEVBuS8oWBEx0q/K0BH+QKBkdotXLhy9jtwOFwF6rKeqHPbsarFL0Aw8gQG6V
E25scgOcDALaRLOWPjBjkeCa2DBO3aA0wKmBHWW3yqke7D0v00AGuSmaCcsnFbjHWehY48pBCGC9
ib165F91jU4eii4rg5JNsi3O0ZEmW07cHXQz9mxEAyjkLUS7C3JEJL7YWfbUGpt1XLKBJzU39M5Y
LffkkzeCpaGuvkccXkqiI8BdmeNsAfmzV1QN/hl8mzlwa8vTAu0lOSHWx6wLW+SieeygEpYlyVR7
l6ja7VurPzDq20XA1FkC9UbkTn+alfeTGgGuoNSNbq3+cYT2CwFw1aWvqscfIiwp+49jq/fOPEjE
eQS7ChRofnUrPygm3/4jFulo3bVLIlrE4vCfujXyTzdFWNu8vHVBXjg6B1ymZGfd/ImySerQ69+V
jMxOm+/NxTvJkDsSuIVVEXAKj6GDi/ZNIFd/L5n3khNq3rkkO4D6f440z5H1s6UfsN/x2gLMqHhf
83dG9t5u1oQxlVVz+d/roRTZkBboqal8dF+TF/yS7NghoyN+KKml3+nctuzMQOszrY2ipY2mG7g0
NFwwWnAORbr6s/6AsOCzgjB0RcQcDHExS/yAuKL9q9RScUg72BMqxdUuNnmcuHjQnyNQeqTIWkof
+WsIWKXKpTi2zseoFKkv1+ld3n2CXssqncMEEMX44b+Oyd9MG9vLnTCGZzK3HccXIjB8VEgakLN+
WJywVgV6y7Nj1FIpsqr960N9HODOeZO70ZIiWUTWpOb01rulgzyJdU1PJnk79GNSyLizmTSYFR3b
kaUckn84bGv1tZGe5iMTwVHrG1Kp5b/n7bgXY9DlANn0Kj1fs43O2X6AkXRTNpodSN7uZCR5Xqsy
l8kbBGBj7A2Slna9KB8duhW/J2CIfi3GR7JFprQy1bCgHKx9tBoceEsdlsXaTQQUJYkZe3EM0DV9
ykrb8d23j/PG3GdVG4Uqd3ns5qE48e85In6W3juWHj8dPLGeyITYx0tnAzFEE882ZNq6LrYkGI/h
4pTWCKKiYFrrgG45UmLs4SfxCsYaVKC++hgAStMzKxSSBUAjjAP6TgidgYo6u8McGeewprN7Rqvr
1DlCrp0QTcvHK0cfZNESuUiawskhcQNqOZOjd1v3UoREN8bJOTzWywsxnNZoq48ULatqNSHnxSqr
Hzy8aKUTULXZT+tGTWscWljlxIacPDntkRf4HjhOQoUAUMgl/gsxEtWUAUF7979tNkmTgWtwm2oQ
WG+NfYSa9G65BSbxPB8wzmdThmO4tgPI78kX0OUviZHGSX37KLyzNSB40WUlFjjoASNDovAtb92U
3k4GN/hfPAgGlqf7cb5sV0AC3G91PBoRn3UhD4OY3VDhfS8vSPwz1YX4vxLVDN1CBnSz3+fHublZ
7VeYKCBAIVJnhpezqALu3w19j3NoKDxXNVjKprhDWXI/PuPZF6fQN35mPIitK2xT//JQxbV9OLMc
f/kbPM9roMqtBtCqBaaGEo42FvnYYAotUJn9wj5AVD4oip4F1LtyvdMTzoW7q2KiSwWFCaCzxIKs
OnfNDFb2KpwWdUTOTSzj4M4A9vcfRHHd82D/90iKWjMm0G94PPdcPvvoB/b1n8waclX/6OySs/Gs
8JoiQ/FUJlAR/RFWaLjPrVwuxf3hN7YJL3uAHcGjOTMbpShHZbZBnug86mV2MUK19oGn0DjmyylS
1DSrLJCsrDKYshctzpY/35Aq3dZR6UfIsHRYytwFG5No5KzwQKVJAoM+kaxU45kq7iUpgiKZziPq
sTEurv3Uk7DLXqcqwTpj251BfdkKxZjTVGwi+w3hN/1imcTO9CVaolwcyeL7avoJN7FVUsxh+FDD
uX+8V837HYZRnwYGjo4xBdFsgVB6nTgFJ2RgGSoR+YaE2mFfwPgbp2KDvq//5VqPRSdyCXZio9Ij
IthHF9YWRNJ3dZDykNVBfMkVfiE0Jw+2WVmhEPhu9HNouhtLPuRPAOuYgD+xnm82CGpGD5mqH5xg
Sbjf0F3Gf0afUMKonGJMWZWa69/5J7rTdSU0etrxbdYf+opvQFgVj8Y+KOGzawupHQYV1mxVAeS2
In+7O5zDcBC+XTk1d7Ozy5N3l/olLPCK0jSyNJA6v4wzZex6JmX0q3fKZAJ8GqX+G6pM2CSUjy+t
H4qNt+8BOCocZisb3vw+PRg7ZrPEk0P54Aaq93fy73I3cg9M/D9wbFtvGqCawHUvBEOhlatG1ZrC
FfvPpx3ZZ+sa6tzQcDThDITCqnuBr4RP5UNJ0aBGRIMY1ICPBOfCSUuF0DRNSO5wH4C99Yrv+1Mf
WocQXPAwIt4Ioevg45SqRP2Ay7YtVY0XhU+3W65rhsBoQCzzGguEfiHXxiPNVWxYxsFL662lJFd2
HK7vv0yvVsIvmayrLAdVANhNy5Xg98CiYmfnTSsNjfQYrFTXgNRz03PxEOAJ9Z9tExbpU7LSlbhk
U4tShd0saUvVecR3OQ+VJ3Cwh/tP6QJyE2Tc5NjATZXzgPJyYo3fdIy+av2XK59rd3xicqjpJ0aA
sjhOlRbLd1V4s99yPqMj3hlezEaC1BlUNFENPr/vxugM9lJek7U5cUhm2TiTDGg7PbmJYkFWZqgu
QITvaOBdWkBYy7/g1WwrKgWauVQrDhgXJVTEHgDNO1NU+OAAOCUDMKriESql8bwIxzZPtNIqXDIO
GGf1ULGKePS1CJO6HLXFC+g+uEdt+FD7PlOvt9JTacqIJ4iR4Mdhys5mD35VfPzdaJZpZi2UNHZI
GbSS8otVpWsV2v8wnYFD821O31D3tBhWqBH3NinNAbL4RY6vw/0orzrPGDA3oNsn64zhJJtd0nk3
ff6lB+XHpeP+ItrNQNWjQ+B5LtLpddWRbV6gcJnfeOjPLM0dkt0md+0HkKRWZsMZ6q28IYqwX16X
XjOF9IHfjCpy9e651LQY7OsGtLpOKkEPenxhhsBUDpuo8YCcD1GhjeWUnytLWO7tcIZ5fyTO/Gjm
kKdjbO8q7d+wxyg3crMLvrHyY6EtzZTijtqpwCd3/Las9h8P4XnWyZ2zapph6QHzrTs9PKlW4lC0
RQyoa81ZqSdMLG8ueolEcRUBBfQYZkZB5Xq0g48KXsARx0sxWeClZNJTz6prwUDERZwasy9i+oKP
5MF59/6/LqMmKIWwnpYoXWs79kLWMlqeb38+doazsGSyPNl7r97q3PoOwhKyx0ef3y/gYnk88IzU
i57tn7mxRaS+WUIStSAQmRrb1tgF6BZzT/kzeq1Xq4G6la9J2nXs0/p0GYNQw5UtjdU6ILHf9l1v
t8rolWRhMzpJVQimlbqgB7fsjjzKyNuW+byxPeh3Y22be4mRTjGkCESOCoFf9vMXCrxL/aHBdCeT
zBz/jiPn0zpUAlK3j3o/ECumciI+rea89qxm4yg1sTg7NAif2lriJkJP0XGMgvO3iWRJpNsGVXUT
NuI4VWo0DpLKmcGSD6YrnoYeIjTzm37tbZgimXWO0xR4XayvPSnQC7AhiszWYTl3+LzaWrUkkJiH
ITbmJCPofkuKMSyCwEnAEc+fyzOXTZz+5C4SNJbEUCbEsoYi+8/HRsWaIF24lrUWf9T50tJIe7Ug
SzfRrM50nQo/ShrNG4i1VcD0GU3VKyJ1TmTM193x4+328od1M+ng1QnFQZEVDXzL75MSAIjasiyy
PXygWN29V1jihKoE/TweIPTXCOzStdF+C9izo58vWKggvr19FKlcBWAhr+BrRjMVeduI1lZQAelt
zV9+Rr2VJTf+i92itOY53TstIxEOERs4XUjGgRqTHfrqVpFCEk4cZz/JPDf/4cMv+a+PXjHfJIWM
2GpVuKoLCrAvi6HDqAnA7z8IZfbAkterBF/G9ghdmwAod0pOgup9yO3aXjRmzcdNqw3adpA3u4/A
+HFX4RhrmXD89ykjp3BUzauPeQRXm9148YnRmkTCKO8nPz7HGgLrqd0UoiE6g4IRT/gkNd1ZaIT2
FUi4TLNnoWUs8r7ElipUV38OIJY9/1KPqYu9U97tCL12Iazhd7ZNX1KIY03wZtH6rzktpjClMIdg
AwYm0VTmsSEmFMKBFx3kEJf05w+XO8bk+lNQgO5PY/MYuPyhc+hM4BkViVoAnx0kY5OlnPHGg3rS
E1Ym02ltUW6MtmPGA50Rw9b3xULi9QrLUV0d8RQ0SaOxv96tF/R5sr9o3jB5DRwwpAKNhBnuOMBE
jEPOjfkltF/8/eaNWlok0JEShVg/J4PFlhFTWECNEATdqhBLwM4N4eyd/TWs2i9z81bMYKhbKEsy
m9Oy70eS4tWpFqky0aNwVdWWt3u6NeNdGnJmcQzj0n2/MvL91cjKF6l9fMO/AnU7wmqMugit7lki
E+RRjMW7qMQIgAHxCFpYm4I6qZOo22Qg9+qL7FfFos5Icor4P3/PPoKdMhHCpYNNei+jP2ebQrYo
R+QNcsZ6h8TfZMKRz9clcCnRfM3IoFloQ1y+moQ7KB1Sv/C2OT0HqincZZxl4HlJCPsWKr/oJDqq
AKmPV5haczL/hab+sktwbT/yxeYQJd0skZ6i6XavJl7RXCCcS+x9e4FvgTX7dNSqc2JT6uW/6H3z
DY/VO3qH2A32N9DbhOR9YzW+pzcnFcQPdWQ3+ckTp92+GWbTsVp2iImI88LWCWm0BS7aBzKCXhPe
nCyvGlvyPNhlMnxrKYWk0f0sb8hi6yBqeDMTtSDL+OfnqOhjo/cLJfeQmGFobRBLLk80zMJgC8jX
WPL5ZaacVkn0zB2yuELdOjeW3cHD5pZlRwansPYL+mKv0d3eVKUrFk72E9FYJGLi3l2Ep0/WouNx
V5A8f79NqeFVmFTujTezS/QWpwQC03y0jCk1lSo53R0sOlphey5HRkdyhnxBDm5vCPk97pEAI9y9
Gk1FUNEeczfb7uULJ0zYP5GzIsmjnoucKZIvnwqxWqHmJykXhHpi9L4BCzT+WKdZDzKu2wyRNBDd
tTU4Q3VomLiWtmL1Erq0PUKgWYvbGXCnY23VEv2peyDcBNTchHvAE39rSP+Mm/K4wnVE87NwV+4r
LIYMqQweFFZZXHXP8OftoqJYvmy+5GatFcJHZo/m5LX1dmE0WQsOGhMy6AujfnLwb4u5qRGz3zFh
9EOt77cVBZoBcxGrSh9PCCdTnjaRPr2P59mUarAOC61955J5QaXR2rVT6GdZ+yAaGjQI4USlVJzn
JUfv8dQKKQy2gmrLF14ERrQ0X+rZghNaoXQKP6tFBz1wNABJtnyJEAPDd/MDmv1SGCQKIeZnovD1
rmV7SZ/yIZ4psCfX/45AApRrzVqzp+FxaUeQBHS+mr7jKyT6ldfRL0QyGfSUK1vrgdqAArSCb7xN
6n4soNwz87FAAr7HbrMMyc7lyJxaLw9UASq18IDG600GfvptIMPLBs/T3rfrNB4Ed4lokRBJcUeG
BME0WkwiuaCEat5QvvUcUThqqUVeAF5zkNzMitvlHVa+FfhqN1kTucrkFxucoOyddIURqFSob8Xr
WQkC/e3jBbPXFQz03KGNGuA8VDPmNE7WTOEhG0YCSuc1W1kXSoAC+moJnKXwBZBxiFzz/1wg0fs0
FtF6AJlCuyinvzWZsni8WDS64k0zjZyRFllzW+gmL0IK73FPw5SQVi9O0WbLh94pFvyzHtXjKwWg
vnsxlF0mndVpjcRzSuoNXxME+Uv3HqmrB6B6c2uqUxvoU5DyNF3UipKL4TJLExCzc4Q31er1azEE
QQlDIfAZ+juuR8xIvvk/R0h3sCpzrommJLxR4HDLoE07ClOlmbmifRa996uetQJcqkRwWIVUVPPZ
fAgsVNC0vps1Sw0Effgn5XRRbVSRfZ3uQSjlAAiYcGwC4KvMqbAHl+ZB394bHoc7vQtvtzBVMwYd
+gWflNuZW0uJmziczBYDKkY9XLadVoaM2FiFgX3iMDLaOjkeToed3Mtp7gut/rJU5DAg9JU+emYX
x0CLGnTxAvhoyIL87MOtj6f5Ro46DBuDusHwAoWa1PJ3zntlBWrc1RWQi4I4OKlX90ND8BP7GBAa
5ExH2BPlC3CsYMH2iCbV0e7lN8LTmbk18wFR9rgf0dAFLyuHNfNC7p7YF5mq12oQRm322BWBm0uF
8CR5KNe4qtcaucZ5TuwGeFmAcSFaQ5uDig7FVCdMJPpkbv2PEcTGTczC0rv8v3CJJqBDZ5BTugSk
quNv7Cbhb0Py3M3Nw5oOdAkrBxvIbUZE43Gt7BSpZ9VuPItTi+I4V5gcUQ1BMKHxWRxlbod2gVw/
WpffEyOQAUn8K3ciakCDxks4Rt/1/sOKuAJClhuXjpGmIRoBDWaco3Qpb4TThNf8gc0pryNBBelP
XjNrxn+1hQZ5IJD8axCSvpl5dBd63pKhvIojs8KmGO0vr4sddqUzpO0s3rI7QX/IirVdtico/waI
VbDDCFj29ddxbgW/zlaf6xhuANg32Pu6Dp02pTdGRh/TdC2jvV4Pyj13mAIHXiFDOkC3qwguQyGZ
AnPKuXUnsFOl4QuCv9DYuWT2PQZsedLtUvvB5Unzm4595Ky/Gfjbdd+JNzd677IEJoKkEdqQREUh
fW3FbLRUfP0Qtz5USD3Eog0mpJJ7xME2A7RSYWIeUeNXBfm4newILAY+W29tKLYbm0eFpXV5KLlA
Nu6SHRZLrKcmtpRXPrMg5rqky4cVZ91GosDsX2D2wA8K686lrXA47GzOw1Vj9V6Ak4dmeapsi5Q+
d3k0V3OqP0aUfh6FNCtG0Ei5J8m0lRZg0GBRmBssNhG52d0kv2XCtsUS07VwF8EQe7x1Q8saW3ls
eUOubv7xrW5GvYhPxu903X/Nx9l+K3zJmo1KmKKxdrhzIlrvTk3FNmqLRpzCNwMnbmvv5r0mH4zS
FAFx2ga/ouKmuxH9NbUAv1CEDQ+bAVT9s67e1gI6LBgmjp2Q42D8kBu6Llagv8w6oVbkl62jEdO9
aCW8gB1wP1pfqctFztQ1UhkZJbUHVbNcTDxeBb22KzveYlvfYgvauYPY3Ps6ElU+XZj5wu5rO7l+
N4kK7qniyrVscZy8KISodSscY4o/JW9N7h3Qrssjpj2fiYbkTTcuUF3cobgSGgegXmqpWI/t0wXT
JKH91ZQ2Gg96hsHjPJ2Lhk6/kVLWp+dRv3MAsy9peLW1S1fUXiqFY2ebHLpJTbLYvuHAWrg3/kei
fnbpjgfrCEdpBAFO1dtt1i0sJZ2xH+yWwWPtRaTYvd+RZ3AtX7rc1yok8bFF2SKVExSt8gGBtVLp
p30Rq58llDqzmNuNF/un7idymq6SRrJbNyUqZI+th3XpCBPEBD3qBXeT7SFPQ/ql4wa53sBEQyMd
0WBYTiSdq1TcAItvQGlAXLOoOi581VeVQPVSanN8/LXFN/ZIdEtV2yFa5Kwp8CS95U6O3SBJFXQp
J50vOdr820uHAYpWN6yG1CwJ1ErT/R+Rnc/KtExl9eq1eQ6T9+9Y39Ruv1pahJC5Txh4iCMwzp5L
HjRA41gXqUUH8sdaC3NZad+wmhCEj5aixrlnMgChgbpOPEtmw4wAAQUbeUPMkCywD/vP7+E3GN+x
JElxlzgum2USmo7viLNvpFEOiE6s6A79HkiezNloGRhw9RUr3nDbC0ZBxeD6E8gLEuyYT/kt7EAx
ntjwWNotzqzEwI0qs/4HEBUlEMqk0uon4+L0pZk9tTZOIcpEgl4BR21LpxD4XDYlIreMnUdEa9lD
DsT0cvtKYdH0SeWKUO+sGZgAf8ujb29CTq7XgirAW8BgrXb1Mx2iyhTpfJmryAPKDBSNWzutOC5J
W7LbNpNF9I3Wx7PdXFTHj63WcmvXHvms6zVXbPiNTVqvr20KDS2rOq7sq2lvIl/CGbP26uIoQHwJ
O612s+wskWVEcruJ+7nwBOIVmODevaIKg7GTPNYX8/GscGPlyta3+LcnVbxmDbis+ekO8RUB04ui
UfdtEr7UXC5UML6B5z3f5KlCKv05r6I6nCsBAM8aFiYnmrUcjrTk4pmtfRvXuvkkXabajvrxKdpb
zLIQhkrNgBrodBOJZlGHUGq4tr9ThQtsCEBiWtCR5BqIGL9tqCiBcoQYyka+dtknK3jPRwbpMq6L
ex+2AJiOGfO7jvyJcNFRrO5NGi0az+iL2DNK+wXTUlO/Jy2TDHUXpLfI9ZrJTvLwqFhvqSBT+OXB
sGvaNs244C3DYp3OUpGKMGazQdqJyRSEcnmYYaEj9efPBYa8OC/RXrCjEqk53j8+Q/5HfV/p0YKJ
FJBTNxPNlSqQUlb7YqR7E+cx2qd0IW0Kg6brA1A6TPYOYzKC75DInS+tpOBYBwOnZbJd4OwFqdqo
p9Lvn1Q8BEa06ugrmB/OCO0ZilUW6stGzKoTzC3gdOlfqa3nOPWF+xMn9O2bciE0xiARxr0LA61H
LMmeNBky4Ptt1wbaUNBACi5YC/tV7w8qxwyPGKU1zuHzywq7oXHORxM0n18tFk9MflkaecBsynDS
PeqqcHJeBRJeVt2eV+uq0cxZZ2zzIdhZx0/BZdB4WaJYeSk91JJ8jONOh+5lqvcgSOyGLM0ckIqF
KtZ2f6uNwbHAprEAXkgDgKY18Hi37CAZu3xRTSFtHu7lQaNX3KifhzzPar0KJJUe2f00o1XfeKcg
uSYBJ2lmfcNAG41AMIhrJy8WlIailCvaPZ3+oHTisBwRLHAl1aobt/8YJx6lEgUp6KwmwMU+KYgS
6HnVhWOTWJBOj7q3J5fyRuANo2a6LzouRFVYmfuGSQcdt48QnYK4Vy3tzRGlzGAoBCAL0djL1C6H
Ntmoov54KaJPcjvhnW618F+cYttVYD5AdB5cjtNgOxd+0F7qTQewrqLFaOQwgemZ+sdAWm2I+7Xt
tkL/lce2Ic1GZkWFHxbiyJdGhucCuP3b/i9dTVFkpA8xT2ExduqVMk6qEel1EV53/ZEYhgJ9oTjV
SbjC0JQEPIqkyEn0ET0IW2gmCv4ixFcsxhEOD7aybi9mguAv9+AzOZkkizuX+/95z+JPwM/rlMlH
CAneTLFnXrAl2SBE7bU83lmmR5s49RYHltQ/ayb+mX5E3XD9XjTuIuEZYSw/ccC+lpT92MdKhodf
F8xflOJjfW7dxRD+Mcej+kaSQdFYfb8g8BED0/v76ReXT/atdWEWBlGjYTBHRrpGdqeGFG2eFvhF
esx4RZVD5KL2yL53xgPcWXWna8+Bdm1w7pl/5XHrpLezw8CbfsJFR5zIGZIPQPT+928bqL2SDPpa
8UPbxZKRKoYfF4Rox/fgk+LFx/uLQ2V7JjeSwgRXBTwo9U8lCZLwNUlQyIpmz2PEYI4xUdhBJkeb
kctb9XNY6d5fojdOaZztfxT3u4Mpv8cGXMlIAjp/+4H/dHJlcQ0+n0ZAJzouTDkF0e4rjr9PCoe/
pISEYkL6VwstHM+VGogv6TrMvV1pUTNfUz8yJZ76rkGw+XRKIKTiCRBFLo64phVor/Mwk9HptO0y
Xz2qNUXCyU7yYTzQWbLjHTm0WhESIzu94mrwB9DPcDWX9WepGGqxety2znE9N1HPb8XPxZttr/oB
XZw7GDbveorHWJIbUDYqyrZplKwuXAimFTvdZpuorKG97M9p3ui6GcD3RBAy5QKq/DcYgvzf6lAZ
gE/MwEYt/jK8mxS/6pPi5pCDiWvRMS7yN6Ztzs2jDYZiyzy+K8THP0SA+2Pyxjys0fDOBDfjEdYJ
54RU+0h0EX38g6tsXm1M2B4xoHCc7bDYu8iJ2xjm43qwfnCYiGpDxpYunvwP/G4seyVq1wVy4C9a
0cHLbN2t7hMeaXQHTR6tktWE3jZhx1iQeeq1MBICvDdr0emTtTIBzbOlX60bUhtwg3w3CuDyobUL
XH28LNRqt+hpwkEMG94nXag7U1oFoZeEMDAv1URzvk+r937Mbm4LSZPwwaZtHPAT2w1uCPnqEVGx
x3em33XvAxItQvRyN/PajfbUHnAlE91MzQPHmnjUijBBGPhVXPMJjrDxK3wQAcjYqVhomTvH9xBU
NZGHJ5lqw1QYVQOprNbQjPmgZHc6xdMOlFCNDq1Gy+R/JWgX5u9gMTx9Qe/BKK1xTWCh75xFEcy9
2MP++WIa6Ae/fPeBMeZYkS3U4zFTDpjalTKkaa7GVTIAr3rsvTcduiTnxX2iNmh9HeqBJ0OGZvnm
XoyCjsLDaQr6LKZg9DJ+g8yVDCGHmDIQSelB7hmvDKgL7Elj03d8fABmrQyMFe0tL08cjTt26LK5
5STJ77ue2gu+McePn6EhzyHk33cocCj4wtuSx0rg0O/KEmmVS4lUzUgTo9HI7dooPdmra1bmrEzf
o4xQ8qp2rDFOE36lJIH73YO9SPnighs5O2FL1dGEbAYrEpiv+1AgdzfbMdeUPbbwH65wOldJnifC
Fj3L8B81L1SXntXT0qz/qLVoKIKdNulR2j7YpojLhH+db34Zy22JiUaW36eH49n1+CKO5FxSH9rD
+59DZm3bjsqckqQ5ep5fEiuq5K5gpU6Z1/VTXjzlSK20hmknhSYndwLN9s5N6cmykGX45NzyAIV5
/EFuoyL8o7jcf8p43UO6C2PXiRgpzey6PSfoZ/Xr0YCEIwwyAF09Y0DOE22B4OKQo203XCgM1JWx
WmJkPAhsuij/kO4+/P+pAOfd/9bZnZeqcOjHOef3bcYGkanzVG13CYiWMmau3/A1XX5r6RclXHe8
pmjK8bWAWzxiEyA/tvrsXgqab3ebirhlpbtDXUQz/v+eIbz89Z4Jyg+j5rmqJNaD0m05B4BnM4D/
K3j4oTwAmYB5y8aK7qYUhL3O2y61NBN5z24daIoSOredBnteKSD+8hbTw9awMpT7MDqtrk6hltxz
RNBnhVhsT6PTR1sSU1aR0SnwPCyGqsyRnPvkydBSSi9TWrYk85t9GznmjY+XlAJ+YZuHwcTfCMp+
+Lo4CiKNrkF9L9Qt8iVDk5BjkzX9RXzsVtCUi+JXM43RvvP25tI6EmiC9pHOr5pbZ5tIo8kUOg14
/YiNSDBK+RMCGPWbZs+QK4WNJUp+PXvT8r7tY3URIVknYUxS6x68+I4l5OnDTozSKDzrgwK4SOBW
bCjC3SnCRNcmtnfAjIMJEJHppPhwhn584qPg+K99FKJubcplERe+j4RzE6fP7HT15GXnflVEnaLh
BrimIDvmFspbpj9DA1c4g2tbugCjvi4JBnm7Qc9mWrbo2bHCGg9MLXDvNgkO9kYttCpfufYopzEQ
NnTq4kFeUa3/jzqtFgugvEeq+ST1ZSo3lffW+M4Ic4R7USxdK0cGgGnegXIUR2XxVHqzuj6gqldb
qskCrTB8XjQUsx3tGHdyYbDHA/3qxS0KNvmvW7P1cKLXVktb+Gvrmo+kaAIoAUNKtYMq6j5PFOxj
Twk6eetwrtisH3l0lZvKdrTEP9LpcEUfqKvkHJ7SB3y91t/XUbKQJypY+UWs42pvycisexMAO1Xy
3GPdE7yWr0bpheO25njCEx+A4iTABSo11Y/JRI0aU5HdYl4LMA45g1rbtl7f2OXf6utMCU2p7yxE
KJFfmOi/dwifLYqrK0J9PZsobzBo0GslALDKYXYrRpxPnnBXbQzaL3Aivwv6s6EPDX+yRftanJUS
YtHkMQz3KloWmaL/Jhn+RF3zb0NtogWcGX73oHSeGyysbRlq36heV+hCQSSU9p6kZ/nbkCMQHEbX
alR5yiSzOfI5adFrTm6Oddqfr7o5lB3seBI1d8LWfODK/iTcD1wjIQZCiJSiOL8S2rqaMHUlZYXP
FRzTuMt9YjgsIgzNzNHkYdmlZmszF6DdhYsMKOJ+RQzhAqIJM/ORlkmUkrD7QhzS6C+dYeooURfj
wEL1opxwTQkXbef6E+1Vro1haDneLStcqQ7V/qcN4/B2LloD2yfZjyJjozlB2t4efl+1nsBGsbcn
RvgCaRbfIl940JqhZy7l6t3AK+9wdM8+tCl5GSvX8TCICEdSbLjIdBH+z5Uo6g51Lg470dCa2PtB
2SKJYUXAxmcuKxgtcdu07VU2xHJAmo/hKdjGujs35D4HNITTwhuOOUOE9mSqDZGTP0ga245u6Go0
HYLw87MxgmrrD2ypUk0p/bFvXbZ+cDuhqdKXucthOniYbGN8xDnqevuo/enDjsE8rgrIvx5teMLk
TSYjbWwBGQpvhGHW49YjpZ6s5iXca3uevVwF0pIO3bQQy6rQkeanKVxD5mYHwoisJg9bZr3oCiS1
T5O3ILEYVYmWuV0Jy5z0w+GDwlxZAxkOuL5v8lDsj/Z55U3ShGu8FtoIMftcfDkZTV7fZzLmpESW
CFWTLVxustg9WdOdBEfZ1/mjJ14Rhr1TR30Chvrj4xjvKPrTnaVFsQu8t3KzcpGDrMpVHt1s/qO+
nBTxBOPWKM3x2LE669EtmFt9MXmg4eCavr90EIb6dxikbG3smXVjuELRvB/crVwbcr7LlmT5wlze
Yamnav5wcnphKvuakrHqD8EUCxDTmKT/+8vOrSzHCWIWN2O03MI0hRnKTbXdMhC7Hw4hHQ3DEg+Q
zeGjpkWqfJr45jq7BFPVLyPSxiTbpO6EtBZBlK7ERZtues23IBnl+aie2JjdSUI3PVlWSjEDXAiv
6OYB99d57NiUuTLlRz5eyQ30mHNuGaIM1wKD5v46pLtUiQ3yIQgqrHXFK+nRE9j81PYk3kng4IqC
CcjzNssBnhMByzUvWLlZQDLuSWT25vpSzzd6+rXC2/4cAMT2ZrsImqS7Z4sB3LuZvf1lfnKYl8Mg
DnQwau/E6Tgh+pfosCfZkXiBlAHnNxPQ/HtxT9W1Wwetui3BTt9ytW8dTQJaIF9mM568POc05632
6nqmxY+4GugwcVrV4BJazbDMuuIQsVTYEGIguzb37Y4R/fAEWFVujnYMZMG8VyFXAZxCJyB82lst
8GMXSYWE0KRDuXuMcxRsk/dktTS1hqJXQcq5jjHG/g7ALyjGlZ3JILQPCdyQPI3gcE43WXVyQH+y
DrHuvczd74LxDNKxS4D+drmbkwwU1HxVeuaPFCS/kI0f1kcOz7hqxSWqhFlTZm94wne3TAvBjZPV
MlI3w5HjQxzk9+aRMIw5W00nvtITuhGN0k7xnbfVGLBeVdnYgN05/Fu3GCO0igMJ74V/O1ZvphgN
06G9/3Rm3G5HWazHEOgn8JlpHWF5ljalKd8ytU/hgsixpZ6HatB+/OFB0g7TIHNEWjyzDmoTgIk0
85NTQzV5HwyYiBzuL1Y4NDfuIUJr7kbworaFH39AgHz79B/u9TLHuHNYpL1j4wuMF7qSa3+WOclH
GT//i7oUc75AUgvBiTgAYF4a1DsbydGl6raBFUDAWECqTzGVB0O4ves+iZcN33fWaA5dvkHnLz0T
448AbWhr7wobo9huEaLh41H6JRWbS97BKF7zVH73aD9Nj2uuQIoexP2u8o8VPJs2MyItRNJtLECL
WdPggDm/KfWbhzEPfaLGVqpuDk8jOzpFGDbXCQPvlmOIan/CaEgSI+VFukdcyfBdTIcmtMpecIJn
JPtZ3TNQJAu1NvaBxW5awsJZc16y2hYv5KWBpdfniaJTtPyCIo/Gz8KqHvw8TeQ+2lal3kdAJsPO
rN0wtFqwGS9rgP1Z/RoF8kgCSih11aHzxzIk2mG/Gl7oNeD6qcl72ZuJuSMAHh+MV0H4zF/nivZ9
AGixsDbtM8seDGteozfaCBVOuZCd3UbqNsLU0Rai5Q/QGLXJFcyeIMaAQoQ224h0DCaZBPQVzBWo
zqG9RtDo3UHQTltzMcOfQanQqsaTNr+zJFPkn8qJqMvZjgM321g2dJ+oQBzMI0Nj0RW9c8knkFnx
WHd5Qpf1aZPyLwcg+sTxr5GZlNFGyNd/YVSmG3kCMTCUnhkYql/uvd6lh7+HAp4rNgSxNDgz5gte
ylzKfBG7e36x3wf4uWL0aCqCLqVZKywZ+OmWxr6izUmperw2fMDBStgaTL5afVcy3idjje9ntWCp
hsyEupXZfBtbjuaMrhrRqfv4wxlxJnLk5wURzY6PhkSJCx4qmMOYU4h4Kci4RawAy4+07HFNe9Za
ae4ovDkPPKCmcSqU7BxL9Uo9qv2U/AFuiStcGBsMQqxL86qrPTqeNnNZe0vptsaLX1L864GVINY/
i0BORxuvCJfyVb9Z96iLQSCrPZrssF05IGbaM124B5HWw3IptsSllVlAnDeFbfx0FQvc1gCyYSWR
vKWTM3lX7cu+e4xOa7f5oChM1PybC8yHHNHmHnQ87vzIK3NoAsZKCRdyiUiNFUNLgs4XL9kxwYPG
GhU8QS0n9+cUkhFfXaK2DWP9OeFKmZe/RjUssq9JBGCuQXkAuDmuD32sxHj7C8WgXrjkaeTiGQNM
7ReMnfMpb+4BlJ29fFJYDK4gEIZJkbzFXZ7s/3okr+lt5rNtYbLfHHlWvvO9C1x7LTi7XOOGwBpU
O7AxyZ7gz33pfTvR+YEDVP57ipJjYCqmBuxRic2Jq1DcEbXzkrwVWQzsBmVQUq9bvcBu7hVNNz9v
fA+GbVFaGNzb21ynhRLVIdwesfLc1EelEj/iVDiqxuy0T5vgyVMlIpGXi6P69IlOU/jXasDzhjNj
cJbjEqx1Znkrwz1nI7er6t1cc2cUGMsFBB0ADUf0wJIH5P7e32SurVjYkL7t7YA5JvtDRF7UHKWW
aj1iOfckFKmuAFQtyoQal+amH3XKOXsv+SXPBdM6jo7TOKiqscjNvoHFuDp7GPI2xH8XVcY8u999
1Na0Y2/AvjOsijy/bOni86rH5d2VCybL7/aU4wba8yY29S5+ekm/AzyJqXZhR2F9MtEtoD6GNu2h
PaKmL9rDJU+lnQ1Ft/gu7Ijoy9J4Fe5FU1R1wm5KFOK/zvUgcMgZsCAtj3LCUmAyRBtnwiq7PAGD
QP0khGBMBnuIdpulpqV54uvbLjYAF27/Fyi+uDg6d1fupGQqJaCkZ4ohZWSsOxjiAH8Z484G9QvC
XEFEkEJXJ4yIUrG7Hr3XQ6QL7MUN27UmUDybL8yyPdNmsZDKWW//AETIWQ3ivzF4j9ON+BVaes/P
G5aEPEgEfLOX3aVFlWa5xxNxMtHygd4m5dG/YNJDGq/CKDhabwiWO6vlc1lUQoG8GRbojzezcVtd
AqdjWCqvsbGHpGA/CiXk+3GmWOIijCyvQV78rQ9FWE15TlTXSPngP8MKXdEFZgpFSNyzDQpZyJgz
1FMDcw5q0hK9udlh2CeumzDum8U97QeSzj7q8SRJ1wPVFX88LCsKQwft3pbjnBzU8eZkP+DkpmW8
0w6cf43Mhm01fBIkvRiZ129YgqB4NdxL6xZJvBXk+VuIMI9rPLIhwpTD2eLUa3EKlbtsLTpPXhWC
jxoqgQyXJyDa3UKHCFOBthVljFMQ2xNQc4UsFi+mOhRlmMmpdW95BiTLNaASzs6zgcgI+6pNjNlC
jxkleil7gOPgQLvzB7hTfFB/kotOCF2cmu/TEtt0VGkSIhc0cKfkKZirbP8VD/b+XNdSp2kJgk/H
oOJjuWjQ/RKUqVOoyi1B2JC5JqRrUUH6jTa03a2lN5rY/8R4MoIC9qd7jJwPA7rLvQIurCMGh/FM
Xp3O5sj2BXrDPy8xh0I3D/TRazyOOb27+jHMKdU6WWpGRiR1trWUKjtODaPLqAf3l0KqTE0x/ITL
kvR2BUiEj8ETHifyNBNfX4AN2w6a09uXqjnluKCGVMFRPE9PKhocCcEV5rs8eog4ohUecmg/XL+p
4r+ZMnHQ0HRc4frY1AzQKhxtRymDHp2xu9jn8/oVrOFZ81pPhJedii+i87RXdRap2ag8Ixhxf3qk
7rVEUpVp++XR3/pP7l1mfishq79NPTkN7bUKNvyzBW4t5V/ikUsw247N9NKiu2kiCsevJ2zWYzSI
k72zPhznsUmNQZWhuxn8qXw+/fm19qK4Jb6kTQ8VmzCMd0LDC9LECqBZwL1jYUk67PmDdmYW2PI5
cNVrfF1taHt6cw/2VdYEOw5w9sOOz6ljkl3ftwup8t4hFpkPtqsacBZFyTyc8axdDUhDjoqJg8Y0
/bU/VIo2GgS9gw4reHCS/lawBr3twC+fqt7ItPevuQEB7Y509zPxI//KnwCTsMIishrMzJtzs6OL
sqH/PVkWGUvePMjeM0HFnf+tBcLI9mCq96v0QPAUeCKrxf3BeQvNS+EN6JRZhSqEN8SSnnYzhCa6
m5A7QKpPU6o5Hrz/GYFYhLghZ5NBZ/i5jMuqW7gTtUOK/WOSaimC2dRi/WPvgsBwo5jorJO7s74C
zLifSTH/0ExjIRI9PtCs5Z/BGml4JPYpOwyt7SqZ5CT7vkmfNcI5rZRpJU7KUkIFzl30GEXrHz3/
+caCdxu9ImuUImdoAOxwwQlYPHOmDz3DKpDoKJpOQoG73VittxNnQPW+R5SHqHBIN1nKrSF3/QVU
oQ5mqomQ5LhuONlpMFaqbjfXOSmN+DjYiSR4oLrNVmpnuXYPhqu2bm039In1vN4e1nSTNtiWkA5W
SmPeSBEAMICTncxBsULPWHSmdTAx7SmGouhfqQmPInEB/mDZ2BDu2lVg8eFup59ZbdH7tbeNaM6l
3GMuE2mKF/JcVrnvCtfytwTtlzuFdDN+vwHYmnIk+RqnGzAboeluhcn9y22Ck+9dq0j8/72tjew4
33wh3y0Cw79EHFGKWVggioCbjH9uT6u+cGDyurrnsn77Uh69eeoFE959+vxVobVqG2DugHRPdoC/
cxig2QZeywV2k10eUze0q3/mtajzP7cGcR+BJKKsuVM8cUBkTk9UkXqu2UMikNrH9vF1TqiGqGYz
DfRwN4YAa8vBZItqDyUhBxdbC0A0yer858BknELpev3msRQ5r27WrKl3cgx5f/IPgrtcbvc6Bzri
yNiF07jGRosifwEgzooAbwc3knu4r/u2nwbsrbWADWznGa3HMVRWgXxXw4W6zDUivJMzqs3pu0KW
yBCa3NbOBeZfC6uhARAnx9DnvwdzAZV3xUwSisDz1GRauucYl4yY2h4nPrSb5xVJw74204l0Cwhw
Nerp7yO8KpCCPQGM+ozoVifqkVNcMx4b0/QeTvf+Q/62VeXv18z4RoMJGqvxGpR63gSgyXCf+CGP
QUjK5sahAmXmb7bCm4WnXUOzTmBFjc2pb1SL5w2ppBOA8IeLO2xBaN4MkBzUCL5GoNgvE8z4mU0a
Z+HbGHebiGW3+8pIeHL5uM5Gy1UT1dqeAf0Cs9cPon+mGgxx6oV+F1LtnSWqO+fcTv5FMPMWkLEC
5c9sX7Gg2C/SuMzq4oI370zehj0ojbq/jPWcnBEXMrivvmT2EOH5fIFhJD2A7QlpNSBLBqqjq8ea
Xx38lWdfsSHpmayHxiHnIUEYiOkG7UHZabz63lgauB7IA7y5Ut1317YvSsw2R+l+kO+eSRVguNBa
iGtle28nxStTDwWih7hfE6aX2a6kxZWYLssdRFYpy8YH3bc1ZNukehM0L7Bq7laWpAfqbXNttuse
hUEcq2tMouIQfm7Q43t24hh7kR/w6E9nbaOvuOH4WCwwYdDCh8+i7BkSmTULYgr1RjTbcoP9BMiF
KvScZGXzVkrOr9bQ+vugl+ijajOOKdIytzhocY7QpAyVYCmCjUUpnU7DdpTsya6o3C5QobUYJ3pY
28eYrkH6h/YApAvA5MT4q5ebj/whx5GmoajhJcZyxlKPfUixezKvbtmKC0un94Y57RPgGnMwUOX1
vMGYSxFMuvM83InH44uGgepxaMi3O6RiSzV/Q0UQcv5ueH+6+YSXUh0XMMYmPbmAC1hEnyDmnsp+
pLzfZBEh5fd67j3q0e0lYP5AeLwnOYPSC6sB2C8+Lc38CxL1kFSD7DsKYxFM5450hhpQ6a7fNO/P
vlrKsZkoYQosys8aUYCMRONq2y6vkSiQ53Kiqn5O3UbqDI+mvibvtHSZKx42zxx6aIJFCDCCTI5u
GOw6fi4IlzlIhotrT4R9DQCzgnKq0+fR6HNJDiQ5E06xH0WmfUFIhg/t0LAf5/Bjasmu8XCOOlhD
Uv9xIrnIVU+ctb1phEh0h3eJblQkJ/3sQXwMuB5F0K0iLjiRXIwAcoAtYOZ8giABsy2ASm/gDkU4
HGROnUAJSLM85U4PcWQXBYNl8T5aO0dlfZW5GZKuYydgqzBoqfKulQjJVJdus8Bn8kfl2k7JnXed
tHFcuh781DGRotUs/9y+KJm0WuJofr8ey89xPX2wpXDJ+EzUGC3INKQOOyGs/fB+CHiviT5k57vE
wDOcplqg7zhYlSXCRKh1lCoBhQMENjZ6y7hgC4CH/4XqV60P2LTq3+XczENci0T3dp2W03yl4ICJ
ND96qxOXi9DBAJsK96LkW8RIP3PjIVQGfaeQefebgthnxJCm9Z+v4cQyHdUDuyajd1vvZm0s/nV5
/QTv/2PJgcRu8Yup95LGr2Oi0FH6atQZLihocoo1BUJjY/LHOf+ITQaCM5BvXgVl7+nwOlP9EOby
obNC1Y3YPOG2RWZ1kulr5phyk2jsSunBDBYXgwiyS8fUutHzey2GW3q7S1s5un3nh6thWXL9MUUA
mZglspGQBMXOhr2Gu61hhE5ukuysoSM112PBSmDxglYaR6WCsXCygoTSWBaZCQBUHiFczEcGApna
UErtzpf2ypWUXA9oiWjaWh1AS8m1zQBQYCBT5eTYcGGASP2N1DdwWaSB8J3R/0YypaCv2gsYZ3Mx
qDOYRlf2SrxMJ15mFtq3Zd37tkl/u7yzYsKAWIodHVd9FxZVnrr70UDl5KGk5rYYdMu7QIZeT0UR
tp1ztl8FfOMUfA6h8bDnaacqoFhqj+1aGGoxLzasufbeFItbbet2YBzVIIyhXo9GPpIxrGCsHpTD
fXTnE8+pwB4G+a+X0l+uH6L9MZiHDw5nR5qLMWcwwdtTxGTyTjKaucA5uLgB2KGUQmUpeNDwAThb
LqJK7TfVUSYgWc3A/E1r0nyMWlbs9H2GGeChiEZf7X/rTMH746QvF+a0BFoNUxYDUG+iBq49xupw
lxdwutYAZdzYVYBFzBGsKVLMuru3AVIrclaoHJni/b3jf8AoXNo4rfD6dl07nybSvDl9orKmjbfg
pIp52/q/EAVGZ4Mx0So+AXcj/QATMFM9bAIV8d2s9hZYTrlpxmheQ8pCjSZTkeL7a02sMSmJsaDH
BxUSp6uPVyfpfJR3dPD8zVjL/nHoJ8ZVtux6QsoeVOFLRg3JS2lMCqJ/7zYf9U78pvgu3ElClFP4
IK7jofkt6MnytMv4Y9TIICCDQO5/Tjlyk5hSa1dNSrWRhNXfXgkhklmboQeRmw1mNRrJEdmoOAr9
nDfhiHPZa3TxH0cnvkkzfh5gH8Y5u1VmTGYjb15Wcgnk25oRPh3ovlLjtEKeK/7O08A6SGgUOsxg
eJzJNvjqaWZG9GKazUNHUcXYbnieWYAJ/lw1IMV33CC51IZor/N+E7Sj05/QDNkWmpqp8wrnvwq5
diCnGDj5ZctT5UTrqXAn+6zY0oMJdoMTLP2KFyEpBBPACre/AsaQokfcBMU9Lgfl0wT7Vy8hrR5U
JdiCZ7GlC2YGJtCqdnyfftpLGpYJbxXEw1zvGCsP9e/7VS6mea3204RXzozR9VM9paE1Anwiw09M
wa26fNBBKaoP7Vls+wnhx4t/7E97n7qdfeWHrr0uIz65vvurKjeH0AoQv3cfRPFlVL/l9wXFyzB+
FWme9Z4qb0xzmnNonTt3amB12WJlR6QoYDDSNIsMcuxkU4/w6jVz+nwZldhx1DX/gnG8be8MLesy
ew5+oxQgvgj3LkeBE8jlmOe8okVLA2WmQjdzVUNVApig4gqu50AdHs2fyDfVkXPbQFeEPPo1HFfY
L8hMEfzxFDK6dE3ROairpH7aAm6W0uRNC4vDwWJ5op4fese+Em6V/tEqp0KB3cqsJ8hxA3QClkKi
ubpt50679/5FeHvyMbNl5pDuHtJJqE7qbkYR78dnD8qVwcShXcPp+GK1CDdpJG8KsssJBx/lmUo6
P7HH1DtCXfgI+bvngYcKe5QUqxBW/QsBfEhmgY2s53jH3izN58dpUia+8E+jOBGo0E31hT5MROC2
x9fGjo3UPdR8yDZ5GSDMxQHpwqAcDlY8e6dptzlGjDQM2CBQVEvgY55xty2h4KtEIlx7IFnPjRQw
LAQxuHqyk2FYsRS5sVedD6Fgfx5KgiqVMoPO1Nq/KhVGQ6Ay27CuTPOoyDA9thzvWYPE9zZ0JYGQ
lmAr9/jBBDSNShwjQiiptM0K95ztoth7YU+9Lns1sgHGJKpufWD3wLXjrwXncCkIrcf/3wUjtuku
4fDutkdtVRQNADvw4KBhwuYgcnSNcMJBBtW1IwPUrh7840o6m9iYbs3jeWX0qjDHMmBG/J5bjB0A
CHt7jb8gBdl4ilVauk0nrCDDSGVFY70Hq1P4/O9CADSaLX66mbLFj1/6K3XqwV6pA1lhErzfbGyY
uEdA98AiLee/0cilXWCEJPWh2dNmkxZai9M7IbHif6dmXGniolp9koCVf7x9tEtAiNgVFJSKNOwI
KvPHND2TuRef2ozwExqQn2emv/5KYX6G5dx8tSrYyFazFK0gVB6tnTEwo2cl7at8lFqC7tLf5qcD
lbrF35DDI8dbfUjgI0HPbUkuTiHHZxN7B4cDLhKR6nlTVYPCvwwAKs7NX7d3/H5K9HqoWjGK0ZJI
NUSQFm7H7aXKrA7C8RHjyf7WG1A7Yd07M07rRm7ZKWUKRYz5KxYnjrk2sXDABD8jQY0tM9fW0I1Q
PaQKMNOxC6bG16TIgaXbLUwq4i9oxlN4LXfsZ/ZDQe1jbCCfqEhKa00EsOfNcoagZOuAgIbIryMn
81iqdhaKIGBjSgLXWqzc28UoA1cTgxtFn73b2OD2d9gWvIDgYIiTAQyJ1b3se1aakTnrRyeavi9+
2fPqeQnSaLC6eaQxXTFwofqAv4masiVRuEdPa3Eecp4LrkfXCb9Xf3djAe9su+S7XTAGAYzAlM0j
N7kC6s2ynGzeUKAvYG4agTsACok2R8SSvcJpxeIMEA+v41UW1aPUOpCU0lUpuyDDAM/BB7f6qblu
pm0J4pS7DD6VMPt1DXyPxF5w+sa+K/CxoIgVlzZndKGs7U2ZPZ/Bg602IIhGNyMbM8tqLkbCzkkz
gDIruLd2Szo1FZ2TCUM6SFJVN8KAUeBh/QNn33QHpMfCTsARTrr+uemo1PFBSQa83zI+Y9q9FunQ
Oe314kb8kA/4L5GUPhG3OD/pA+elTH/MNdaHqCsWPhabXPGuSEOaW3Rqdvc0oig6YpK8JkeXvOMO
vo/eYa/a/ISGqrcFhpoTXl8xDHRCBkx9eQ3dhfE4rY8cE4fJrkkny/fojppR9cMc1y3e7wkmlfh1
0Tb2fjnuu9VqJOlVKz+nOZF2a3nS/gKnNyIQLuxogY8zAQZWwnsg4asywY0ldaSwGOVYs0SqWthu
lGyq/V48ucsKGHrXKZL7yGyvIUGh4CjRnrCHkwqZexDfz5AwS56XGa51cC9vTUy9MEJKTIvUd9QC
LwyUyLrim6W8dBKLDzNEu+iwmD04MmDyfHto9soCtS1k5uUWigwD4cxM8UXpzsSNXy+EWpB1RcWk
GFOxLlJxoyzR+yC1fmF0dvyOZySbCYg4LSvHSY9+MwScDGNwB84VVj1w6nKhIZ7DU/DIrxapV0vs
iqGJ5bzUs0txzBVveelGbUjdR7Wufi9/HTEOTnD5+SI9r+Opj8nlce8bRT5vO/joqEywTwthWBPJ
w5x3dDh4ZHbWUxkIk+VfdhDpfEFt9aYutem1VoDM7quEHUdia0YMEHa+pl1X8kccRYAjM56LutCx
ksOPJv+Euq/LME51OloBLSyqkvtOI3bKM4f89ooZ++Sjb5sm3v5LCp2Ayr7Pjvxx0Lx/LrklS85a
XfTQzFycWqWWkA8hftW0D1v5TjN/5i1cVHbP7fi5RHn5nrevgHqjrdTt1dk2VZ7Jdj0VvgQG5kVT
wP8A1zoqIXq+ollAXxnL15gcwucDRIAYIcj/fLzkfbWodmwbNWo6hJhrp4VWAhx2CBm8Pby86rTJ
vMp9VTqyjsDTvyHLV5NQycIGeQD82WcErAiqw/gWlfa0GAAGJj9x5FCU6SpXSZIZrQ334PVB0Zuy
q/qW+xSHrq3cHQ84RTb0DelMDfItt0+K7p4FJ+EP+jIQYdGpf1qfbjYUa0zHXOat+6fNj3oaWXlU
P21XYIf09MsFJ0YQ+LNQ83x/DguYTntVywJFjs7vE2TTe32nlb3txrdVNhUcEe/dXK0hBSA4Dyxc
I4QGtKn20uJMUZcufcGS/u1b7RJPRkqVfp5Ix8tK3gU6q0tYXu2IUYq1IXFWz8HjdBqIfWhXxxKC
l7T5PEHvfAcbu2k9JUb80ZdYeD65HXHD26eZX6MCbUWzIHY4Z3gcCvNqqJeiqchDcplJSLi3fqXO
CxqrbFokqBxoGWlsrzTL7kvP7MKXHJsuwIwfVdHy+ugsLnMePNdjjbCNyRUV9Itb/NmrTgjuF0gP
IIWn+l7EG7uDElhtWGT49Dm4vmLhB03UyNDrP2Tcw4UPz80NYOxsQmMDKrssjs3tLcjCnG/f1B8+
PehGY+jzh1PTDuBjDweNz1Nd0yp5tzMC8C1oORx1fHO0QmymOCtJAHmFOWsVSZc0cwIkjqrHw0UO
lAMC2w402K/lEDBDhaexd7NQcGKTediYkEnobLcUGg7C6bC07s0Ugb8MksJ4EaSGUHkjmwGsSJ+D
kppQuqv1q6AUpcF1l0MNnL1hnB6nM2iBtyVkx7iPVFRp3NTohlox2I17qkAJE8r2oK4cm65mY79j
giLYgW3Lclpw4bFCkgkQ8rzZ1dZNVGz94jFO5Jo245OZNlI/3y2Y7SfYhxQp/bx8e0WHBseJv9iv
yRiTIFkOa4iByh66WyA+kcxlj0Ug7iU4NxSJKuus/Px+WSNVpVrz1EaVL2zIN1Rc195rIKw8sJso
SWHcAnjmLz+lvW/Wz+0zeDcpEvZbRSoIE1QwpXvJ83AzkTj3G0ylRkV8FbjgpJl4upddHykdF++s
9LNyPRPAwrTRkiHa+um4KikJHAfmXyhsPj0SVNW7qn13c5eSXa+H+hSBrKi3F7xuUBKHOasM3CUw
rDqg1+/T4yVR2LKAxcgv2Q2UA+jKnjpdv3w4H3E7GdUv03uflOeuIr5gPvwYsl7y+x6u4N2Xxoam
itStZQd4hZAzBAsz/jcEl8Uhrv6qwqDMAZcLR+MICXru5xxWud941H+f2ZCKHAwrhYxhV36cH2J+
R1CTMB1Yo2dSwt665+SQeGZO9WE8+I4T6nv+QzEvOe+HfPlCLENt1YK+WZtNQ8+HLlwh030nxzjV
T76hNkRYZPS5uV8GDk5BwvalguIZWE46JUnk0pwkWGKQlUzDlw99WKnS1dmL1/zz2yZwJPH6NqlJ
mg70Pyv1pqIh0QvuwStnC6oZ5pTP1MmoRJMci7n3520jVJI/VIdDZsQwH2wJruFfCA+SAEzZZPpT
v0w1bVAIbl35JEY28OgNvqKGGQ6a/zDDFKh9hWYNusv/EKFqZbl54bl3RTCgr8YlMTOYaDaQoOmN
V3W0/AlHXgEAaKm7rglPUo3ueR+cTIu29tY2GKDdUa2t/M3WK1nTS3Pa+peIg+NrDRTGWD5K8FBi
NBdcy8KU/rqDZRMrwVY9rV1Cz1e/aEV/a8lmnXUgwZTm2f2KgTh5EKPCyLq6P94yLvA2MM+pSNWf
5hrqfkY3DUdcQAeg7Bnn2H9qZX5z/gVrEQITz178VgZtA24YAGvDM5NYYIGJtqRgC9poHg7g+T7d
ZVMZwJ8ak3zL0hhj69MgJsTlDOVBa3Kn8MQ/WAbtn6rS/rgfZh/Lf0tHQTLDOBaPNYo5bF4MCN1R
YG5RzQ+xcpqCVoDokmNXrFHDAKnWdex6P2z6nBTmv8cNkp+IgSIqgG6oeF3gVfrqS/c7EgFRAmQN
7xLfQyddz8LK8jW1t8qur6ojBpx4tlgIX3tb6O214frrS5Txnil4uNBxuanr/k033//o/xE0JCHi
PGgeocoJ1wJDf0z+BuWpCtCEtx5v8qoQcorB+yMCEOaZvY7TLIJ0fymSSJl7CfR7YPiM44Wz1ye7
D0mVt2mufBcJSblVaGVlNMR5BySNnuDNQJmEyyQ1pu9hZCcfvO/Bj74Q2Syr3hUH9kEGpxd1eDdS
j+5mZxh/WJWuHApYjCY5Uz/1F2pFoFtebUH4znZAJuU3yEku4O0HulgvxKfMZyRrXcTWP+8IcFd8
cOeadB9qWZ405DQm3WjkjScEBNxsOszUSJXkxV090T/qQnCz4oauHhIRKrsS4jJLg3W5tgzWZYaA
l1JVGzgIMX1IW6HsPs5/R9dsUiRvFcJ2yTb3rPizdFpzr3qpp8LfH04H2yv6vujVzuU4clsp+UAU
wJcE2PFcnDgFg9ZALi8nNAbqCrXLkfE01OglBgDnZLYhyptCx1vaQHy/zCUSvL/IsCe+h155BSKY
7ZB20xs9cYMk1OjlNoazAhM+OU4I09qSjdh0ZUrtuXFBEGd4P/rKTzo8raI66ZcoVJaiEjZuRyXU
FUtsigt5GYw3pVCV3OW2Hal/fhP3Pe7gvQYOD79Trln+bOtnXnoAHj/gftIthUpZZmNQtnOL3B9z
NmGB4vbO6IpKlozZJjj/bEe7GDqGzRvlxgfIICJXa/OxV96YuitbmK4mAt7ZdLrqYuQwzE5ZRJ2F
IprGNhm1TSySNGgNqRxPBs6hy1hFU0PDRztyEi8UAAOnGj3jlBzzKGwsRyJXZgyE7b6rdRHrm3Ml
4pMHxI4cnuCUzsh6tuQEjSGDWpavsFpErzxN+eVuQCLHejtKheXIt2+cWVR8VnhvsV452/BRLd+b
4Z9jwTkPf4zgRz3zSKvWD+we3yWUQjBt5YE1LR454GgolwkDnf9A16VNBhLtW41zv9rqMqKW9wsV
4FBERz8tC3FIILFKL+7biIW+A83jj4VjEJrBv4kgn+PwuKFm6XxRuT1q5vV3iWHvIe73IKJckqcM
DebqHqrJKE9GlsizPE0Cf5oYJYzIPkuzNt6Sb5u567JR/o6kqe1IvpD1mQuNG+uj35D+GOQ49plO
KTiadtIYkCEdUM2FtLrSG9n+RI5b4u0RE8R4c/A4znTdzwyhVbLMNKWQLrOxyKrMMRxbsW9k7AgE
aVjejubddywH6z/RlI1R4A/TokCyhnNyRLekNsobAsmzffEvo9MQYkbhDd+qP7M7lNde8WyoXwHE
AZAmSmd7zZ4N9QQEbqlmdOEGQq4WSiNPMbMcjuJvKaqAjVoZM5OrcMBlTiQ+L1hAQIdBDj5LI5iJ
EKqXQxEAhvB/zEgLoSmWTJDYqdhdkE9po/Ntfb6cJ8VF1BLMGLmOmVWdBOUxs4rGXFB3yz6XYW1F
VV1E/o0rFzIwaXbTx2j+ghPp71HajX3SZPb/ocOJc8u0OMOhR4kBcjg5g3V5LLOKA2kZ6WqDDJ0X
VgBOqtOAXBIxn5djXM/9iiTjHznLDX1kfg8QRQ6IRGG4YK18LdeAgiaNdC2w6rBXUA8lWrJ6T+Bz
7v2wKhXdI5nHSvPykK/LmnuXqXFpkm9C+UxDn7IGgvxWPAho1901kjc5c6kQI8qFu/nqCacJ3XV6
O1/0ID4PUC0MIU9UnX8it9UH+fgcwY2yMlj4KrqHPl+HGMPdVCgkyIFTVr2JikG5xQuKDxtpnmyD
LXKcM2h+2fbkBcMyRuhmBJYpoAYrWgPgUnOhmph52IfNTX0MPEKyJsO952pVberzTAJolkLEiYyF
ns1JmkHqPHwy+NE/bsy5M7xYh8GGe8d3M7VggR02ATLh9ZaenYpCpbh4qdKndAMd18TuEnEwi4Ja
G+E5PdToLpzPUWWE8BHbGi4/TKZLtrWltRJcwFYHQfxB6tSFtWHOT0KxPj71GQuhHuWm1EndD3Kj
s/n6ca5cw2X9bZEhc1m8VwT2kA11UdmXuCbYXf2ljfye7aWSc4YWnjWGkN0Zi3F7PX3+ym3VzCTS
nQzY0kFRTff+eA+Jr/bRxEphXuTlKIKe63S6FLlKDU/na35/wU6yqSSdj5sFTFR6tj01x4vxjpaF
BJ4ji0ByvG0vanVorGsreK2RVIfpKGAHyTE7AVYc3sELQ0J6NLIDMpr/HbIPOQFdH27m60xyTKkB
8Ktqx6uvPOyHVPQU8wrGJteFQr+2Q10CM54JaKrqQRRUa4KS8EOC9sTmhEqX541hFmrDWs/KO/8l
FXbzD5QSO9LpvMReTKd+ojJUjqdm8+IMuCCcqwr4KzWK2iiZ6VrUmkHKDBiUX794xud/G/M3owwz
KDtyhn9AU0ueJ0UeSGN/4n/MnOAWpHTrwctUhm8qpcdoU5zYIQR6PzLJDSZ4q6j+4phmMNmwT6Pk
QYfiGF68gVllWkUetZ5gKgq9NkFAyC6BvmawcZSwGMOgGfDUTVN7OrQuc/TI9Zirfo3z5jEj/fHt
vULe9QOJIlqPAOlzsAsK1ttzA7alP/OyqGJ+aH/S+/FwNXUwcmTN3+P11tFVWB+GGfRCnBUMwsg9
hfzvB5pfYr/GM0kAV3IAZ4xo7jEVSJ+LHkeEKHAvlhAmAoYwTw59rfvpWCgWQ/BopfoRb8Vt+ZP1
PwesY1HsKEcH9bgzlvdjKH1bCjXfc9LiDuIzMvtSX3Ynp/mbnLrHclmG2xoNOq6uLKvPfLdzTloy
NiMeiRcbbmK0dyiAcLQAkJJXE6tp5X+HVD7kvV98ZaQfJZceI4tOa0m5UE9a6rZBtYrzdobJusJk
urSzlFTdQXT3N/50ggYvZ9q4Ki9vSLy3riWjoqRSxQh4KIuIdoXIr8caTzVjGq5OFne6bicnO23Z
l4YG/7beMamgA8VKPrxwvQXTh3cgK71g5ms4FnYbIU4ngXK5sYjQzJtLVmkZUp29xsLkuxaPvVaZ
7VATm2RwBLEJEWXyOFWsFTfow9sGErcfe6eJ8HbLNXX4bCW/t80aPg6TzH/4GjmY13xpEMjEIAbn
Z6N3a+X+eeX39ZF8/pMNRmGWndsQao8BIEIBwwodNrspz39KgBNAs2Fmzb8MSgs6V7JbrBkeCfZn
cojrDrgc5oddzPiScrDKdaej44KG3CmCJMfeD4IG4vRwnXtwz8bZdicfLb+Z3V9z5ckb7jbuYFUa
x2GVnwc/YtKSF9UGHiI3omFOFBUJ5MVUM5fE3glsp8urnU7Ydd1ZxRAUDGk1ZnUGY369/m6T6FrK
NXEFutsE2X3Ug5TmKo5Juf7wNUugL1o95vNY1uVYUsVwKgBK/TInVHY2N6R4ZTVKAB+o4Heo0e+R
k4PTwdIjgh56cO2iJ54yuVK0pglQ1bnik2b0RDDsshOWs3Dyty58A3ZAHif+XXHIxC+0OjrJl++b
KM9AW8e1STadrnxQrc9ijfW9uxRKMNWaj9jjbX52WP8TreMDl+kB7rdj7i//kF2T6xjUzbOmdPV9
ktA0aDR331UIWn+u7y6/F1dKp1H0cNB4aSVUt6AKHVs2uPfeqZQS6NVZH/+htq/SU+q7WCPh/HoQ
pHlFf7TnegtJ5qx7zUgMCmS630zNcNusPRFhkXBMTffhEX6luv8SPd4MaKlEpKmFHYLP1SSJhuyP
7Leq91Ru7xftiDVm8NF0SXNgjGq6y9Pn5pVtFKmH1n+J0bnJ0VrA+wPqKpvBJ9pXaZyx8TXtufwG
POKojyrrfMN3mITIV9G4f3mIavu/PeJByp/KbiQrc9w7A9mJLORutzDLgfJMIBR7PgZGKPJU+TEW
kb6VmP93NYHWI4lyEWHEapTnJAAPjG/DVPtF3X9y9ChZxQVxopO0UAvsRbpXB8yOoHczu6+WNt52
HMNhU+sK90IMI6gRAmmAHoHpDkNj/U9FcKE0jdYW1LqXL4mur4R5sOqRGhbp/M7GOfbIFBixO/Nl
Nm/LqnbzCph1b4o8ixF1iO0XmjZn7DdsxNfhTVV709E32WG5mBxCUHslPbElC/knXQVd1IwgT4OM
uHSJgz0zrUMQiZQFZvl7PmZ2B+KxmZgMJI3m/v+AWAx3PUPIObk0syC/B1DXNDhKaqag8V3HOiR4
1NiIx/aroCPVRhFxcZPj8vEOBSctyv34ikvEqj7gpNHEmjtZ+ilX1BduG6MMMTHd955cO2H6hxS9
XAfgJbPoLKzzFxiumdRKs7tK8YWiTFI5BtsXtE3WIKAV4zZWRaMhetwCwSwFuFyHfDtkHKDPX/m3
dBFeRf6Oy8pMNF8mrLj0WiANjbukJDM+JlFQ6T2n7X39N2lYhryN/66vEHRKwxvFKTJieWkUOj2i
52RETy9h8jbxrtikhzKL7mxaGbK118aYqSdgys82QneQ8dllxnXGzJMzq8wFa0Gwm89OBHOZxXxI
E84pNUYMwzMkzdQxkTCgr2J9IaSrxBqew/mX8gh030IG5UH1upvUudmBGEOaolclomKeatq6o1fL
ZrKq+Hd25VbaMadvWm1AMiSKsxL1N1eB7y+oTFC942Ds0FFniAolZCdwW2a/3/qn2cxZXdGc2oTO
76Al+bUhTL1s5rkA3SPhJnYyzRwB/YjkDdwF9U6AKzUTcPgqQCQOCpNy5kwP6TpK4/KEgV7F1CUZ
XNBYLCboomIozf69AHv0rmM2Rg0VnZGZaaMpXkw40RbnohhcLtNCsCs1IN2wrLbWxcUuYMfXovfu
PhtVy9OIjLY1MBbNxfl/PEff2nk9clMj8FUqW8eohhCpxwRZrtJlnM1nU4N/sYc4tu1MgNp4xGwo
O8V45r7RoKmy6u7ifqSLnf9A9uZZ8zphuSRiFoR7MaCxswuS1h+jqK+FfG0zKL/dhG7f7QxQpR43
5KiJ9IdwLIJLU/LidBVw9CEZG4mrAyfJXxiA+MioPOrMQU6O51CUGJYwlvcYdfqhpEAnUgrQqF3t
h5YLGgDaYtNDOrUeZI7uyaaw79DYej9aEPoamegX3rTheJVAVbUJmuN3llbCNSHKbMdUYbAXlzvp
2P8tNsvO4VGVRI8sfRA27ElvE6NNOzmiPzNwaKMPTNeSXek5ce/qVBLmBbnRl+dXVHA+6BkkIEII
CZV/X51TYS3pUFWrJbtWJJLc8glR6vaHH+zCT4sqsZFN0eRCQ2lFQk5VTgn2J9jwZqEbh9ZXHzUo
8MW1qld88z+KFag/9E9WJR/lQlVTnVgjy9slTFNwZNtH2x2pTtsKhnIU6YV0euc1fOjZFoVQUTTT
PiovJJMHu109Vl1PhhGyTviqKjfArFxtUvmWtC4n0Y2fvlD87k5AcQbHP2R/s01CWbl9aLpqnqlr
BXZ4iiVCFJ1a7CeAnN8eQSjx3o8+BUduTs/6samwTA7RJsbpRHmTeeCzcDgfDgW9/HYuiUCpZuV+
eXTu8TljM1IE9qzgYxvpBCDX0jpqB4w9lG8G2zMb/SJ7TrEqMeripYO6F+tINKoeGckeKXL9Lf9R
kLoxtoWKyhjBkpyJybIIpZGHRVvP5j3EJabPJSyK8toMLWAW1aGdfTrg7V65Qcl2Vd7kR83Tr/4u
Eikhbe8xifn5B3hVCe2TryixhPUOhKKAJxpDBo2Q8AhSnCw4/lc6+0z4haizaFRfqc18pEAIv1Ol
bKiMUulfHE24PhxB+KxWE0ZZgT8+tuqnRQ1tcce8THSg97xAr4rPAzPJ2aHyrFWnLy3WMDLhHqe/
o1R0gvauJ8IZmZ+VzHzO9oaD7laJSh/qeg7a/W0OlWg8P8PYK15tjhOxBT9iD/55njMsCmOgFjrg
ZlepqMQOSnZQKyh/71Q7S6lTKSv6cUFhschXl21XfJAexi1dPlPvXHgLRZ6zHCObhzOxtIv2uRv9
6zrnetY+J8CMiQIPX3bO/gCU5toUMLfVy67WLl98w/y+QPl52r3IVy3ZanbRro9NqnDOF1DQnhK5
P3W5dvoNDoPAicxSGyvQFjL4Vk0gOYd+7m/B2hWIJsd1+XJxB7etiVQAfE2WZb76Ia9iCFJT4B+A
2Ha1M8RTrfcJcp9qTlEbZemDfe4X4zbH9NXiloNsNv367CB8CJTI9ZdmoPobVw5oyIwhyCfezEQ2
aHJynQdBNSAwSye2jPENLVWiiEzdS01QsevxrEYSoAhTamO1k5DdrIwazWlxLzSEhyIJ/WfPGpJe
N6JeQ6QB7QF0B5X8xG7RNN5fAgVM1WV+Sqtl3wPJgKBqTEZEs3HzKGviHJHxesN51wP7COZNCkxf
pSWlSYsUOEjvVSILoax7EctLeGMrIj5UVKab+G8hWq3e5baq+2jOebHvZroGGJwKHSVooFwPGY+u
RC2D5wa7P1dBzVFfas8jRwqEnhs3fKevgLjeXHatVvU0y7ihEeQs2eKiJGTm816FHMM3Coi3URgY
2lmMumMtKvbhIytjUcQMZsyrZwRThNiuRLfG1LjLgXc/51l3ti87S9UWOUHrxbRoYuWC+QznEie7
HMrs6mTR3M0r/ryt3C7JdkUK1ddq+YU4647NHOB/xPWV1P14qECuaLfDtxFOohrQTWWqh3u1UfDo
Cy7DxRQmNTrCDzOCRbNLRxDATiyD6U0+5rhuh5ejYVQ4ieQWL4StlS7EHmXxkR8u+DFhE4LGHg02
e11K2tIiNugInaCQfJ6VWD8TX40NTKoZrTsRe9tYVxWzbdGpB+ERLsgfE9h4xLg+wO/1unlm2BSh
E8mNZE2INWBXblZpzfcNnMm09NdrMAVRPeznGTim4qTCN8rsR1Ceh88P15IuM22V32hzG5pqQV4l
zc3fKauYXdG+vII1OJ50hPk3wIxFYnfvWzPJqXWNafTsXKbHmHEU9Cytwz54jOOUQo3XSlTpW13X
SnnV1zSydFkHN56qUk3OagAVoi1ryoV3MTSfzCmj7vVXhteDW44PDe3u3b9ye3wrWCWIMUTjgXXr
oMeS81RtCfyirAztBDAyGAB3GJDXUJ19sg+Cf+xRH7qM/q7G9OPBrAlujaMsRhyOmGNAURPAdfpi
xXJRiBBvedFVxSXEGTlU6v7HMcIEOvih4AE3FJm36vOLjQxASWBL0bKZSK/Q8AHZyz9GKqQaIvGn
hhAI9CehQfLVmIKZ/UeMaB887wsN3NAT0PiOATo7StvNmpSpW1bxe2AaeDjHS1MNxLi4M65ndObF
4Q9YldpSH6u1ERbF5gf7VTehE2WGnsVh4MiM96mxbo5JvIB/w8eEfMa0nAz2AC9hscvO5Ct7/P8z
gj+y96C8klcQUtcUM2Esv+6af77iXU3QFBo/Kk8cvs8111Zg3FQRWp2Bo9by+h2r5In1FGI3K+NU
o5oiv5iYh13VB/pwWrRlQfUbw3mbSVlkPdq3CLTcfAk3I3ZaHLfEH39fOIVWqPZ888K9hf7CXjl5
jqefcBQIgj2qcyk7oIamH8WM8/X+hDIW69LOnCDGXUurlM8FFBTbayTeIY7ar0tqsOGt4qZB1zl7
cfaO6TSormyZ/b3j4zsUhIBmQ7qzISRHr7Rmc6AXsW8NcbFPQyxbmsqLLtIx+UMpw/14goVlFoKl
mnTjzvot76byQt5L1DBmiSO1BmcXU+/sGIJu7H8T7VEkYr4tu4jLAcHXZAh+8bhL1CGCRemUWQa9
vMHgNTN3llFmFdM7gKg23uZbd+tFSgDD1Jupj+zDXjuQ3d/smzidquNJ3lyZIxGhTQHRqirS8GuX
fPRGnplt/0qqwcNq19HyZdDftWu6HdGopn5sujhG7X1bJOCrnVRyOU8KRLfHJg5rmB7UkYy2eN3t
Gldm054aw79/TqqnZ4/U5u9r71yrxUhdYfvo0g1HeQ7kyhJNNspy9vE2q33s8WkC/dhL0b196yAq
8CPI9XgC3OaeZKwb+WaL3+wYDM5xKoDeTQ0wG4K9K1paSEoYKFIf/7gcmq2DpHhX4DoKf0/J/9DF
u+52pEAdWJKrOZ7xpv4ERW9xJVpZOjYcTR+1HI7wRJq+kMA3So+sw0Z6nOmaGoVQqlM7/2EaLWNk
6ITrCd8JfiW0zviV8W/nwBvsxobOm2hutJ6dVCcKtZsdz16leeVs2EAsUoG+PV0vuoclVyrgq5ia
wDyu2zKDR64LMTZjuQXxZIeVUpG8feHTclN0aHVPcSXMS9mYL8OKVdl/p46IsYQgG8EDxDT0r8LG
izq5PFEVGe9dHXRpa9TcjAjjp5dArO3Jl2mCE4mbnVZguyvkTgOoZ+s6w0FKVGYtS9HAdOzkfgs5
oUeoMTEkj0J4meeiIBM1uLj31tn1vRKUkuZefrB7jJmoMSGkncCYiBbKP1iKLJlbUh6Dzy+XSzf0
Q04ka3Mo1JQtQdXOIwCIvIUHAXVSU+E9Bd6krpCJOC+jE/75sP+xGXKb1w2ttuWNvB+iBU0p2HNm
UCREkxmwB82yAnmFqAIIW5HaSOLVup3TCOqiXPfsMcvAI1l4cxb/QS78M3AItsRBj2qGMQmMtCV9
bZDZ/7rccyN+hS3xS8JT0hgTlaS2o5vPpqThMJqc0KkXaUrIPvI7mgCtJQZ5s3U3gLz6xjaodN3y
limq3HbAtLWaMBn2tCg6bSlxhO6aHi0HV2rhnRXLBxAfc6ECUryxV9OM0LSDOYLfP0Cmc+XpABTd
nfzi9sl4/hPbvrDsnNNUJJmx9e2sbj1+BpUvotHfeUc0rfuSzoaNu+q9EzuHIvLsZ3N+4vPi7D+z
h+vc7o+vJ7h0oEQxbSiCYgVHIHoJQAqd2X0XwdPIMCPzXlwc2ht4gZaEK1XOm6Bec/8IeANyIfdz
pZfDLfV4A4OH45pXnp6HWD1KUAApFDxX6w70/75yD0oXQ/y17lDspgrqPj5wCIbNLkSzzsq74YDH
Ui4V47yObJazxy5PYmQI55IMWJTrGZqmY1NLzi1pZC+mGBhXh5N0bdDaQ4+u0fC9xUiicXMCVUi9
eUL9vfQdo00YPRrN0Txb9yzSGpWTR+JzJ7lfr14MKN9/8sf8OEfq4xXQfoP8qrDGB6SmDQs+GOSE
L2KH6ctZ660ejDV4MTAibgRvmzPyzXr+3L5qGrq+XwgXRj6FfnBr8JXFSTIywCHUIcutjJB6A8JT
WR5A4YesuOWNbCv8tAANQvZJaGAvPzbRVdHkR1FJ75Kk4ea3NjHSndK+RayfSF2TcBZ5dgXw/kEZ
Njtpayk7prElZqegMRqQAf8VxTqxBelEn7UMXJxVbWqMpfl9tR5RYfZlucjuB18FlG5akKgNopRG
vgye7Atnp6yTgJjmmUyp/xR1Pa6IRKloZZZUnA+fkw68nc0d/m6g36FJSPM1Ym3c1U4C8O+Apkom
08QpFkGeZZ8tuFN+vcEsMhZiuLj04ToOXrRKzFITKN5yYcFh1XIni04NfjE646tqu7zicyAmkWG7
pEgS0woXTvLtUwFqXhUVZgskHKj0WFnebPoBwp91ImNIxZjgc9hA/TaZQOMsg95DMW5A2rG1oPzk
5sFu/EYfDwKiLKOXu1TMvI6vjEGtgGMdaqBDktn71cNKBULlVNFFta+4V+nscKEQOhy4OJCdKF8S
H9fgE8DqOqeL+AXb8XV5SDnsZ7t0F+vPoWLP1dkawFOQE0hSginsz38HvJOrE0jFTCa97wOusdyL
j+o25K+d3SkkVR69V9KUzgSpbqCPE5TDurQSViW4kq5iiNfGosQExjJ5EZH7brOpV/5XD1NQ2z6g
g2/Q4CjWYC6LbXSoznORvrw52vOKxbGDIaU6K1v45sBgR1KiQkQP1QLuw2Eb/3z9sRA7VWItDscD
1NPFYtEt4crR4fuBK5AROG29aKZw70sEbQ3Kpl6d5r7WTSrhPbTqW0LK9NrrJF+hxM0QLJGlwiAb
Q9pQOXRPWqkeCjiRnrphRgTS0mPCWA3TCqSFBErIzJgo2pxpjnmuSb9Ao0XmX3jX0Xb3eTewfmKR
l3VqrAsHej7ffvhqsr1MPSYO4hPiddzYsPra77gRo82r4RQCfOOYzvZFXmJef87YY9VQIs2+0dhH
pLfhgG52zUt49Wnk4JVSuspWIc1KwvNNUkzQV6WkNB5zxn76Gelm9azVG8+7z4ZPnYTuBQng6QfR
8rsK3ClNnaIFI8H22UfgrODhvPnyhHKslREwkIsizi61b7M9poIkcJC7bPfw1QhiskvG6xehYAAq
Bl2rTISBVhBnOlvtvO0UmvNMkF6i44ovYjDU+JKTGTmVo8/NshaTi3sg6HjoZN2JntYPwd+CAA90
n4YaaP37iMQMmUc9uVTZY9U/NV9/Ocd6n4ID5QH8LD/W33AVDunJ5G8CITYMvvuxG8qmB5ebuU0p
FkxKt6xGdTlXZa8ubEA6myfZW8BQbH+0BeS22mDzsYpp9R3kUoKnrvK+vsXUGMI3rpm0SqdiJkJR
ARh7vQuC+RLBho8mDHYEkD0aPPcov0slnRqFcDI6deceaFWtfqydhwZSdMhhs1h66CtRhvoFprPE
2v9qyRvklyUtcCeRAxX6ssabS+EdvUuBtFR//zNHU7eXijXtcLLbOzoW6wbaSkuyOJHbllGwQj9J
4bpte13A0WVP4TAXRXtt69r8VmcPn+JwPCPuZzBMcza43zlz7lPUf4AJMbRIBOsHIhaBxVCwMxid
sMPZwHrPG0VMAeauJnoBdUb14K/ExyFbqz1d6eB8htU/nzGn971r0nadUwqnFJFmGtAdKSOjppcT
LcNfqv5LcgerkdMzK562hML2H9Jg1asuTs9K0lqlVSFww5iHnVbFzqXGp5YDsLjGFuuyorpkxDOe
11FCndF4RMnZHgjMsxW4CFeaCzYZ1V16X6AdWYw/WauXTBLBTRL7k2VOzjHNHqnIiagkbb+oR6Tj
Re0AnlpPqH/v/1uZNk+BrESd9YtyPTG6oYCM9b8jifzVj6/BmgBHsBap8EF6ydiRdvIZoRF0u+Sa
/8qMFuadAdt0xQeyQU2FAewqyA9RjE1MfD1/KLjq39n/Rtt3lozs02OmqvV2TkyFUfE6Qevl96ZN
5D1ENKbpHX+HdFGgt3e89dHLM8bDTkU6kFQVQHNFrZG5juYV6LEavUPnDHGZsIVnHrAyEZMJanQF
tyBU5CUi7KxGrXlvyKRTy3tmnN8vMrHxKnL80Dz8MLRSEATiWPi6L5xSfxKO4NiqENfQ4eFVYkT7
QIovAUMz3rRtll50i56mdqAjdxes35gCrZf0FFccpWr9A8YXDIfDPRils+t4T7zcQuqtHxkVWSGb
bhPODprxqXdnkoXf22M28YopDADGNWCJ9P/DqAeiLfmMcYCEEG2qFSwPVaLgmrssiyBy4SdoFZbY
ZetQSDnbX3ZuVEYuwjD2oqAFPTr+dk+siFtMcvOuWs4nqwsUwfxu7vZPvJ0vyBdzreQRexTWKSyq
g8B13W80byD+uEr0iggJnXkMll3lRXfx8Dxkq2JSafn/yx++kpyi/AYb0xDExZCQj+gh6kCfIG2l
9YAwh/2Jq5/H52BC8Xz5dSQD29Ry6sSkUnUtcnzU0J9Czd0ErLpydiJCaWQWgL2eJxrv87UrTQoJ
75YnVZ0HVciAR/01XQThD0f79D0qyNadfOH3ASS6qiOzJX1L0Lk4zVWWUigVBuugnQJPaqu7McM+
VtD4FNbIbC1aVvvjLVN6wR/aIIaVHa37C3JFbbeUXKasV3BVNZsCHNa6JJxeUk4XUludt4fWCj0o
c39J3YE3JaGHZGUSMuBwd7SvjDT8NzXQ7W7TZjNFBhD9f+OepNCnbCSWMsYaWg1/iQRHgaw4y5C9
BbOK1d19NfdQTtOk0CdFA3Ap6/tRCKchiKLcS5YjWBUafaUFLT1bG/VsuglgByBBe9Pk8kf0IUih
Nztu9zmW7O8fUap6OnZHi9baz6SBoYM9as87R2Gt032UyWZtFdaZ+kWSdF7GeQX1Ir1NncFo1uoX
R1C2buzBigHSfpGEdCyx/KC1sGe1ZJ0K1DbinIE0ne0oC4p+3AuVETYUq249SiExLMlFdMBO8HEI
klz4YDKqoY/sAnTCVl7Ap+MLnpuk3HBaOhoGzHHa3uVND/zYnJMNhedPMZ0JAfB2Bb0D0+BnXM3q
ffn2UY3CI9iy9IxHq19CcjHSWa+PWijb4eUQYGED6I3uGb5MRNOh8jO2GfpSEA36xwi9yxjzdCOn
RZnpJYoGLpP/gqRlBhiSUcAkQogWjgU9cvs0UiqN2s/fPuNmH/CdgLWlweAUkycEuMPEdVemBAWp
4eMuV3gEh5tBFGuKoT5G5EysgDq0ZsNjib0R/fLoY1qpnPvBm5tGvZdgS991IrH9KiA1isPvoY1x
UQPQ/0QzGluMpRzw57by08EjLYJ4ZYDFvCOvOY7HhPKUJHV8PzRuWX0nyNyDvUK+p4vNiPcioCVs
S+d92EpvoeCTqGb2t6XpR/8RKIlB/8RdMuRsqWPm03oFF/yYUr1djqMgoxPccR1JWF6rs6/jM3/s
Umyy5MjrX+UxOlsMMyfruV4GaCDkXiz5KlcMCYMKplnj4ilQy+wbirFB4lNGuozy+m3yrPRnlrP6
6ZqkgAnJ4VHdFskUSwy8WT2ClQ3uV8r6wXC1ido7qBPFBA28z4ltxsbXtZwC14H18wZEazDDE7BW
5zcRMdjdY+nY2RGXnBUdOXgdA8NKaoI1bGDXGd5XtL7YbExCyZ7j3ttLWvqCkNozOJvEdtdyOloe
vX3DXL6wGzME5DFzrFIAs7kfo4mzOcjzht/vMxqCA4Z/1OPM3MS10LKpA2Q9Uw5Rf4bj2M8Fu/1r
ILZ2Yhe8o/1NK1HswF71KbFNA1nG4sl+fydyTkSh9gl+agkX8w6qRu20kn1hcP3+hahTngNDlZM9
r+i1n7W/G3yo9iUQV7D0CuqGJm7nkHG3UiXVg6d0yha32YoHWah5J7rh8/89U601e6zy+lLSMITT
REeeZI7POCSFlPxBisVjQ6vmxm1kLKy7dZ9DhqEoA6TaPyOe8ND7nfGOa+74sz85DckIy3YofFLI
z4XMM6Wlj8zvyrkzFg1FKWn2P42Nnby5TREiAGFqM0ugVbx50+nbtGzvilMY/cIZYboYm7OFqn5H
L+voJ5yKhSlFjo9r3Mau5IkIlPamuogzokRm1aYkCCDPHYpKYnmHqeMGEHiFZtR3aXZxj/KwfLQN
Ztx01EQk4AAri04+z1eInJ3Mtn9DMphim8msCyyKXwdeJGWBfzTvxsY5wG0sdgTQcDkW0ZxXbslp
OzCmef6xlBBRwUwpSNlnNOqELNSndMJwNCenk/iJheoOg9XH1fVCbjGcW4jD0BvkDDKGT0i78HoI
/l5brkHDJ4bi16qxlPHWt1BoD5s6RL72iHgjdJyGbxg6pMz6o9n/WS03ezLjg2D6ZxGc12PYNsht
nHxOqAEngCtuc03HFxazXHl6RTnavYxQcseMe2NrVYJl4tBo6M4n5J1/+cv2g2+SPQe2lD3tLPca
iiRCXEC7Vkr0ncKg9bkjG4IA8cE1oqObNfyonVToz/tj41H7KtuRdCfucrSe+2usLwJ32BbFoxEh
KguBnBTY+sxzWTZnjEvKW0Vmg93k10x+5Qj/yR2t98qVRnXEBXyj2p+OAtM5Oz5UUjZlB9gyJ8h+
vFmlCSDDcC/SgOve5lfWmjiaF2OE0gG4FjuxnWrhyAQCwILBZP61n7+XfyT9ZZ1Vc9JdSDESdmUj
d92r/tsOp7UClcjVdAh99duoGkV/pWFLVGzadaC1CPzrT+NyAeWYNzLXjI7M5Epl3VbKSvG9GvoC
SFwRXJdM4AGdzWtRwrlzD9myzQaEzYhle4XIIiDjnx12+BNHFl+Ck4XdCpUtDlJE6gFpMdPJzLWQ
56pQ5Ltn3bnIwGye2SafrHF602kjJ32H8IPuhc7eaSesuBRCMGKbAoeMEKACH5iueOCn4ChoC/MY
e6owoUxtLG65Monb9B0NoeQqz/YLsq1cVguHnNzz5yopFND+5pJIY3DkUM42zs0GIzrQFv98oC4Y
KW88iW36i7/5xZzVZF0yY3cGEz0RjcCOGsnGP/FNq0rfRTbBlLH8cn9AtYJDbQ1z2UzBZaCzfAu4
v/QKK2+mQSPbWX2MWWSIFrnsJH4scE0BJTJDu4VOjQWJphB+JgqJ42DTt+SK9MUXDu070KRj3MXi
AOAYS62ILZPvXF9uDugLj+iLu8HiTI8h4ZBNtRloJ4Tr9GwduTsStBSk42OltWJbejev50hnMKDo
aSv17b6DzMzdyxGV5ADUg6G0qm2zmApOwsVyz49v1+Db6kleohakZ4Zn/YhC4ie8tgz8T1Cqd4MJ
8cXRCkrv5GO1avRrmXc4uG48Lp7CLHydGL+6Zce+d7VL/piEdUZUMQ9uuteL6HWY6F42UtTrej+V
xwj5+FK3GOohUKrFbPZO2P2Kj1AANVO4z+xT/mirNL1kvkZqYK5nLrPsGEleQR3r5W3H8Ah4LZeK
sq992NcX6N9KM8yORENs1z9VWWyKOSu3KRcZK5UUKss7Jg2gAG9Dhi1WDhFkwpNaRWxC3dN+XNNL
QS0aBPuIsQW6ffgL2LNOOuFSP8CS1UUlnYZ82XKnM46lLNdqLXyNWW4m91/bSHwhlHLKUnD0m3x2
ZVkKnxwRFm1v+mtvgNGcKn8UMfhJFNqbRoBnmpYus8vw3Y2oscpi6pEv+PlWAmEwrbcIOuRXKpAn
J6a4kxex/5PsdmYRVQ0iIYzGGizKzjeuskppRfb7D/dLxZAiljjUHKvpG1zgCyTbGsNIynQH+vEb
P8Zs2jaSBl7lg5xnIMKyi8566CG5I8Am7o/jLQaSKdWug2Zo9RffAXAEHHunJzwFVBJ22DoKzQMe
+RAMiHEMk8KHOQ9bXDWUOBQtJAs+RinTNa3/gt5qA2rJjhCdnIDVAcrKzyrZVZphgLG5xXiV1YD1
RtXWhBRjYE5OposkC01QLgMd5TwKjuzGkBck1zumhlT61XYvp81YPjnFRIrhC0lThdFq2XdD53iK
5G7aHpEsJknLBpIqshGQCfw5xS4E2gQxCKDOMws0M3zk1UoaME8if8coJQEvCiwF1N8oZ4nOlkr3
XAd2MBRjOr5VJ5xD0PE/MUGAjViPfLcHg1o9DwGjMThWJi0T+hU+hg94Rz2q113zja4ft1arPEUr
qf8PxysHXLwfPzvMf+WSN/dQZbpIKLCZmXZVqaZleh2HQYlSJ5nODcOrlUYXkJa1MIJ+BZpDcVkE
FUIu3Y5L467di0AyEf0qxU+JSrdTQZbOA42VINhG+GJrc5KMJ8nbqKTj1dWSaKgyqk57vLYxtnkO
QN7uLJaXPn7yFFkWNP2Uo57Wl1fGy4clxM/9kFSyYC89j9/5gkBbcwKujQfppECzrJZohNfAfj0E
kkCOMg11ohqKxZnQyXFHmBv8G8vgw6J9uc/7Csk3Me2XxmS9mV+isi8KUiE2kEuX/vzXnjqiEWlD
VnERdIkJs0iYcnkpn30rp7tB5adOfnildxk1aAILgqXTw/ha8U/lY2RuB1uF/zaTcib3E925V1/t
5dLhJNRtsQPMgZHSQ/08x33R5C9nsXu00Of7oypkFZ06RrShjiSMprAfxJKBMDCtnJE6KNcBXJVZ
+x6YdwleV10AezkoICGhXnnntYPbBTMXKYEf0Zxjr4ERl9ibt6QqZRTu6VXyYbFMuwbJmXv8ly5z
MOdvs99NFlE4f+yRSGguLwlAVERocZtsRySOvMxSB+b7Q/g0qJ50uZbRrAN9nQZJdt/iFuzNy84Z
YG5zKlxAIgHuH103we2ODYhzg6pYdF73whT0gym4fXUi13Cq6LbNt3ZkkJWxokBOmfcsvHXQdOhG
+QTicKZXpXL1fBpXe4WWjhV3MHTMm63FVrHncstigzDzv0EqaTAY1tUGl4/Y/sHtMKL4/KpL8r9F
AmpwzvIk5At7PI4D30JWY+JlzYDWCNvZ/RYfR8dJuKyf1a/kW6+5VVbkgrxOTsQi52hDc2Jy3CXJ
7Nt/rkPT/dxEE2vCgbeGWeb2R8mxiRqfUINbjU+/MYAI21lYxkM3w79Y2XYxUmlAgWLDQE/UTr/2
1v26mDeEly8BXiOaXW/Omtb9datt5syyMdivQTFa3BwLu79VXe77rlj+pEswZj3blssHwOI/zKlK
Nn5AMxh3sFa0fEoojV1aaUNBwMJDpOXQKmuOdWIqUq1vKleI9a2KfzjocEOayJ3v0aqxCzgsjZiJ
AavWdu/3S8hI34OshOb2/iD43G4TWl1q8M6IM84J0nEohJncdR5aCol6rxHB/CnaV3YYAqPsq4gv
UAgOw+mqDkAnQTUca5Lz0Wd1qD5ITyIDpO5UYqC56aUJaJmOZlQ94jLTS/832ySMHA2Bye1Gh+Ur
eaiGfQkya7gVixf1k5WvICaH/R2zEQhQsApooZmvgNQa1M9D6D0D0Ro8shyArl4gpcpdH1UQLv9W
03Pm19azHSTNXpo5Y7naYKqAWG9jTZGRMTJz2u4kQng3iiXCDDNC/zf5qxnjAiKzo/5so5MALFPs
Qagx9Y6pagXrOvl7IVqB4E+lUxWIlgXa/uMtFsdGQwjrC81ULS9ieqLb8KCAb1FxltsJDvc3r/3T
/go4fhaCGDmeeLWCHW3sTqDI7pWQ092muvpFgtMdYHl+tWSPnuzpA072X2oitZZHp5aJBdnyM9TN
mcN33T8hO2KKItDqX6CJGQljZnlZ1Z+EJKpt81PC/Eqn+d7nfGQpCjAqhKSjkX4k3NwLTgDmNGVi
9x61Trrise/shIfGTDKOXOB+1KSSVqC8aNSjGkYK4J+IAKv1TJCKs38SuXJUeStnN7+5LuFGasxY
4QGHeqv0D4+WMEHQ9Uh3tnkPklwANicyjPokPSYxSBL9we8eOREI2cbgj8t8nyHeOIUPOYZOL5nR
AZDSLUTBI5G69l9mJbHrFIUULfuNpay9aXeVJGv0W2b4uFLSh9Owi9MsXvON1rq4a0r7KVzxXgxU
PslipyrU7eBg2qNhSKjYGLFYuqXhZ3q3SOh9jwTU7cHa6AtgXH1fJ4jbVqO2lbKzRM1TV22LTBsA
jos3n4Hf0pQ5ekMzMlr54aR763/W25X/RDiBD3CxI6HvHUSp4He/8u3iWSNwxWCGrujaN85uKFva
4CrB7RaijYJDSGdfgjCI1ONDBdnLe6sy682+IukARUcK9T7Sg0CwwCgE4X+2aE5NpvLsVMTPUeId
35ThnTzR8tIJy0v/SXsOZwpkY0zkC/e9utfU+nYeA8LHUJHoW7uU2Wnyy3wzKpGw5BsD006gGLrJ
dWP6+B3ziVxN+s+S9c4PfLq2oBBXEGjsB03dV13NvoqWbxvj/oH6DZrU4flKmxm9TXOQ1g/JVAO7
dBsqntHvgqqcfpVOsLnYCminaHjz0p7hbuQ4GXTPQWgxAV/hpL2c3S6FEuwfAMBHG+jIp3UUiRbY
60BkTd2gFPLL219lyWq6kuAe0Z2TlRmGuFwkFybKUxz8HYUnZdpY0mk3fb6VVEcoyEQdMkxI7Iyf
eazDcOo52NnCk+wiu/xds/3rbuGAn/J6dpzcM3UWprjX9E2j/UygohNpeLRpEnyVstjU8rKz8aGk
K8Ft8ZX4kfmK3x40vKSv2yr6XWZWx4dpPZO3NLy4RK6NXjt14fve7JV0agsgBshbMz624lzZr79t
jOgdaqyoN7iqwRetoNCrhdGMZDI184dp57R7UwmHVURb7JHtGEQr/nWVkUvIKOpGEAZCjCPO8lF9
z0hL61f6gzIdNtKXwKQufdm55UIC06Zz975VYF93laWfd7JON8vL8rXO1hcQRB5YciL407HHXpQ3
E5Rf2xVzQ/hDhSrAAgp/16fqXlBMcFdYIB10IurEVqdeFtEpGu1xpLJd17Yn29/cw7QbUf2NF0Vp
QSkwihUjCMuOJcanr6B5bSJq8/oC83rRL/GoNpB9kNJmUps4egcL3yOcdfJyyFhrhJ3PqO0f3zMR
ExhlnInNj9LSKjBzP2KPiZc3GtkFY+ysawCGF4O8syHC1XJ7WZzbL+sWKZCfn9sIShQB7abFWExx
4xVQVnc+mDztqerQo35jfp2jIB8D5oT4XCsR5FeqcuDAOW55VDuhEYDpBgiKWRjoCq1+lwcWNnTk
nlIfmvccUIS2l23WH/08gduMflCaT3hYVNPZcza42aAYo2IH4MO9xA8H9X30tJ5UCLdcquVr4Npl
J3afzTp7RCIii1W/wGHK6gC69dyhGm2owv0dg4GEgSR5RYCgKAzuVQzk6HRIjCqcpAep1xfNT7oa
S6UhapF2w1xSqcWbUTZdNsBD0oTRdKsLnNjbueoXIPI/WGpOEfnCR8EETliRnbAIWVjWbg8yNMLh
K/VaC1nwxXMvGKwtX42l+0/px9keFqSzMezx8UQ98WMF9Rv70W6ytfqsrLnsR7gOhZQDVWIhEEf4
6bNIApbfbU2b6Mn8Zb1GsqIdmh+Q7/w+WGBHQO5spn7nRVLgoq9UOv7ddgC4CW1n0KjacvOx9QoQ
jsZcJxDtPoITtWFL4YVbJD608w5fQaUtMKy3zbdc/hmPnBBDe27g2yRqRlEFmfX/JmdtS09CBUAQ
dS5lbLQ1nIKdlJFGg0k7HzghLJUsnj8qPrCRtdtLPm++f2SlkpTchCffUnZrnnAqm45i4EH3rOV7
PdwME1gO6+Pxkm3HRwbIyGo7M9HYfoYQbjhMYh/5FaJ6j+juLGEFA2Vu4FOmug44f3VYxxjiy5Tj
lDHSG1srezSsvTNrdNbBlKgKV4U2qZ0ucSvuGcRAT8FP6qai2igJrW1mrHeFp1A+jlD1B0ojPWXh
rdxGJU1skbtA1G8GeMSH2B/f2232QPApw4gkjs8p0UU+kI2WYN5dHQL5BF1AhJadfTQgf/3UQ0UY
Do5KE5ynhcaysdrGwAH8Y7pOC99NJtbAgLmwV4lYIe5vZf5kqYjX45OPVtgedjKBpAEpot92YO2e
6H4pQR3GpWqBoATsT6WVWFMHNw5j21dBGUvKfGRle84qosrwsK64OZxNL5tMangMgrUACBbc1+FW
Xe+jJtziRUlELWJVWNWrIbUm3J/UqEE/VSXYdKo6HZFHhzOpYYYEbJvFFDIYl3xkCpn63PtjTQJd
m96YnyrGktmxAB7GpaEhPR9gNMpVmEtgQDDb5kGpQ1EWESMxmZu8sgVVsI39xw/dAciRjh1Epi1S
kwj+FySoukJC7XZnJ8YJ3QxnjV7gmSqySwBM55NNpAw71b0YQNz6CnbpG+TB/VMGaINJxJjQ9jBm
1YHL+3kwB8WMScDgQsobVWdZtNwwUitp/fiMPNk2EMrsYkFCjoslpzDdR+uxu+zqYPtY/nK27mwG
kqFA6DX2+h3FxXBmcdbUNmaNQ+Z5NrT7kaAiC16tD2hLBZin6zaCkUtKXKdoE5r7lW89iUihLO0Q
f+XXqyJNZHdrZoX34NEpSnosWWkTIlsqTaj2LRBDG+HT9PATMyQ+KF33dG7O9trpgsFdmXmMlkIx
wvjf9MVRO2/76Bmg9/jUI1qrsOchXH6FvkFN+6BQNsv8bO2ckBzXqFwIWiJZPHMDfntAtn0sBOJI
VERDnd+rSdOpjh7fV7Y1/qC9W1vBkbMTvMCzru1bHTs1UjHbQAs5X346lJZfUq4hEYzFqEO4X1PX
m7QtlOLAyUZledx4dC1TzEsYVcdsXLkIaLWSoBU1kILpe/HApPXnlGURln5LkjTol4fS5bxppi7u
Xhr0VyRuSiMZ6f2Y93ib2+oP7rGsNnXhyrLojnlzyM8nAv0pGXspHdfwpK/MpBKYro4ENZc1enCR
yScuQ3PJYmXZf4NbUSzuq0ywmCENCD6ZOcKwNTowyXioO7SGWQLELJhRCRTvzMHyVUit+tO3imCT
P10ydgp18NU4wkB/HDecW5M8CLNl2uxibn0oxPhopTrVhzjbOe9Yqkjrbi7X56XbvN/Q4AvmfW60
bfNFdgE3LH+GL+gM4tY4hD2TUhUd3uGSaeNYGxZgSgkVG4MD+RD8PtEAuymh4hMOGAEhljE8KB1b
AjVVv34Ho18VUM/7LD21BKBcWVOgJW9cubxqUCUjn1cC4+3k29kNgWIwjl/nUAgMcFh2m01YVBOJ
JwNm+vxZ96Dbcw9ZkDjaE71cwdrscrfY2TRACJ1c4OsN/sLoBKyMma+z9Fk9Diikz5C+gml2iPhy
/Ycjd9Du7tSeOzS1yXpi9OvVZhFs/VlGiYNGL0hn/UjQR/Ci2UhIeRrQ6zrtzp3XG9fNXLhXXn09
NH3tq7thsF8UO+hSXpUK7f/R8q8OyCbvzpjEt4GmaL/fPuyfbjNd8+Ja9eZxQTVhcy0ivW+INsQR
eBV5qqUPkdu5WpoW6LC4K7FS5qHN6c0oRONeUSmGgyiF7b1tsdvJEtudn9sCAOGHfaCIdJ5VqkDu
f4PB69xXIIu5PoK2IrAPqhGDoP+CryNJji/tC2troT8hOlKWFjQiAYYV4TMgY6aOclUWZSf67+OB
5A1J7pSi7VqBxKk7tF89TDXPVCr0uVBRIj66ePpjuhYg1r6MRCLzG5HzUd94ZlFNdWhPYY44qevI
qH6812CUCnvwueVH42nzVK1HBTl2Tu8mjKuHqmruaji+VO7TTdgfyhhTkkjA7++d8/BV6T7qMF5i
Kt5Bvm+rUE0vvsdcQALCFyIbBnXYBxTYDsF8czPZrrRWDrD1vnZqAErZtoq9vnHH0qOjN1eXzM8a
vj2iojDUZa9lapDCTQUY8+u1TmM5s3KuUs67HgkeXiHl1As9ajSQLp0jfDW7LsBZTacuxulw3Bht
slGid0Ws3VsO+spAsEPYo6HUThCPH5aNXGreQKtuPoWJjHmhj0fGVfIERWq4coWt5B0sF6srQxCK
2arxZiw8niwbJCo5dCmAZpqcDiD6vbzSmVCT9WOW61dJoHJcF6yPh+i3ubff/Q/TvJ5MHDmpwnxK
6qgC52Z0njsA7OLjBvwg9ssR0r8ldeCTdHHAzWATM/0aHmrf1r5f2fR1ViJjs8HBMBg2I0F26Nqc
AJ4ISJPrFisNkl0UTKbmZaonkybsQhtgOV4Wf3l4PGz1aDuHjy95PQ3t7gOG3QgxyBT0PuoQQeqB
NXDfylmUmypeeatte4dgf1zWws/iq33d2y/20snCwKtx/Sqlp4m6xC5xc9Hh56PtC8VW02xDvn9K
/qF/2MExbzBH3ObDJALy+tM8QNmSTZrcChz120wTmdzeMZMPXa+paSZcpJOsANMuEiDfVbgd2NhF
G2gO3rQkVSLjCgaTeP+QcP/ABANz3V2sxX8+RLHz41F8bXLqDmJWDf0gr3OEqK3w4xrIZGFWt4x3
ZGo4m2TlLnwR+CjXkke2KDglgXuNvJTLuzbOBBHoZC/Eyy9be6NrLn44+XXBRjPDMC7ko7J0Knh8
xwdHe/SX2z+cpk45m76YHtjI6VO6tbil0vUGSkcSZ/JgfVRDL/yQvQQx83HyIoIc+rXSRXYVaRyV
zvmd3xgdOsxDYWuGX1Bcy1FobgFrE92GRiDCreujDu/izWPv2ugzT/slSBeoGrxVG6C4v7N8wi2Z
Pf/fz8jT7fQvzv1II8oD48OFQYYTVnf6e7TWyBRRGL0PJq9OwL/cLexVKIvlQxuVXerFThEIBwrP
TbDyNRzeC/TiSHFkDgwzyxOZdkH6lRWMfV0X9OmhkOS7SEOPN07upef5ciVCwT82MgC8nMJkB3rl
ntTDo/dxLYPcT4V/TNpESeMC+QAqInicTMoQLIE/8TVKZHVQY5aaHVy7VTrM7xN4OER1X3euUxmZ
CIz7ZzfD4qkBKYHu34waF5W6hCZRwaSk5ze1lmBZQsZc87MWnjM4sN+371fNCqu2CEAYV/RoQ/xx
Oh4ogofrBL3wrJu4sjNTeOvTKkc3CooSuP7T+AyuBXf9otF1pMn7m5Ts49KTy1avo6Zrko9asX/3
Pojx0Cz/c4MiARMTvrcD8WlVA6RfFvBmy2m9InOoO6FYMzqY5Rcb+V6CvqqDf0aLtTONw2LE4mmX
VgRxJzn5ucQhvvrzq7etJj+taNwYEsbimO30/zdG5q7dSzHj+LxC2+mFxR1kGsZjfVjFOAICDWWm
EVzhnLQa+LOJMz+poLhuABN8d+SJ1SzxBYvaXbEnS9F+y/MgLm9+T5QkE6X0uArTIWG3D1c4FiuH
GpE2c/Yr3xo/n2SXBayW3nHr1h6JUNXC//xzb+ZsPolCUl5ErdeSospvglikxykAM1Ady2ADlRvH
qYWvFIR3HsXGJ6XYvPrUEQOuHdXyCmJvvSCvrwjWVIlAHo9+RS7Vmi79XEmsNm0KkOD5gHzc1jqF
3san3tocX+sZ9ydxb1E+Fq5zgrCm7nB3SlGmU0wWNXhRTcuHvt48gmu5jofmHyqvR+y/TasTwYr7
dlxIuSWuVlQ4Oab1sf/EDoSgnDw63N3H4fGMxJPHr9MSsYF7Mcb/qkkGPBhLsOVaflecK7F0e4iZ
iK7b5eyVu3prlQP4w/WMO/le0NB1l/rIgsunlCf1wKUx9pCmOMGlq1Z2CDnnWzcCMl8Fqnl0n0nC
8ls6e7PLgcWx0bRDkJoNbmptmxrMR9ZJ/CBxJRJVfTanWvPwvzpKe6H142V+p4cugfWF1lL9QLs/
Ts5396rAYY0TRXHvilqbAaHswYEf3EHlCmaHyTQKiUteIxNtZCigLnTLuShLZzCgLf407juTQpow
4O+33T/GQLBb3peQEN/Jolgh6JHMrjhrd/EzAYpZx254dK9WjKdbixwzi8oHqXg/8g5kOGzuNn0S
t0XnaGJ53AKoVkJakOF88BegQ1DsPFdqhdYAZAOTG21+y6uP+HJWgC80n1m/fFQRP4xKgKOHXtTf
GzLTnxyzXSylvsUqUfP8r9ZAmfAWk58lQqphAB6cyc1OKpCUlyh8G8utJVfr8rSECGhHZT2abJ1z
sBnNsbwwYCIqcR2dr5D6AkeygH7+uUFNjnzvBQ3vHxykmbkpXcu6j7AXUxII/JprTTrSoiK3uZ3g
r5oJLL/vCLlza5Nr1ZdbtN8pqeVqri5ATJBinQzDh92/P6yJp6c3XHTvty9CCP8qzJwOhIKOrQ6k
mbf0GGgZiuaIs6OChSPvJC6WLZCRQcateQZHWlpkHcJVj3cmAW9uio3WeypLqsvA9mwmVlw0ETy4
h9O3thVPIK1dBxMmkLaGzCG8yFB2uXT0+gpeh9kFpu00PPe+5mnM/WDiD3f/7PvkOFPvwvC24fTs
Cd8j1f9vw/QzJj8Z3tqBgAq2VuPxj/QhmaL5wpNp2LAwHMFM/kc9E5+ds3pkoywBsR2TZUP0Ltjs
PUfqEyPtKc/uOmRUTLrfPoeAiO+MaE6O/B95LLmn9Lzll+Ikv5ShOG3iWNeH6oga2JWjmRk1RIp5
QxUD5EAoTqkhygrtq8babEgfvtFtL1OD9tiTJXXSIAWsEjDhJbBXn7yty7F+cuGx7DMp342dYyLx
KHf4AbkQsHBD6CqH9GIViUYdiMuNgnZfdkjv80/RC78Nww1IK4WCCTQ0w7lVjcf8guekLQRlNRVW
AkMOoemoYN4tGEWZIdPoI8SGKprLhjFc3vVGA6Ix3zcwh49Vb6PNKF7g1o4M/QpyPZ2Cn5C0+JbH
l5KxaABZUNuO51/IIWKfuyE8lPvOfBjtT8m59KPBU+AFLchUJWZbVHl1nQH9s9sfvep6UH6k5aw8
e+HPpVQuDcpF7kMGvBFM7BkPnL4gkmXQNAbvRuTDYyt+LxpPYGWIH3oIy2vhsCpVrOfcl/QQno00
qHHAkJohjVu6gzji2cmrtMO+6N7Xa1lLQ7L12eFsbvSSPI685q4eg9doIhggOxYOEoTwfGqi615e
+y20mnzyljBQ4eGdDVrWFS+jJabtoP5sZmQ98ZuBiMQZ+lNE2t+pX8JDRWysMEyn3jgc+f0idcYK
FnvdN4UZ4l1DD0xwiqHDc2uZfw/8rhCu1QyfVf088uljfOifxmH8Yi89r19PPP9XhgnP0l3jGF8y
Kjw64is0gHouXaCF6X15WHt490OvhD4oxyoTXZbIJLR1c9chV4ilRKP+/5QEQCD4bzdzNkvJwUT2
jKYLqSnJO1fMBwZ1yrsjWAX3HwuSnFTWcGC8tK7H4OHL42yH6ihAr83REaLqHOS48S36tQX3ZGSQ
ByNQz0C0wvLDVlaNozrd3cHBa4vCZcOMUFnW56vl8OzTi03g7APZKLrIwm1ojR5XtJDfqINKrXc9
lWUiKC+RQ7dNRVaNXZvFNG+7haLf1D2SHwvTtswqrrcETZgb0406VIM4SFfvgAAkpXkco4tOUmG9
O2PpbcfkN/fsRO3iuitS7tYijfvORuWFb+bfYQjo5JKZ1+/axkfH5mfC7NZP+yrFJMDlmpkwps2a
qKfOqmOXd9FyL3eyzpsyzNzUJXfM+S94ujwJQ3kZGW6kgTIx4SRyrabAtwQ7D4W7z2CXU6T13EI9
yNM20NNI5H+5KWU4boTzJ0uXrZqgq5IOPlJsPjzSwf0k8Kp5EL2O6k5ZkljpHdZ8SQjeGWDH+3Vp
URFNII+4V5oklpv/pdTbbzwnrybwRsb4vqL3BZe9PKv9AF4RUm9rBp0jS1umBeWqrDDEVbUhGjjJ
MgMEuwwy6p1+39NUAJKsaiSULub+Pc70P/v9RXngBmNqUVT6rPy944le9Os8LcLE+dWkXLkxLD92
atR/Wa/0QuSAXqKBg7qw436ya9KiYVz2pYjEc1S0cINohHD39XZwNQ/Jg4D98MmuJxpA0fPkgynj
ErBx3WPdSy00acvakLo3MtnEPXY7y+/odpOemtsQaIQFG2bOFBedlahgaOTPhiHzcA6eydjV9oNn
f90ldB+9piKqP79u0zpoTfnSEX2sHKc8jimPtAg/Pe7IIgaHQWkhV8oV2icgdkcTLz1dyq7PPCl3
IYKNWUlh0nvHciSnGoBx1KAbcUxGKvG19Ds2cV5ReSy0Ej9e9kDUQ+hwbBSAIMWWRqv1+IUWyLYS
SK3T2gU/6QTE1Bx2fOnlKy02274LY1W9ly2QtK5X3KOvOOJJCx06tJkpqgwtRfnI5apxn1maY9ph
VtXLuasHSOOnzYhxVhlFKlnLQvknRPpC90WIzg9K8Rr4p/byVRf4a1V22/w57C7Kl1Wgcp8rbTew
Km4ENZwjPXodkToCb4MQJ77W+8HjH7MbjYhHHS+NmmDq1VDh26xvQ8ps2iHOaRtEw+QbQphr46Ty
itFnbbd66xQlNjyg0w88iRqlf7NlvB5UG7QkiFcSBkZV7bxgF1CNWsc5DnqbsKGX3UiMBx4AfSld
X/FN7bOqADYfqlgXAYVi0lCCm8aZq8lCYzjyR08z6d/8fQmtYz4toozJt6uQhi4ButzatHzlC2pv
y7UTeBYR/DBE4c/5iiq42sbHS0ZvWNsXw1qicPtown4hgmvNB92zn8bMLP2raEi9tCAD0VtXGjXY
sfeE63AiCJKAuMJks6ugLt29r2vWqEBWujfEfW4iREZKBAdcL84oDPTQU6Zcmubp1OwRo8PHrzuR
llzSosFT7DFVMA6PFOAyYxY0NwtxfNoTJhJyYuLNWwTb6v5GappB0FCu+4KvsoyPwPsUtgsGCTzu
oNTb9XTzodRV5tHxoElotVm3WfHgMPGU1PdJGyX3J4Zr889GtrymyEkVwxTJLJJVkOWAou+iVwwq
+3cvtipu5zf3ozjomKphtGdnD+6dopWT17KmMMtd9RVzMIn+yfn0LhUgdsItIBFFsTl/Cf93csA5
W91hlAnpJlTICGNeQ0y+uhVCIzidCur0e4ul1WUDH+OV72zZSvNcs0eoLNk8kFHsFkZHa8vCnhbp
sFtvKb//IQGKBZLAFFi9oXzSfRJEOYaLQFs/5mFBrz5dVGZ4r0n8qktNqrovJBLTpfodH8d5Lpin
yjTQSgSWg1peoioQFCPxTXiPxuKkKn9YlVVeo4Ts8ByrFqHS15KO6Bg9zXjcitkDasbhAhA5Z3m2
lCXRZuZB3EsRTLqm4Oh5IHdOQaJ4ngGCf5SC9NobLzT1A1pWop47MP7zV1oCESPYGzCB+3oZvTKD
SUakx7KIfSi5Sb2e2nMGy7cFqXaN5g0C5AaeP3n3w27Rt/JzOO0nEi2oaWEWW59pLoJrmrAlkV+3
Znxu0w+Uo6DyhOkYQjx30IIrTfZsYKqYYlBDYiZGpe776Xy9FtunoFZOT8tYzm11oNOVUXgbuPUc
g7a4hiLI4yssG/bTR1nLqU9zDWA29SL43BSkxvlqQGYeoxAu8MkoAVfM+DfjjtI5mIAOOXeBe51v
UBC0uaaReLSzTJHX223p+hRtZIbaTsEubeLUhYgaOZXbMZC2+3U/LDxpKuVCePfAXzy5hcYEG109
fktzRN06zyiDNZdLzWXlD60ahsRucwf5rWtUbt7XHRceIk3mAnID7uPXYgCA+xvLyhOJZ+zC3MGf
1rYjoYYaLxrFpgvX/zKbP6SP5J0EXLOoVYwgs4EAdRlIdzTqJMPrkxDcd/RZQr5hpMAqy1DALOyr
O8M4xYRvOb+qc52oBKF0ejPcNgbLZDQfiHaxk/yfoZOfmA1pb7oSjnb/EZ10IVygs2UrZJW6A+V9
AR0YsqgxMyMkCRYjcwObPXvH7rXFgRHsMCG/qDbhS/LV/TpcotNa3I3DEjWgKn7Aa8yrGoy8E+dk
9MF1kKuNdxwXYet04N2htzdV8RJhdbNoiFVWCFGq/BfOzOVkF2/1662OT8/TKhqzQtt1692wuUT9
lYCC5TEcXAU0R+cBcYXg2SgAgwMdg7IHjkeMXwVGoE5jD6GJgLeODpIGT6rkDNZXxx6pnFuQBuUA
bK6pT5ETy5EQNCTXTXf2uRMzH+rRoejm1getQfW8Tb5Kq9EZ9yW2lLFa2OesAIOZ9yPbVVjMrOX+
zU+/E46dnCnTd77GhtbhGIe/dKQd2VXNmDxkuNi92GLteDQgslKlduSJbfRhpkQOC2hxfIG2HshU
ujwdxcwRIScd9jir/rRZlDi54QDAmex/hDixsW2Ov1t/A3mah8rDnRbzxuqmQV0ulZmWAyl7zqwz
uPQ1jowcSrxlJ2fbVM6NyXshbLIh61FJcJtCfowkFT6nYaWUIzVFyrWvN8xOPZi443D3ufZDwJnj
7hejuMgLyUTf3ax0mksEHXt34PBJrWhzVhfutzad63mXUxVXz0o6gp5wa+nx3Taxw+uRtzs67lz+
1sbF+Fa0WYJKz7VtUQX+IhVDuIPpw/RTNohc9MYutorY03xO6Gck2/Tw+6i0+36Rck9JKQqX8lPS
Nz/PJBHje8Dju8cVByN1nVt+KHSQmjncRt4ry1yvUmBqhb+FFwh+3WnVHfR3ZK6B6tvcOmiJUU/P
TkpWdHrCTx0Fh4zSz2mzoE2MMDaR96E/sn6u4tIWr78sux5oGitecmb9L82W4IfsnC11uhTjjMU0
29vZo+gW9mTt/9eC/lMQP/dzBpvpuNNBMo16A+lRdnuwbraxtovMCPjn4AzVoOXcLBWFkWN6Oxz+
RNiYcJkLvVf0lkzjFYjIPqosXZehJrG0nBs1I38R3UFzaltsZLWYPAoaVUdUrkBmkkXbJWxTeYKh
92rWpuWzKwdatywrVSQ4zwFChIDADkkL0aeV0XbD0gMmaeb/40l0jKrYolPs9P9j5KmndUkHfqvN
5nektBOf0dyTq61x5DRroW3j210cOeNRZpx6Ezk3hGG7LwhcSMDPjWpt4P9CYt0D71BDWI+s14ke
q6NamtL9lPVHtvPk3H+qFMFsgghl5Ecdog4z+pf91oqnMr81UEnw4vY9EJ+by/rihI2EOnOjErb3
Y5PTGw9Yxifgq3Vhw/cpoGNiGCFi8SMYH4CqiqTftcO5mR8BcpcqPc3ZM6vjw18dkyhfJ2bHKn+u
sBCnRmTAZGxpLSo4ZnoJbaWHb1UVjKwXxr4mWjMmcwB2iuq32lTfc9Dch7tRI03Mq+GanmjP0+xC
Y+7BKRtj6LA7fROXhApGAnKV+TkAjFDPKia/SFgKi9WVQvwyoSfdvw6IbuVgyr7Ka06XJqfSLcQg
MHVetyk8E+IVEvcQbF4Nq0UV5dhBpiy8BaWc/wK6MVG5sIZhE8jwelopgNoXwM4WQBMJuvwCrnQu
g+MPkxUEKn02HcJFjYBMb9aNR4nvkoSmKowKXoo/OenPWFuvJeR8YGNEZTdc7ZxfAWoBctwicWx3
zYMACqOeiClpY/pvs5fnnvEUTDu7k2OEBpz6sip2cHtT/OdaRdAkyLL+s9A0fBLsGbsdn8b0z579
te+6I6VKd4Y5y4TYCZGzgQfZnOtOsLTddazm5ZcLy0th3hpXFdjdNv04gRhEAjp3ZT0nfRZ9Xpbj
GFc0fOu6KpFFnfzWh0aKBn/Dp2L/yv9yghDTDbe8zRhFcYUXszJxaMOb0/nZ0qfWN7Kd15JpgKAv
aBr7L+qkwO17bGNqlLmJlPmR8h/3IPtIpEgdQSgh5ZgyOZBphfuOLVGxo52WUEYyrpXxTQxhkBK2
fOyKdtBHkCLFfz0gSSYsRt+Q9i5eWrlETiYsZY7y+nlMJsbnctfcdtDnEysVhFZGfavXpjrsc5wc
RAPP52118v3SuvETKKBa5VkL4ESInmJhyb0G524qfev6yNByPfpZdbJqJ0JOsuJck5Yaxx1YdkHf
BLqhZOJBl+JaKWR/7e4Nqq/AOT7AA1TzHCa2A56GkoUSx11c29FP1KpU+OgcuZYQ/2mq7FHNpeTR
c2icH4cd0PiFOjEwyXe9ejuA5MzicSkRk3Dssqadja8pAWlqNGzQIO+f6Vau22hL/2r3vJwEmn8W
h6NQcTEOeXPemp2KKjQIXVF7XPyrZxtlhKCQaunyXdnp2POF9TLywAKx/tDfTBbKhOQWm5TShXPj
uMowvkJSy0sn+V0QZpiVfYkME0B0W8nyB6ZeI6qygosgDYyGdPCrHLvKWNTAyavvm07i6xMixize
eQi9rF2oqRaNv7VEEcpLclujmDu+wcSYRKKPl1Tfpiw55BIVRKjLFCbK5dx6ArqOw0NN/n/5PnXu
Z91rGa24PtIJ1t/JTULzpEUhW4IGUMivpLyZ4vlLwQ97notJwE3aDL9tIHMsWB/swrQbTQtJtMOR
RLaSxUz0BJIug1XyRRyLeUPjCMfcRNupiP1ebNYyFJo7rPfTCjoVjKd+a7xECHjL6JIWy6d6Zrqt
P2BzPtpQCOFazV5P4V8czAq4UoFM7U9cNzhHOVIgh4ahSwqNiKWAIZz2Ym3BeZRDslpBAjrwHBkg
4W5v4VGhmuvAh3SY8aNL4r4oj1ROYI8Y3NHBHZ/qzMq6bM29z3YLRDp4s2PqaH+2k+BkQZXP6Uba
aNpqolY/KXWg4w1kPQ0lU9Sf4V+gmv3wseS+5Aqjw6WUqzMcU6ctDQoxmOzwMgVe7ZlNZ7ACi0xL
1wTFasQLS+cv+pQZ78HPqIiCbz96+hkYfgp/ezMVDzaNTTnA0QEbPnYYXJrnQfsXRSJRArYH1ta4
2OHmWWKDmXurUsaEkP8f88phpi3l8pY2Z9+GafNNwmeDEv5evz12HL0jxSDhyGBwGK5J1wjKxLC8
huqRr7DqVmNXMv3bANCSs57SO8HbS3oZt+lxG3xA6ZBkmBHurLyiIPgq/RmvHcOcm8lJTIpLvLkx
9jfzhqikSFhYzyhuQ8AvzoeIAMs8O7Edpq16uAwYiVXANwRTq3uzG3fZAxowcKHyxg+jGySI0Boe
uC6ueLnzsx6bEkiVt2SXNzutgi1a9KyZrmQqb2rjUv0PM8EpCkGk1CJv9J5JLC3XHywMNyuV8B3v
u0/e3Tc8DwP0BVDkQK+ZcT+tAhajKA7O/ly7MiYt//7fIbCj8ZehuCPY1dsiKn2WZB8WEy8c3Hir
vEcGez8z+zhp1orpoPdc5dx7rJIvv80hux7D4kWcpPbtL7RW24WnLClvp8DW8FAlqXLy0v4GGU9y
BHsmRqnDLOrLjdttHkJ6yWNIo0lo6pxVwWQi0uE0lnb/VK5UoZLB7Jsi90uG0gdsUExS2ScO6W9O
Ozi3kB7mCbO54+QO/rjh58nwAM32OJJZJ7lfhPnk0VfTxJL6DDP3gPNW7pZHt+qif2rsKshkZ9Ky
iGSlWnAnQu8ykb3jlvuX7pyqOwcvRfO3SaXt/fpruC4GTclHVbNY3102lsyYs0I/Y+Ubagc4lD6D
xAii+MTpAGoI35KrJ8gLNO3Q0Y3tqJ2QsmlSXmq4AuqIIQnU49t5ThyursMbgW1VCtYbSpfK9KpY
gjFfAxr9ivMTBx1nalRkRPnfzev7LZ7EPNWQSNGRG9MCueVCDq4i85xbqOYK3/NlQpThyBsm4oOx
ADLlLmTExF1qvLlwmLKMMA+CglV+vR3YdhIlWhMWbzvslx2JjOaDdhnT5bZY3uXmr/S2MvK/eY5S
7F1b5ZEAfYhcAhvTDH77Za4fulUUh5XX7jtgoj4yglB0BMwHd3KNdvTrlMF2QSklrjPyEDAQku5I
Ptzm4KduAEe6FK8TO9/hEyEDfEVkNPiNU9q88w6cK4u4hiWI0T9GPrYjLt88YJCh2M8VvjrQm9oy
3kxK22bFDtQ7u2CM+4QmCHXcimIcQph3ix2HOEVRb2mJpEO1J5RLisOr/i/VT2vN2FNtzc2QrdvT
LDVFLKLO63OzYdJxH/bYGvUUo1pYHhXVbZUqNMvvCswuDHLAXfTeo8wh5UZnFjjanCDYEtdgOOwR
Aru77TrCg98Vgz0XVQlYdDgJgyRNyaeKrohN2HC8svcoHRVOvr03d9fOc9rEAICHqSygmkly7bWx
XbhFP7FIjW+vw3+NrW72SSMbsEZlZ+MF3GmpJtT5/u9kuzfEBe3RD2BRZV9A3bsP5gXUdGd/CR8P
hgIx3hYcPNLiYSOuR38U93QSUoTgEH1afd8ObJh38Kk2hRcR4qcrheiO4K3pvppWy4VMpveEfwfB
1sQkVr6GAxgEP4Ji2TjNXi9tEQWUfjlqOggstLM13SRpzTIkSrAztk9X+jvNtFsipZzx2p33akMG
QChiKHA3ptEh/qfUIt/tzjbivoE8C2BRt1f+n/wdZt2jVdjvEAU2OWkn9mbNU9ESKjy8sao+cgOh
XwjDh0kFUeZblFamKFrgKRfqPR9QOE5t7/IAYKM9t4HDxYIsStKtqK1sRm60UIcH6LjlNC87dQNK
2m+ke++0ey0iFtIKWAR5KkW2ZxIL5XeMqYDvSuOiIvXpNSStDkHezurZL6iqrfTX+vLx6r0ZXJdx
pH086EPMEte0yJvk+1xX4QUQwkxMtrPmG6bovqbQTR6ETGlVlp+v7h1wMXuy6hFNwN8p0i7ksJfe
soIXVACGcfnpQGPYjRupzpDmXF3ToBoH0+DiykzPAMElQQNs/6jCICgEjRpy8RLiWipH3opTgQET
ICT9COahMkE/UfFHsTN0cJzGoId8skDuorRHa2wXCxv/eKrFmMqQbzvUJvoJSvmOU77uFBk0XZrc
DQ9hmdCPpu3uNa6PwiGb6Vh+BDvvrYZ11YJvn7PRG/K5bY5PWion1l0SgTv7juVBn5LFWSVMDa/g
ax8GsD9TSmn9iS31ViIhYwrw/393ZrH2fwMmQ1PYsCY1/QF9GWnjdtGTFuhCXYAD2+jGWnz6D9Ha
TVoIIAVJ78VKZUxAS7Y4r9No3KO33HeGbH140LkPflFF3molpI9D/4IOccNQRv9LsnPBfkhAG0c/
AERJRJhixBgsuWZ1UZsbt+LodrD9zixs4rrpf1ZjuhMG9QrjfXtWNDsg5R8muISMGXXfyRFOS0gW
lXKwgkzg2arVzM4xeY+ZPeGMaLULe5hoW8cwwRKgt9rP756ICfO2niYSLsRruLIrDe07grPh14vU
eNBfm7esCkCCZkzb8tKzP5Hpgj8DRK29JvVK4cF5ZL3qWBiOOaTw+s2i3hwUPh+fsPiCgZ/pEl4r
qu42uHH221iWhBCMDVW4ThMFeXZZATEWJZb4D2x4sBT8lxOA+YCn0JLt9UIpk1mQHDKbeT0PPj7s
fOUpJ08XxNtITIs0vPOIeTtNn2+egHFv9yUSSwL3SHdoEJzURWS/UTDpk10x2kso8oWDAE8EMb0I
Gmnk+6Ak9Isy94O1brvs9WXAmmMnb97pdxID50NTE4GoZJCdnISuPiIW6O0G8ubwhGBKt5ssajtW
jKHLXDlnReQ6sQKZneSg7ekkRKEHGp4hKsvrXXwkmriqOScBafRToBg2ObMH5XsdzTziRTyouvLH
xRdmCLYtv0t2WVfDaPi4LdnpzslbiohqMx1hJnUXRYKWXQygOds/TzNAbH0AIP3PoUZWmNcG20Oc
Y87I200nMmdg2zEHM7f87GHn0BeOYVBCJpO16dBS9/zNIrtj4VPBFNMTdCeEjj6dnXGwv0Ws7hCp
NcpFZG4CLXXW/1G9b1IhBKtfCXCvRaBeXUMXq/eprmkEZ/dpSWanLHVCGWPq4dEwqwgUqjADgIq9
yt2EkkRHKKF2WhZfis4iFRRG3roBhgwjj6mw4kFWb2837jPKsT7YiZEKZkbkun+MRGU1fkPonZwL
eHf5FE00o3n5nSvLZoQaQg96rZfAYLKkL4xxgysOhGGKj8b/UJ6O2cvmahEpeOdQ+Uky8hTIopMF
+u7opvpNgVXU+x9358n598WyCFZ867NCER8wH1wX5KgG51Lc4inK6DMbmYnSaRIrghOLm72ZfRz0
oOTkkEm1UtpOEPwTCoKkqXudgSuQNLyZeT7bJ5KPd1hU3JqqpWu64Knz9uStl4AIQRcdLLLpVJ43
9YkJoZz60wZNl6ilpKP1xsOOWPySRN+Idkf7NT8dM1od7v6AB7DPQd/onoPNQBQjP/rWKO9b8Bfc
93atwHF0xc5ZhmyVeQS2PbkAH9WxuxuatL531npVBLwyRNcVAZjEQGCL2rt2Zxfof9HO5WScNhwj
aJMNhRWO1jTeB5K16g5RrzPBy+eENPHYv/QaJIM4VD22Pnqw59MEqbjGd69+CF2MRZ6r4PG2Ly/R
+TzYId9nW1P+XwCTVdE/1+7P7rJiM87P17Zr38CAiG4ss/RfNN4Fu4xrlY6qjXDNXV74kG4/OeYr
fkkt75hjsbrzugyZ6sbB6ipXKe7ZrXsR9UwJy5q9i3q7HU5TNEO2eD1+eu01rZdpt0aWYQcRqxCd
171hEydzaY6Suaa+e1lTvhm+PrhYQXyoF5CobSMkFDWZQYjjx9ACAJu9kBGtpoyL5JaoBRlNmwKb
W6Si+Jfxmgo50AYHnHccM915NPHs8tRfZEWreYuMDrpiLugvFNNXgl1nSSDGFv1Nv+709VyPeObY
UzYWf6k6gleepJtSo8Y+y6+YVocNz72e59/WYJxCVmV4A7chQgLlyTO+FNZqnnHQDDu6e8QOxDYd
LcTxMRcnq9nb+kbphjbHfDiI52krn5+jbpZyJFiARVLF2PoR9eAgM9gAyli8W+mnMbz1RfzbT7et
IiyQmWHDedPqw45Pa6yooFg+sasPC3+TtmV8lNwpIMGavLIlr/bnRiVhSvUN2lreTxAoDMuJePWm
xeC73GU0lAPT0g5biU8jua6nX/pL/wU7xUzFCUVV9hFBCEFhWG5eUxatmsl+XjPOBKQ0eORPxCiA
Yc4KYLMGCwhowPVDQIop2D1+3fS69vMBx5eTo3wQQboKqRrjwuxUmvB6ZXeaTvqBTRLRMiY/enU0
WscM2MPDg0bUBVcyfZaSmoxQpjdSo1Hbq7iJl6rigIjOh3tRFGx5NKkjmfh5MMb9MAy70ctT/VgY
Pu9l6cZE/Ju+vmAS/L+fbBkWjyMomzIlP89sbGmbujnX116UdpU9aQA8LCyzRZKAnHwAF/C3EZaW
Z5K//C5X7WxjsbvMgDad+W2EU6xouSMPNBzfXGqlwxg5HsoswDHan+zQFu1rNkd4LyrgeU5e+2nb
XtbZHwVchwPDxu5C/ea24hrpPTaUU788lxLcOTh1/HxDdkPQxL/q6FKwSNeO0HCnA7Oj01SYVojB
nPWDTpXpT9ZYNmx8TKhmwmsy3KbWdYN5Hmz05+uYVPaiCzRDRKIUhH60pnIyxTW6+pHa/7DmKjJE
r+vHmlcY1wZQcyeNELhSaCAxZtB87JWBJiEHXGklTgVLJSQDzdMCgOCrRBr8fSKHWld8D8vRQ5Je
efKUoUc02I/SWA4+z7vlPX6/QmJ12+pCJ1xUHQ/gdBsw7KKflcueotH8bAxXtWsDoyCJD+fo3fi8
9JPfP5olVwKDPQbqLEArjzQ+ga2T+7lnF1tNXdsrjb3JLLRnAK1UFabArwbUEOUhum4AanQc76pF
OwpWK008Q8TGkbMghMXyYZQLNTx2MNDxkM9nxEcMwrWAdKcuRTjjTyG02FbWZNoi+0C7bOJwEJQq
A0X4zLUYC+A3qZj7nO8vIqsNDFPq7gWwGpsd4WsMxP0Sqc4JYrV/ZdzC6oX2azmdiX54qJC7AghD
Di6q6R6UJph++ZXH3iEGWZEPgQF6trHGIdlNTz2iOFZdj+/3e0WV8jt4UDbOPtNpFl5M7WyLE8SB
KVsEj92HDxHaEgjAqWh5qTGiE+ZAUn+iKzE8jw/5N4xO3sqeOUdJEvdIMO+yA1CClus2VH5cABzB
rw5EG2Q3BpTvFgDGDJsI7EjAjBjv57fBVC4VAnq5CaMDLUm2OBzPA+b3qangIBkEKj5KIH2MyWyB
Y/f4WSqNl9a6lgcUt2hiI3uge1yfNLLZUBpMKr5vH+sHC42W0iGzByuN57kl50oDuMuGgSOxvXiT
/I5+EqgdHGJ4cQ+esLG1t2crgxTr8cvSKkLevjHXik+bzCqMQOS0A9tzmkdMwoZ8LIlrCCgxmZIP
NdOBjaQBT8RFrkgTU9W6PW3uSRbKBbN8qoByR96RxHmN01EOMXChnjy3qQOJIaYPVeqQXFziJ+9n
ikftLpG+TwzqGtkrRlzEQu/FLTgy5g3Qtmrs/V2OaDkN4LW78tKIhsNvf69uB9fIq+uC6I4eKr+v
+6mSWjmXfXTWJSgP1qC9MWs7Y2dxpnLtdVm/js1NFK17PNkP7OJT15AJ6lwHmphAteZhba9vPt8f
m48XR3RQUGvPKVLk80adxnKTdU81R90tXSKVxBNl4WSV5SW4JxUAF6hNaZbKXcLzcBntSxBwGFhe
/TUDKKta5VdDGPf5ksI9+x8XoGoh0Z6FE+LIsWEjlAmanTVD2P68S/tXGGetCQc/g9Ob/RNnkMnA
DROPkW6qJFeyModK735cz3o8mJTdB7dF1I1RWjFoQYahYXVnbuuFDQmLba2A9PE2+Ek0BmjVqLOF
4mJ0MagQ8VxhfpoAYzr14xOghNFCct+ISitJ7vhmJ5m+Q10cD4IGlDawHxi8X4FotpN3ksBZW5Rs
fSrXqMkjTXqaMOqb+GqJGwDI9KxTFfVEisZOM8/gKJU+dAmXk4Werv4F2vN16xBI/mxpjQ1B9g4A
mbBs2KXgZ2qG4UTZC07MHLnxBwt3fKBNIegPvfCNPbWxilxIOYqe1BFfnBlE3HKHL8u7HkMduvPy
/tNKnaveAXL8Q/T273e1ccPzz4BD+oaU7BG8++dTUGKd07niN0Tm/NGQ0XwiU0j/VWRKSr3H/WAb
QXIpsci/ePz8Lt8OK7nA+DErNyiY/T+UiWAV0f7YmtHVHuA0lY9IHCRBODFDILAjqOcbwdJr2ed1
gb+9c8eAltsVl+agGfvB3fSFo/GpaN4qnoUhlw++W3P1vWsvjgli5T5rYQN6d8lRLIQk2xch6OrQ
Msok6idvGo/b3ytLPNLV8TEYfgBZ/Z2lV/6P1pMRxY5eDnMYZfGsTRZAgSbSOr5CL4qSgSu0qydD
RGe8m0W29P2kR/uALqncSeLbt2oIJbYJuJKD01dnrGrinNkpCcH1YCEABXR0VLyhq7LoGYF57gDy
zMOEHlx1GfOuucOAG6g7sH5d4IEpBhVk54OhrF1YNqSS4tfVm3Rg7VECT1mfPYSTwAiJAYLq37sm
wKLfhz5azzeTOXwOuzMF8MTnKPCjVDkFNpeQ2/BlrPXkGKDFCE4B8rsW9Am95ZrXzvj9ba29NimP
bVpun1Y+0xT4yXSTMYZzyBrpSWQiQsJ9azL2+F5cC+YOBOjEskKJKlzp/whk+SO0jT70zvIj9lVw
wK1Idmr1JNHrOLy5sKREnsHO8KIly2Dn+MQMtHuT9jOGqc6OGz2+4ElsEGqHq5V5KtPo19UUg76g
oRglyy0y8GoWdLuoGM8GV7/4lT+A2lqXO+isg8LpG9oi+QCFZEOoOiBxvGbp2fS+IivC1IJka+TJ
yidoN5IYd1v073O31qmNXY4VVQjFuECBWkjEVTA+TD7ybxZ4M9ezbLI7mNdgS9c9xcnl9DVxw+uV
Taxp7ScclPzHakfkWLv/iXJ73kYLBH+cqFRARMP34EJDaZd3D5nOuUBgmYlVe6vfU0br5TQzQThe
3R4K0S8KK0hE9WHXtxw4ajdy0LDaoPmvqFcT8P6SKGjMOJcBcwmMkk8PCKahAigOgtz/JCE17bxU
3KdQJFOhhrCF1xDAKhcdj4lRJ1BVnqBZFvOG3ent0uuVI4gyXuJMK9bNDsRbc9hjuo288vyNJyfJ
VAEd7V/4zh/B0S1jMEOM6b2pXlMejuGQAGK1OjxsxsLOls8SjtU9Wgk2w/1Eb/Bbn0hEKL/16WGo
5dRA7MKGsXeTr82nxpgqA0+dXsaZZP/1FwJfzVUdifnxSuGWbTAtRt3ZCbnqVPWL+35AEHXqcvtK
7Hnu1Q13QLnEjKLIzuFzE25gyGQ/c5O27ySdw+xfNJTo23ujr9bA3slYvlrABoBdieO8x0j+BEoi
5jZM+Q0dnPq8O/SGkEDlySdL5IVLp1Q71fvN9GdWVerjDNrjm10DA3h9wdAf1kRviSz1jXi8Y3xV
fFHblZ/PDjl5Ijp0NVfn/QiYPvpabWhjHn7CXMnC5Qr72pztd+4Yi4h1y1/yDuBXhPbc/RTBdk93
ktfCrD53QnwMafjfZw0yqFEuhtml9jQG1edTio1ZLfar44vCDZZqbKRU6sLinN7ehcFtI5UDKhur
aeCIzzAxEGOIon9tdtTQAzIQy6bJ7rxW7AifgLYeU2w48devXlpy1cAqrXEJZjJ4HjhOrvgZNxVp
GsoU0/9jxB9NWr37zMc8nitGUFAf4NMfagCyxNwUkaYiyHI8mlK6cBxAvwV3fYgHjwia/XS6uEqt
sbu6SLYBV0/sd0A/q9NNky5FqiBWXH/9W9UNAlIbxEy70WuSwloJ7XTjRAFAZCsFi7qCfQ4N7puJ
okXhMXejVOKm8yW3iWAtmwTw66OHauUidogn1Dre9JLUwYwr1s4shReUJnYi4Ci7ppXZwiwGq0fn
r7yPC3F46RbNEm1GwCWsZq28WgCkHtevXb2vb/7nAJLxfmw1PLegIWsegkE5MQsg9RHUw48+bNfO
QTgO+OUstfJcsOJREVZrdxuCc5rCgmbCs7jcKILM2E20gclnoVOBmwJS8HZFJmtEt8ENCJrPDONY
svrIbJ7gcgNIjmclrXMoq9wTJhbdSIYlbaMPBAZ9I6KkCAzTZyWXkAndxgMY4QIBMIuFsv59Qq8t
In5wHD5qFFlKne4Ia3Zb1joW/UDAKin5tuvPlzOrOZBquT8iV6/UO6S93IY/J9CMusZqQNiX72Qr
/Se1EYw1fhbpoQDxeYXwmqOeLHv21cWDJMKncPlxlX0iFn2E+KStLjRBA60HvahQ26POyD1s9Xaz
Po+K2/j9iG9ZKFulWo77PTIZ5JGtZjtzI4GsEYqnRYwrrK0tL1td7DqiIBKnNkB744OssR2h/uQp
nV8t9cY5HuB5xK7HAhFPYgXR9hDX5YMdUAxFQoXpyGtiIu/WpruxkO97l4hX6Pt+DWQfmZ+jlv3p
OfCOppEujPrdyxkA+lNJsnpC5AhcwHeXJwDZYO1v8RkdXD9IUh8OlwO7bmN0AMGi0KhKKfrZyq4l
rFaqiQgN9aDhq9ennFAQJ0u4DfSl34LzqaXMLwCwViaVhO/tqHxal7sMSS54MIHX34OKoRsrGQel
GzYvqFhXz9Ww56A5q8WLI+kJmuXrN2sqNIhgbppBUMv0qWG0RC9IGoXsOUMTY6HsWR2dd78380CV
ilwiKqXe5wkUP15vblMqSEAhwflJMc2GmKCWwehCmluhlj4Y+u39oIOCojt/J6q7IxZOp+VfXfKK
HH4tYF0dcq368C8DgGoz8wd3XO7/7W/JMnJybvTt42UEsQqxiiDiLpanKfeO5fEgDbnUIblzLcr9
WPXoHo3m1xQ1NUawgWBJukEvp8EquzFxqZojV5o23Gm4isoTE6mASWu+JfBMtUWoxSOd7hCoORYC
OoXmtPZ4A8ZHQP2KGOsUtGQT9Qxg0SpP14wAYASZv0ETPrDLhCoisofLuInKd4FhY5i9+/9pwgxR
5t6wf1fLAiAjkvExbuSNE/tJ0ijZb8DqDhSOSqw5ZMdRqScs/BDKc+X1gxbLimRavGCpkqFLfrMU
RZBaeeLIWsx7ztnEge66mdyBNLxAvISvWzb65V8s+DCWE8fI2CR6tKFrZgWw4monU7d068SH0H1k
5GIsJj8hZLg8T1PBFB1R57UQnj3qerEEox3s1EOJYM7+H2qIuZHcK0Mk72zm36omu6hPiKwWhJjO
a3EvQOMeUuION74lIvfC6RVtF9EX22UGsu15+0ZWJvBvDAA0NHlRzR84H4KyNbmunQosq7ne8L2F
O7e21lHPaF4sVoa2LIyzwa8b4tYN6bDK1itcA8EUpFpxSX3n5K1uVjaJsg+zGKLY2SKBZOUsakPS
aYCfS8A07WbSBoWNIKEYzo3lGSY4WqQpqb4tRYqNJLNG1pVOHKG1f4zy5EL6T53zMYjPZpx5V4PL
iTebxLl2KIOwI0+yN08ANRONqTpk1pV6HZASPV+0y7MskS71oTKxNRoD2dCb3w21W7AEWhPVMX6z
KDnCDKvv5e16oo2Q0Vv5Lpt7BELn85C2D+c8K+ZSc/Kj4a+zfXipe/AUkYk6MwNy3WB44I6E7uPK
lU1hKIuz1x7si3DYfPuYckS518zy89xOZspYVJbaZ+Bav+w4wQE766iJbnODXUGE2k4PS3dqQFL0
kkZ445WgGyOPCe0K15Q5vsGimAgtYNBwGt46h2g0QyneO+SWDTia6DNP2yW0HNFgrR+dHYQrTs6u
DS9EmNLh/RHoMAt+6Xzg4NlI2ORw6RgCiQGabHmXbJWxMgJBkKv1+QDVmpAJDxr9ojdr6bLJOAIA
5eti1vhftfW621Mcft4/mEHFz6Ix+dEI4VucS3j8vgYVfaA/73Kz+EMKbR+k1GFUlUKOmL+a461J
fZW4nk6/or+DTThtdtKpyq1IzgNKFjIno1+wd5FfSUHm4dV1jiuIGcGRp+wbDR8DO+Tm2Okr0b4r
LJ5fZvvnkWpltkjfOUOztbtTVrAe0IIQH5Cd06OhDj3QXjscrxsnkFyo5ndn6GnOjWoXON3Zq03b
4gJ7IcwFXqJVdjD/9C1o4190oEQ2lk8rvz3Cb9v37/duouxUiZAV7Eg2BOyCJ7kkLOupF+vTTmuq
fzGbMhSjOHuBR1Bpg3pX9V7NuS8Df128R/beJ6tL6uS5tnQnaL1dbeaU5mvPcLv89zWPeYrKJ7KX
Bl38KzxE48qg7we5FPIqzACYeVH0Z+H6FuV/4sCYsM/i5JQz8Fi6MIyXAqFWQsGD8INXdNrz5CFp
gDhG1BgTwn9X5TZ4xEruj+a1yEny/Ylh+1yuxKzxQPh8ec4X7C6Mh5B/PlDVpXXfQlxpRj4hvxqS
Zv0fisNM4Zwr7/7jU9HL6SkdejCMyg8v8uaC7X408WbTK2FdpLlzujY2Hk8ZmRLol51uUoov1fek
Mn8RORg3uSoih8zefbRaWd9lEfSamZpAVT1yQ3OKsGselaZF/HSsgIkswXo4pwlfyE0SKhxl71gd
JGCehUnk7vh1dDvs4xmtYzGbKvABtZj5IW/v092Ah8aQ6oIejlc0TNdpPhqbmmoxgEkTRNijqZEy
NDkBb5QACXlyEGH0AeeQi0OKLXRKKhbNOQfPXaQF32yoTIQbhiwhasiL41k4Cdt4FRYOHDHcdC3M
cSOoTzXzCTIf76rxPlAX282VQa3SkaZ96FeMkJloU+TieozlRCcE39G39KpP49eYreOtEg1J4eOR
vgnHhQfxIdNsqH4JUnYD7o6V25/0aDf0C8OZMkrNWfaW54l9eM3GB2j1gWTTkqvV+G2FtftTDt5Z
9/9FrFtROV6V2HXRyQqJhI4zgh+89a8kP4ag8jdKIhqr6JKrVgGzfvIH0C4zsMatWSqgf7soLGm3
zVIjppZgV/JjxqrqsI7bHPH80cnHCnJm1abngS7V0H5PSvZ1U7EBXFDzQX4HzqdRLlGx+7M1R0dx
3azZ4NQuNFtlfTtiy1xhgyKO3i9/4pvgPVm48f9GTHn08h5BOwKwzoyHCKcmZsCrPHoUWEw8Z5nU
eQ2nARptHgdhsedTna3zHe9VxTvhiq27pa5KLJc3tdnWtrT5mQi66nYPgKxCJa52GL1iT8S4pYrK
BOuDmqn7GtQ29CYBzJ+e5Ndd/lmtB4UDE+XpDldCxsBJ3eD3HnsWh7i5e/+70ZI57xA6GKhh8A4O
Y5L9bahPYfAyOoKI0MzcWozE2EElohGbk3ddVwGXTodKkIXDdp244toJESs+sTJKGns1ZonFV1gK
HUbJs2ISfVlkoX+TVKFkcV3ZPEXqqvxrieajD9lHRebawjXIlY2EBLzKL3+gKPKlCgBcEwcKTLmm
xTGzI3KehqBGhYcJTYO8cKqrIKviTzARU3LyZ58/FvRsg1ptQYquBzV8kTooudSa/EOal9d3jGVU
tRf0W0cU0ZUsx53mfMJimXD5WslDWA8SzGwS4EQ816TpAHq2jipko7vC7MYp3ZZTyV89roYTrHAG
WY6dmmHq9/TJMLuAz/0O/mOyvZAIqKv88EeDPr7MubnzvQdFn6rjy7z8YKhD2yR1VG7OQ4SIP4wr
1pRTvrJNaGA9dfg3gNRvx2xWOI2JNtUxF3B5g57zeL8XZHQXzmTdNBxhkDEs4rbhLniDcHXrFoxJ
cWk7CwS2rSAvaRmXEzajUlJUQ3CRMRPapySODZWooYttdek6PKl9mTOdnwT5qCN1XcByamPkMPvI
Ay5EcrtXiu5KxKbOp8utGWDODBJ2BZH5KhARWkl0wdbXSVsKd0cL62odPYkU7HNbSH0Mfh7Qh9i8
BXLlc6E8MvPMyeEZ+a2aqtOIKH0RinKXD+qKwfqaPUwCtzeU1WlKo4+6Kz/iJRVjMiynrHLtt/nL
k2LAFdyaOovxhl8IN4zxOioK6EBaFvcv2rSZPkW0HvzhwwNTfVTTNFhS/c6s1jy4RVv5EgZgBuWP
FrGZ1fTf4N676sy5xAVBh2gJwcWEe4pYxMP4O/qeUF95bBjnH+tNcvIlcQSYmqFTwCiqOckblnM7
oxkNxsSuXLZufu3+jAF8diCbc7UrqKvfVE2Yjn9FewFYjAT/0xmKXtEmgfdlmb0JtVUiEkxjlSg9
3dh8sQMIdh1C5nOy+A1XFUO9ac5vmtMLGJuw3E7TNarRJscGA9ybmmrlEnrYrjpCgcK2WwcJP2uD
IkObnPdLyc31ApYj7wGXVO2FRg8VoMWeUvlgf3v0nDfwXUuqCxx2UKGN6fSj5e5OBEVyg0gC2obu
8iDv01qXuf3Eox9hnXCowOIweCN9i53qV0ln0QTCRpuQxmh9yhtJMj2NAIs6uQzmz/mi4kra3vlK
1y4ZeHmCs9TX+zBo5IcJ1DFBdeZPOBBKWNIN6TKKnJsr3JO4JYStqoyPivLYWRmgnl6oyD1gH/69
XpW8y1mA3VxyllzWdARLA6C6/ysjz9J4z+JdH1T+yLQ3JT2C0rlSz4i0Lx3ZcQBrcJ6O/Y0lJm23
5lHMpXbptkJLCTo1PKGzURn/tA1C1PMpQmRJU7nn5rNYJnm80dEHSInHDOTiF2kMcaf5PY9vJewl
0EOb2R9U2fJnIMi/Kb+yX0gvdTE5xVqWZjEfrQ6bXbe9FjTsxQcG0D/rFlrcW+aHm8hXn9jvNji9
VCZWKfjuE/37yC3qUVYgdTNqLvWbEhCCGjFSvI4LjqjBBdu6rfWS4IGmWwUV2t3o6evxYN7Tal6j
666xqKztt7HoFutgaR1GJ2jKhbJ2gZVj4AapcUAvm6qhvxzsPZF5mShd3xKrT1YU3VNSBicTty0Q
G0jpHLX0PinXs04yceVrp9zHL7K0IVbf5g5T+FiKP3fD/EKioscGLLaEFSjwrxh1v7+vsXxnu6RC
eQn7zVd9F+FSBAGsZ1cGBS2DnZL/TY1i2d5fPAMZGdrzeGa6dS8n7Vp32m59qWVAGtzH2iRhW4n6
DCWy8fAxz6G7C9At6Y5m3ZMJv0jmBC7be4TB4wyrZezZ2F9s+Zd2Y6EA1WHWJpS0LpytaIkTL5HA
Lub8iYan70yXXMxliVs1H7O/u3o9o4XG8+AanxiEN9fVNb9xBbMFetZQ6grKi5g4R8pOUMAsPgjM
tnjIOYgVa57QCUTsgWXErLfUHenbrcN/DOL1aMua91qGuLkxQiC6svqMTAp/g0yMfZ/5vOrHHo9n
DnJf/EafMTCPY1E1EK+T2AyG/S6qdBcGS94YkNE6cJyGk+kFpElDBFz5bO9cZAz96aEjus+CEk5Y
qWalCTAr8I+u/OX0TI7JcuqI916AlcDnwbTh2CcBQQWHlyzsVx/zde1VTo3R6AhQKWp88pNlaWc+
4u6IKXyPPeJBQKwk82hVKNZZELQhjrAh50fgfMnygMlmxBuowCXUEyrrR1vjcgZIqmxKAHtn4Co1
hiSj2pfIowz6rWSwsqIjD+DZJdCR3lfqBhvIr3iIg5LZ8LmM7z0BxyjF5egZ4JwiOyAYQz2m7nI4
sVb1LaQrhklfySGBEQChNMWGLgQhGlQuC6q6azm91MYewfF2R0PaosMcoS0770NzkkBSAF1mofAg
capV6qEUYllZEzljBjla3r6SREqFR+IaTvtVKQ1e7yLgP7r+UpPA/ZpOiYAb1ZsQL6k+nsYz/uqR
7ieC9Kg1iT1QibKl+p9ZTlxK/7okgFsD7VdH6zd5nha6AP6RuJTwpjR2SIXhhXSuB6ar31UOWth3
/zRV56ZqcjMZahECHqSghQ9CzyOOTtdmAmN7Jkaho5XSQ6qFUxlg+eTcBIcF4/Qayl5g2BHJxdPJ
LP2WwCpKrS+nA5vwiz1At3tUsnLW+2hvTxX1vbAONdB/UIzJdj7aOE8/PAvoMkjfn+ZnMKMdzFVr
uLeKCtIAAwrp3NRrwZ57e6pMvam3GcyAhYY6y9Dnhin97PKFXHXNQIOeblFODwycrzugphera8WR
gYeRB5eokHQ7UJppK160XwAJvL7DTOYiNcINzgOuGf+u/sGfpGFsZ46GRS99is/eLAqfO8RXZCdb
vhuJ6VBCSXjvh1k2KBP3X7a9qR5l3XqG7zbeL5yMOBxm3gacEw3BoObW5o6z4vkSH40Xgxa7A9xx
wCjnUqgBzjPXbbhL642Iio0Dh+28MbhiBeT5PjBWZsXVggdDSgVhV0STcTYIhu901WrvmKai3iuS
Zb26fKpJIs72CDQab+JCvY0KF5bRYLHvTFj5uBv9q+z1EsmFIzWKwc8pLOcM28gcmVGctJWjXWSj
6mfXKn7j0Gx5SvWvkNqu9UYXVB3OE/+uDjkrC3Wi8hZCKKI4W714x+XOJlxKpyI9EuEDz24ihd0D
QmSVP2Esbde8Tbd2FohRFA8/f6e4g14zCsDcwTltFHZYx9JW3SQiELNsbo2S/JgbumsCbHJtezIf
/HEAtHEn2DlzyEP97k2317YIrbkvJE5x3tVwDFBrQC9zkO/m6fDSJaKzcqMchLej7AIkWSxNm6IE
XkZHPfMKdvx+K9rvK/6/bxmzDt2IhqEZY8nhr66upovO2YBZelcg9+5mALS8Wkjup5por0WTnlVD
eCgqLjhsmUrZFJPYJrV+HWPV7b7tS5jNgB+gkHINIRPE0WdkH4J7MFIbRxALu2gWNY/04pAXE0dW
zcmD0ZZ0y+LThYkVqyYkpJayL9PbqZXCgRehIfKkPOf6KkTG4fK6hT/YjqMIInvmSlO11XLv1b77
3vsopSZ6+SwLnLOKXFQBiCW9svtjUqglSkBb7flCP70121cOS5y/6kbLRey/rC1HdsHKHUaO95Lh
bMnsMAKPK8yvi9yztpFpzEgJeRnoSOey2jiSz8Gtr6M/XYxX8F253ixNEPIbdfQZrk8nNuC1xCqq
ferkb3vuwT3/WOXz4KkxPW/TzpZ7WRwlXH/OS5yf/eCgqNLNfvJuVjhZwa7x+/w6mZQNzlIavCgV
y4KAwBTTPKWifrYqbW/1ZMDbl+SP3ure4PRUOIpoNQR/xmhcvkq3pOY6hyUaNrNAAkAX1uVwrjLg
9AYLTZjFRQon9xhYnAEhkSVcTWJ882FawcHHsoohZh2zSn2kLPowHaiDihwRBUQWyXbU9QX6dPSE
piKv6sD3hEdgqB4H15zTb+PJ+22kDh5Ez2xfISw8DRuR8fg4QvRJaGbjfpH3qb0xytRl4jt6x3sr
U+Om7rDRo0Id9J6rjsRJIxO9icRmwiRQFWIJDz61GcQvndgZ6rfVFtLsPCjPx4lqdhMpvIqCpgPG
QpAIZW+fg7pEUNvL7XnZ0yQZ5smuOygXTF8d/2MxKsRzDKJMpH3SS/Ij/I3P4RnO2bpnpeE7aT9N
XdL3SkJQMw3ikkx27CSfiRKvS6emvoQEL+l5F2U0URobpzZ2dFgnTlvnsBdN0vwm3ZookU/ESzZO
W5XDvHK1B7pkyvpX27qRQCTAKE53Y2kq2/XBn4nb9ed8BLjszEDWI2p1dPMxvN451IfpQQRzck9D
MGKNzPcO27Qe6EBKb+uxhk7hNwkJwifGVIbafxL/0Tzc7vzJwSdwVB/eE2Ybps339GqrXsYUXMuc
4oShuIlAfpmY8beVXMF5p7fDtjWvcSiEBaoUqztwy34cVgnbJ54SEm6NVAOmEz/CuyYyvZRqqESu
W2HYhcSsuN0MSxhiSSyQS1ZFru/76e/yzv0fQZxkHOvUTfiZKdLzH3zhqUPw6ocPlYBiO5Y29LB4
zUfdBn4eXt8jzh7Xi1GD9d5R71N9kwLUoT4zUihnWjHyPJ0xQMYDyllbGvxnQlpP0Sqea5Ko2hr2
TdTqz3O2Cyacdvl4JSHaiWsdlwhcP0nGx3BVdExqpavLk052S4eNrx05JBSOdiXFVziENLkGTCTn
pEkF/CDwaJBtgathBuJQn74xF78qbZ/K1ZCRTPHGd2l5Wi1Ud759rtOGg24oQRH9koPjMCbcd1rN
bZD5hAUk9yhOOJDsItO42XitQTKCf0qHfOKn7sHzBTikfZc1JZuCIHsbf+wOwat0ivWImPLu+03X
+tXsq8oqQeKytYw2oyqlrMIaXGKRt8vl/g26IfaJJOeZSREXX5eeQGYnbe4ej0Nssv6wKhQhdTbu
nNk6vM0FOaDh0/bTSLdjxfb+bB7sGY8gBJ+a9cHgZoC/Oq+S5bArsMgFqdIQ2NxlmSQPWwM75JS/
rxZnqx+H/DwyipcQuL/kxjoWrskOgH7wwrzPs5iEVekV8GV8vdn/cK/SWPm7MzjSBMOANRAmpa/m
h7VE1itP/sFb4WtjlRO8zxE+GCIpA733xgHypMgkuJBKlwwJhxcfzBnWrEztfuF3A3T88G8ncfly
iG+5IOi36SbefK3syiuA1U5hFh/hHp3r85+mGKqcGqjG0bFW8u3TCFNYKly+ivOtLS4dyYnuCT+b
z2uZvtt+dcQeyd1SdIm6xguTb6/C9hM3pj0r2xkRD+jkVpqmn6pfMxvj69sXIrf90JtIIKUfDXt8
ar3QDefGOZMjzM9UtHIQVg8Ypv8fz/32/S6bshO9JDjTPxa9uF0Xx5A3Jr21s3Qs34ltdOnUmbo4
ZSD0XIWN0WQ5gaKkioWm/tlkuqEVedsa7des5X9jzC9pz+S+JFiI0nrzcl9rgCPMV5cMVpeDFC2V
e7YqEyFJVGF338PlODUrR/AwUal3TzPgsKoHSodfsoX2OGsYMMpy4Il/28dtHCHuzfyxIgmBDgXF
TARYZ0IICwlV1FcA+XRy8MOY/3QCJrrwYG8/P7qXOrmUJ7DyNukcx+g2PxTkpHFnROYQyG+gvRlJ
GsmYOfysr1VUFpnvLb/FrX8GRbrpB7rP2GalSHn1GTjQRb+y6t/rW3A5YwsKkN2dvFw0vx+kaKu8
5wsFeLVnerE6QQcsxDu+x1roU0FV8mg8Yy8wkDDTy4pL2pthf3GphanBkS3EeHhkr4Ewt/PV4YxL
Me9YZsuYeQ9HIrrzmyVBzaueHg2BAXfK1nif7zsAp1B//1JLp+AHs9CQD/jsLtOAuCbbMrwW3TUf
13qHR9sRGruZhL4wyR0Sy31xsbD+3G/2ECtq2MP69PC/H5hBsfWQaozi70sW+UCB4RDe35UaoGpr
DqF8anJwmiWhA6H8ll3x4bqR/GHE+hXEv2lh7CtXKQGxqPVQBsnfZKQd1QmzdH9sKq87ZHipklV1
QmeK2xDOKbseSP0w+xPwszduJu/ky/PKR16D6vMJmASem08r45J8RXIVwyfS7/izTvFJdirbIbB+
+Uaw2uq3eyusXKKQSYl8Wzl5P6UCGZLrAEuj6L2+n5bRMiuWtqRvEvbs2xzpv+6MNMp554pAhb5C
MasWtYNTiUPZz1Ai7c3P9lg2VtGG1/beIrM5xQ95DfMMJvn863xlEycs6v98bxGTY5aBp8/K/nFl
pCPpR7frkdljk6TRi6MGa9ChCTXpkyY0N0ar8OHQfWQ/jg77Yf+ilhcjSw/5Ka3kknVB4dBWLSlZ
gtrFGnxeVVjL8vhs+xxSNfN+ApceD4HTF6k08+aGB15fIOCpUczH9ELrGNMmYFnt9tvvO8mcZyIg
Ugjka7iBs81108SFIHnC0Rh1XJiPbpt9yJxX+sphXmtFTT4XBdh2LtYdTbzXkCsojo+QTR9FuDOk
dlS18FBw9EAW5zxVKPxlg976kzaX9iOhwaZJFgLKUiOvmhkkZDmYJsj8o+CpsSFsun4Xyj+oSMb7
CnxN1IhNmfW4v+46RVgBzO+PN7zl9dAkFp2WPMKT3fCK626wbsjINfEEpsjK+Xqr60ZT1SRiXnC7
3UnoUIFLjBAlr/S4ChVxyKsvZU7onnS4ZXrecRzt4xp9woM7+oZQyj6wks0sE4IQrgNp4eHN+u+p
OzeOhPb6yU7f8sbH7FM97tA6/H4YW+OZqIFCv2DCCrtN+GddIySK8pa7upo63mbZifStOF8LIrO0
8GlfPlmmxIvReQCfRM/QASdtrLdZwrSM6q2620XfYPSJ8NcTkHq6qOkSeEg05OPARDox9vrtuEau
7Se69POD8ks07IP0dC7szim+axYcOsvk668i36rd4eJb/AV0at4pYNstwUy0QgzcqSMjUGpwPavj
e1DXO8LG1LbqE9lJVBBh9DSbsYQd4QIvOknRVY9KDWtWUTzdr2TOcAHAMfg3rJ6lCRjFQV0zQwbX
5Ejv12xQIUcuRgY+1Iouvc1loglHhwpwHuYaAwh1gOBNIi3UGgfXVCcSjV2yeaMZeDrJCqpui5jA
dsA2ntyMV6nxee22va1cBgNAGy6/VlRHAYxnMd3a6QXJA780MKY5a4m204SM15dLPHNPZwoFrQ+S
/AeHz4yEB5LtigkSTuQa03sfce/eyD/daCtSPe3lQ92f10nG5yWa0C7Fwp1uSUWpoUcoF3n1rC70
YePUtDGySvNXUZJ2sTG4ZTyged9nKx8eOvo8UDvwbzTs0qVvuDgGDP4NdBy3HhjrqUiuM0Zs7pjf
MwVqgO/Dol8w5ferU9mTnc2EdeDv4VW0sHI1cUsdWBT9YILmzxfeLgeYjxkXDfyzr+q6Ia1R5dPI
6LjsPhfGaJ9sePYE1ZYtInZkjaqGz2V+wYMV9hLKZyH+GMCyWGtYpvnRLILiwrnJRcMiUgjad7R3
6yfswh5XFeSdlAVGAeRiNGKuf1/kHv47BjfPeml90jrepTSl8R6PhTMlIm0txhpX7epZQIvgsC3H
TUoHtC38W8qZiM4xlmkFB6dEOh3gIRgqnYG5HuVsrUuBh/gxDjfDVL/q8SyVHqtyFZTDgnLDGC6g
jCnO22/0MJPx1SZ9+A2UYHhUAUg3gUKtsw0brsW0nu6qooxam0QYdR2lnk8BbiPdfT1iZRyaXyHL
GahKaquR5g5kCqIsVzHUZkRMNr6wDqB10CKuqsIcNjbmRRIKtFm7taZlzDyF6K6lPh1O0Uyk9RST
FF4ZrBCaDhUHr36p6Lw4qVgI59f+CEILRc0m2iKSKTD0jxcZeya7y7PPVuHuEPCW3PAirgrnlZHp
dpisDRLdEPriGIdvhhP+kumKQgxzDLmIuEoZlWa5fL/FQV4BQ8b/A2FE2HBw/42zHnQT2T89SY4t
CllTobsnUXpkl2b06DH0kfumE/8b+VLc9XGrRcm9q1LzqC1se/4CZMHHLxegP0Ge5qwdG2RK8d30
71z0x4RaQSXdtRVZ7oCiZZUHA1UuJVyYeh1zZVixzJflcuVmyp37xQvS14pG74v7TK9TiFYLPVBU
JsSRqTBH773tp/4lfoZ2DCSbiEk11uzMRQx0fG+vRmINpijto4UNTl31qttiIXe8ps+XiViYGJJq
o4iKHyCkwvnabuytAg0jgf0nkUS8bebTnb5vPIXrDtXlipBRQ42vOBKwDQdzliCpL0HSXMOWCcRn
VEJfLFAWjUxbV0/e2WCUPVebkOmfd8/uuQaugcvIfGT1Ajb51pnAa1O6WE5CO0UovvCASOSGfV15
ubjQa4nvZhHPgV+JiYHlUzFsygB4q/YgP/TcfOt4oIo/T+Wug4hb+ViiBluXjpfcaAKSREhjuU7s
hgaTPZlM74ZzmhcqDdSUZhWQgkvTs57zkYWC5bAF3oDYh3sqe5AXU9hMwuL43vxCVFQIzPmdovX7
2Q9d2364qXo17tdmT5nv6eI0MApcVFQXmdnbs6yEk2tYPD+hQeX6Pv76Qm0uY7m1NnCM3rJ9KhNR
09xxsTq1OidVNhEIA0rQgkFXLPMgzLDN2Jy54Dyt4oVAPk8M0dY8XD7CpB6fAIg9F3gZB/c/vpBd
w6glliCcOdhM+1Ca8hGfDSwqoC3sf7wFR/lJKpOs3Sle0uLYABcxiWEN4UnjYySPDPmNQ/+2TtMm
szTTEhNKr5lcDrDr6qG4+5+3Q/GtY0/FC8vsDnyrKPfOX3xau63s2sQvM7SRCSDBbWAKUAmEElOf
bWSaxvwJ/J3QCaPMB+2T4nrQt6U6FxyF+bZaGzqAcIPTHCRSE15235NY8nkQvaZWeIGrxy55yUFR
kPr9QZGmXeMKI89dEbCbVyNjQyNIPrS03gXo69Ppk8GYFf1qW7+YiyuB8x0YZrgegtwUJupqA1/a
9VdrUwTMFk0FN/co8nGrmh+Zfv14LG5htOZYF937SS8uyYYok3QJpaaB8tuVHuzgkx0bIVBNtf/z
HXcOa2spCQ7fqUvlZMuWFIyezjY/qzWrtKzGcYFMVSK7TNQJtYNemikmmpwmO+SeXHiAxiZ8g70/
gJM+dl9FxVGoW+hLf/R5Su3ib4YNhQggU95I12ck+Ty++T2ggnwlvLy3sUi3xBgiFNfj864xMkv0
Ru2tBnPFWG4XqoIxd4D2vSPEGsmvgWpKQPtBAjoEGH5G/vBqluJjx97r/rLSDGtLpGfHV5qjDdEM
HaCHfxs+liPeYguACcgE6BjbWJFuBIsH/YBVhYYi+b1E4b8YtCj7yeKBy+escnzcHMbCl7tw9kp2
SIiQzTVDozxqb6DYLZL4GASevRQNKNbq7BbbxMBJ5htnhChPBso3BQcx2OTRHGF/iGzmlTcsewEe
1SFJxettzy+Huzf2wFytGwn19+y23u6UfuG7T1RSoa8lcYToe32BWUD9S1qAV/BfGMhtrzE3tivA
HQqoOxkZVrYZrQizGkqWFhIT+Lfc9kXkEqk2qnD4k/HHsZPyChy/3MyglRn7x+1usboxmOf+U+qv
xSZTYQZmKfPvjjViDjVA6ViI79yLxPRvFcrD/5krSa4EZ+NU4iKaT8jy5l3JCvKaTEPv6O4faTrW
DQ+1ZP3DdJWuh8d6QFS+3xesQl9XtNyvzibANE/d7PlhHWb+uuqhqoro2rNbEkINx5UIQ+XQgm/m
WS4tWPHVmWC+dhEV8Uas3xgv0bQSwo4vc500N/MLAxFS0Hqe+xeXoI6dHMy6PtkyaxA+cfRf+xvL
agcuPuHGpVZRJ/x3FAtFnUNCGbmmh7T24dVBli9cvwSR8hh9yNwCtpmAHiHlEJyxgu5ULu1xrcI/
iKTzq/ZXdS364iemkWxP47tfFIBwabsE4OefW8kIyyCQlueKS3Iv+d0Hf9Ktge9zXcL1SVJCYZRn
EkfdbzPG7BebvGKuQFfUXNt5AZrk5BI0Amekn8xX08uH/DC+9F0DYId1kdBZo0g1x6hlS7NpzBcq
gQM5HbmrNSrnImB2JYObBpii//QA7rDpjudLhS4HFTm+Akj4ka0134xpD8rKO60Fotukqv/UCNQe
2unhXc7fECWzIoM4oI1jBemyOk2O9XDGLCyg8Odqw8txmHXjOcWffLw29lAQQPAka2PvjBe7YN4k
5/su50NzYsHvua3OH95J8MgHvANOvnso/kI1X2oBB4v+R25Hrpq+k/bTU+X98MgUDXEkKVrfE6fT
VHYz6pp24l3YYfNUTEaWUyvHrlziXF3/g30VOwxzjONwLlZjRrEzhNDJooaf01EFrHpEzf/Ekmmx
JbH4bv/xxwXs1yzcabmiHawYecPsv4gZO4qnS8pqo937/Y882Bb5rGXl497Y/wLQgZXRsGuhJRAJ
p2Cqjvw7saqqSmVpW8nVacBInT/iqEO5eNFYNZd5L6byTvcQjMA9r1NEQORbIvH4GQ/EJex2nqwB
L7kAffb5nid+NuIl2Ihk3ALGxQJKAgWhvu5jxilAfCPLii/mAEJTs++odVSDLv8jP2W0Xld6ZDrn
FhK8/3BXryLuArxZ2nONuaEMwyixQHCSS81IPFD3zL7SF0CXAS54iW0Hrai1PGMUZmOmdRAVPCbJ
QCcW6e5x2S2aJzWONDx6F6Eq0vEUfUXEdigAVSV/burfTqaQ4rKvMaaJvPrJxOgfIN3gHy9FawDW
26oTSjdhoiav9EHBYcOhR01+6nOVWcdE1HyFY0iEfEsnr6X/GAmacSG546OXeBJ6PqbfpW/22Mni
Seru4+EgB+ig1/skzL6qCjlvVsS2BNPJy7Lc3DOhQ/o6ho3e8ft36l7GMPo1vIpsK6TcvDhQg53W
q/5wJ7RSlp9bm4wm3GcjLi7wD25Zwd6xC5BWpHh2uEC1R5TilIIqTV3y3ZH9QYE5Bbtg2CbTxgup
fOdNcDMApPR/qn6b+yTXmu37wkuQbOGISUitDNe6zzZ8rHK2zmiJ1aNlLHz68vGtw09oWQL7/5/f
AlRo7I/FrMPv5gR70Miu2MSzcSrdTVhx6fcTHFojBt7BPCpH/LZXyI0R8RT+ZPJqdJwwAn5Xfsnp
6T1rKiXK/6MDkhv+bopUdzOo2tfAcPz5y0zHKo+sMwB1TDAJX67iy5/H7VSJKzBNshx2lo1qQDPp
9q3W2c4i0F9YmsWZkNgLWvKZEOASkWdYbGQbc6rz3GxOuIOf104OoqjkoFaFGuQd/QoaQOHPkv0P
If0eX8YGhqOqdmH+GYztC141nmRPvExkr3xH25z1QmbkyUqaCIYefrGj2uihcaX5OT/X2TBpR2Kx
Q+iA3BL8iLBu5nV5aSWy1i4ayF9/F+ac4gMprUDDeXii9YHKfDRSXXS09+c17BrCopKzMF6p2TYA
YcI3a7kIJfy3CAbA3z+EDqIfq4i4+D6wLtbwrHDCQwu29ZxjPhiHp+5hwAsf+AJzUhqD7gR10gfV
z+VwL634qxjxuN+GJyOQLfC5gMVeIo3LYKC2SKoZ9beiuQZ95gfir5B975NKk9KnzaO8XvtdlDyx
DTa+HYbejCZNu2LlGjqK5zLSPBZQ2PTvksf70aIbLIAgMZenqpit925aCX9jlbHwMEFgItRJLfVD
DCW3KRFEwXttmBNW/JZPiiK93Pc9utqRPvFBFbrqoEtJEq5q8/gpL/LkRaXzosPkZGWlZiIlqF1H
/cEwbhak3jrnL0ddfCzw7tuKaiy5owETIosIbaeqSN/ycHnd/R4S38g83vY+xRr5ghx2NzNxhIn+
78gAUEwxWPKHGc7nUZylUS9/Fzk/nSLnGC63/zwDcya/zrcLz5M3W9/dbYtYWpI4Kj9h0rP1jI7k
87bj7qcfXx7H1Ega5QXwPvtgU8HZMnS8uuUzrEnxyR3BK+HsIJpNJ6u+GkONE20qZse37tg9DLTA
4Lte78ZvNk7qITr+z5nUcMxP9oeoCZPNxFZ8FX6mZs8D4LN27CRH/pZyCGkXss/LfEMQ3z675TZN
Nwvj1VYxjfcuYeEJBY8sHr5TtutTM++5SsWAkUaeKVe2SNPCr25NCXFrMycIHMPLNz+g6okupttg
UY3HzlNeJdnxQnqaU3TEDEPxKazKQRoeKyW10O/ltbFZGbFM1zcLBKvHDN9x9wiMhuVLPh5D7XGY
OkPLxDYe9tWAw+MYaHYyZi2M1UFXWCbd7O/CAWjv3rieLHH/D0cneYWeSjLgtAanhP0C8t4I0tw1
EolnCm9SC1LZZxJgNVdCZyXBcgKOOksf8yHtSzu9M8qbyZIPmIo0gvDh5svBcHS02vGirMTxXun7
iVjuUdCRJsJIJVI+syCQPML8WvSfMXP0XNxetuJR56ohLxCH1F/3OQG4Di8cTKvpr30QKOyrWUxH
67wKc1pVujoebPW1zcedIU6lLemGvng1/+t8x5RtSKZKRWez47LJeOoNs23naQa3v70IyNm0jKoL
gx2NvQFOC57Ugm9UusYN4odpg5vTgWQri52sesmhaVUJ1P6IvMag3GEVdYtzxYzaQ9c4aq1i52v9
idSuZzdMvqKt6KozqXNDmffeFezqWJlaZlkUh3+tGj0O/zwdMmdJq7b7GCwjO89VdcYDrQViCgBG
XZPLYTSVaKOt5oWVE1k+b8b3ddjcKISnOMJ9btoUpoBh/t1Hv48qtfrDCkdpd+k8OGzxCHtt9hOi
uZ6KLGHkJGueQ6zrXaSONill8kJRUSK0uCRuXdD0wuKrnaXz9hOq4NfhVqVaPeUU1aX+GLxD1gQx
p9tT0gBOoDsrBqlcV7NwmUtd8kY4fIai1tAa4UwMDfxMLlq8v9mXr2D0mFbac4MuGWQ8oP3N5ixe
qqpj6GJ7pyufSZpMCkKTsHnJL4iy45mf+XoePjQBbniBbAR0zTn9CuIF/fhye0hcK7d5PJmsOHDF
Q4InhYsllsuBKpJHiamEeM0dlCwlTVWc5MNCietbYJeFVLkaeF7yr6p4neC+qTo6fwGxssRVTc6M
3cVhI+YPO+ulbVpI+jTKMMlCLq214IzSCRr2mkSOC6EkeHbTqlv7HuwYy6ONTnPAdtTXn6tu2Kor
ahXLryjpeD69GSNYq6sDmiJJaeR5lcbzSImWNVS+tfQS3Aw2V33c3mrl5Jf2JNO2MekjddCFY0dh
OxfKK0qWLZ6mY9QEpvU5guyYfedSoiz6sQLV7N+SswLl+a3Un13Y2LPfYguijINSk7HVNQCC4fDp
w7yna74zK1tkXv+B1OrRpgGcKNnHEVoBa4fKx0/i7M7+ssIaZCEE1ZTM5nFHVl+FRDljrM83Jp12
G52X6aaw/KC/e/2xTfhiXcCSr1ogYeFcvdbVsUuD1olo1peq5VPPKErOOGYN5/kIr7IY40vTmfhK
dEPVStb21bjEtpMMy8n7bVkATUzJew8NJTHHNDiCtrswL81l0WtQChyCkAwyB/nFuPz/Cpt5xGP3
6mk4BGUnXa2zAqByTL1r7S1/Z0oPWNsJFJs0D39VBO9LKlcKFVCWLYKijTG5YPt4Ml/2Y25zG35x
XWhbvtGxBii/AYIFJqBx76+2+WMsFCY0DIUEFB8CpqtFx42yYmaf7pFQGv2xJotqNydbNOwXWvIM
E+oeHo5h7zbpNaBCNhe3+AYWEtdogbq8Km5SpjRgEId/GzPRPzlgHsyhUpChWsjFx6/kZD3bIG60
Snc89/35M29LkrlaWvbki949RuW0hgRySpzrLV4YgHSXLwlTMXnkd5gb8ChjsHxNPxmNGnVgjUvC
Pys9bh3a2NqkU99W7GHH4Np7PkEAYdnt9U1AUrocVhODBmsTM0XvAj7VFQpmIbwOA1oBwYkzEgdh
fwaPIJ1JgnNIFgd3/VkLNK6OtRtyaER0381c879uS2rdy7u96eyzVYFJuYsJGnHkam2mBgzOViRj
ouSjS2mRgJ6LxTIsJQpBMD6k4yTDxcAtuRZQtEtb5NI4fXK3owfWHB5Z7zI8hVfGBbE8ge20Zezm
6PEIkDOqusxYVkzMHGUHKvHvBmNIWxVzAfgB+AkYfk7JlS1QhcmhhKVVCmlyx3VDXv9QyNKBtoQM
nz6tmg+g2KZT5+5SYQYFN84N2t8TyA/DosZABtCZlozSv1i2NXgc4IrVnc91sFdlttxNOp+gsSAC
Y/83mJY5218Au8rL0J3ClSBU2/3hFC7uFJvIr2575ZU3ne8OyRLozhg8CO1AZkHtomlOwJaFvTxb
8bQEnSwnXIAuFcRf3tiKhHFiDP9opw66Ql4R7i1FQUxX2WCi5gM2uYhbDUsc6uyMJowtP1lFtTjC
6JK6w8rI5qrhIv7khMCi1yxpHFiOMwZDkHR6L/+UD8YfhkCYsW/WoTNA9DzHGVHF9oAb/YDXd9Se
xiureA+LKbjPAI8qQIndb3OKTnhgYQLe2NoFDGN9MSeWzH65MrYcwQPOgXIanaKasUIH1+eh8nP6
g2X20fO/08QwnmjS/Sp9AQUv/kBgtSAJDDmUEXUtfOd82RiTUbxbuShHd+sCt2o2dY84eiXI9U9J
3VImNJ7RL9FnEkfD12ZbmN2leqiQGXhPgNIMSSc+po6SPvAmLQ9GdcD61j2Bt5wiQtI/k4aZ6tce
R2SR+/tLA4Pno9HgiAt94pFbn7cbuRLUrUkFopLJ04l8p33cXDc505ZjFbKnh/uqJecmSwO6EPbm
R31G6QM0JlziiuHP/C2upq+RTNKLc3kypVWk+M/WHGyuB1pDQwGHrk8vz869u8RfX5ZnWG4SNZaF
qgUG7xy898LYnPVIe1KGWvHmPj0ehitbrEJAJRrjcwjdSDWMwU3wvF1Xcft/YQt5wzCOw4qiSvFw
pZQbJQM/AhLS+n9TtVI10H4m9HBpRQcwYPmLRrXKt9WGC9VxEF67i3R+jl+bupj8WTtGX8PQSDpi
AZmLKJrIZtxSS1DAXt5tLXrud7RmVVJEz3PntGCdzqoZaeZXr9JrVPuNSNo9KsBVbSTbtL+25Er8
LNXIoZma8OrkuKuJ9DlwbaDEXQS323VaZvDMmAdAhfqSGbOXiftfzTNzy3X/8VvAyqUbyVGyeoft
CFdqS3+TzDw/cm09cg0H6Z3fp4wcc97wGXfjalKn9Nxd6dY+QZARQAoeB+y1HVzrKdcN+a95LAKL
647S/6qgGiEuLlxED3qjcEDlgqIAvZuqx0lXpenPQkecYd70FYZz24kQ1KKJFQ49ppmHxMu/uxqg
PlzqDeYsT33VJ8mqoDTQJqxrEfoKUtn/FacPIDqPDyYCc44cmpAx/zWCYCXCIqhee2S722uqrHfB
qjoxLY72S+qxAHx7wPPRP5uyrXL7Z9dxAr06NtO4kwjTklX9MYKerouRycRUNcG6pZmQ9HIf0lfy
piApb7B2nq25oP9g2vxD/rmTLxGSfK1OO20AP5vi2ThO6woOwTxDSxeZrFT+Va68nL1WyZNFEMzc
Umf7fu1RE4Dyx8IzivQnOnAvmHpHXfQ0oPc3huy86AcfZ1IO2wW5IlRjcU1mMLo0O1zUNd8x3KPv
PkMa5TNhJs9XUeEp6kScqLTXfVe+J+G1pqJP5js5hD4PgU+pMfw5/a5Jt7hYggE2q69qJ+73370m
Ye3jBCQf+PPUjT8yi3+za/RFluUyB7xaXlAGJl2FKIv89OnBKkdsl/vjIf9x+SF7ioUHSJLpBWFt
5q1sFlpolp1A/gNi2Wp5AzbYzh3jc8Aer0trJuPxqHdoSP8zObzlVUbS194rlFz7jbGI4V3cCyTw
ak773fEemb6NxlKogEAuzpIMp4ej3Amdj7SjPBWyBTia3/ga0C2I9THngGm5aBJT+0nLL7VnPZzO
0t4zLA3nWWxtXvlqplrSnyvGY9Vo+fx5uwCkY9gbL1gpTM8CLuaIsmj+XvE4iiGNv0IpjYx1DXnE
2jx8WT5J8KK/qdddAA16CIWogeSVKLA2INMoGnCp0EJaWDhx8fkbcChfUnsapIa3QNyhAn66vx9s
ul7hUdqqAdAwk+FAyXqWCY4pZr1oNf2ia/W7rBr8WM6cN1wMqEP4LLFWNJxxUTYfZThDd5sLwAaK
DZ9RFrRpS4vO3wA1T8ZFyGI10mjc682UaT8J0CYqewQUqywJzQGdhrmljKKpGVCpDCk/PIZop1Ko
3cpmEwz6vsw2Gn2dqT4Je4JTaNS8TUy9rliqOTQZAjDNbBewInCB3dGw30P8oi6nSTvf4N0+E9CY
0K5PDftZpdplybyf45quG6gGfaXvy6bsK5SIJkk97upvJesysL9iOa8ZZ5j2rI/4/ixiKNhEpCI/
vPCO20VDyBLP8gtypuVbQbhaBMBW7CUml+0RO5QfPcJ5BxiwPa2V/KKJNCwKkBlmR5i2Az8igvxl
3Uq7++ZZyuXfH7LEOSMtcDDpzfSxkivdlXX5ONdswsyRR1wK9u2A5KWQCWzLFF+84GYCfriH+jER
9ycnRz2JoSghN6BMhMFzF/HgrlIo0+tSTJRySxVbj6J2iLs42AXHq0LHAhH+3H6uRNNTozV6SlaD
vB1YJ3k5Lvye1GN6rStHA52gaV6r+j+oQ0zv6LwZhmn72P37dVvlv4cPWhaPZJuJLuR+HM0wnihl
gQxIp5mDjfZ7yabxJgyq8Gkz12q2eSoMzjl70U0WVBUu7s8d2jWL700XssVzcvy5xCD8yPDNEbuO
gEwFI0hz9khgHRDlDrZ0QBbgSWTGRyUoEZOBzrG+SP44mOFr2l0oxnP0jO+81H8aA2eauunNzcMV
AFsWKZySHp8POpmayv1ValQ9k5/4gFEDuy27hlis4NqzgsmSJLCN03qdtJsmudBonvx8/0TYfRTZ
0wKCl/KmJ7MVR9Uip1cPaLiKf00WG0FR/GFFqB7P0grltyAaUCFqbo/4fjrPGVwrUHyY/ytRQGnh
LhlRBlJGIwWVH4jQ9pa01ODpJ0FZPbjXK1VeV+Ot3FmFLDKfY9hIWb08+gpNrvrv5e3bdhYgGuBw
jWxFDw7NAYAzRMJ6Mbx+RYDZJBoXec4aGtR2GfYKtJ7E3RTlqESqiabhivw4GZymtNQuY+C2F8Ep
XZOWEYsrT/O3c+h+SlMpVl+xAAHq+rQCvTjK9yLYIpN/dy6G7I3bgWci3arMDKZTTCfGcdeT4wYE
w7tCsmmGL102/38XrIrUoCV4L4+2T+1CI4jXzKnmYsstH+XyLY0ERLh8wA6RkKLgnpxxy+xTPyD7
NwvBegAxeyCi4GC3QZ6fCbRFRGvTCZmJhscgiLGOTCjHJBLBAjPUteBp0zXZbmZ01opUhYwWunHr
1bINXhUiPK9jksOHovBOUWvakn2VJCzVvumFqNV2DfaFgxfwBZi6pdtxp7VK0Q9MolzK99i7+k4s
an4M90CBMvbnJTB+H3Phtj5k6xbcNpNZo6Mwlh7ps53vQ802Cv4ru2O++lQ8UKewr/M5kW4ZdK9f
QydyGN5qPJGcxdK1pCLb7rD53l9+ZCBaYYwCwNB8DRwdaf+eg+dnneuvHiRE56Ewp4HAK9xTK22b
bjp8/3Gn8p1EFXWeLWtRTWBi3HnqDGQV47TgefWZ19p/qmr1WVIQyCYJoXFBjd60jIGO8TZkYpaT
gnsDRS22QRoSGmF3ExSipAVl9qwFuO88nx8GcMTWUj3sFm5HIiYyrIUpzvzJ10v5k6IZDBD8CpjC
qKt0dUWz2kJV+PDZZ/bq5uCKjLW/JjT+JhdcM5twzOUiA1sknNFtebPWv1t1R6BZfElxH4kUuiNs
aMGhrsQAr90KTvKJU0XN9gIFteGLItETEZfZMb4+MyVFbEvEPiuHwYFetff5B1keRdjxd8JO8jMA
CxUWkRf6F4xgJEM97n7Bb/tklf0wczJjE/FHrP3Ko0dNaZQVmvwuFg+3EzGfqCF3UNoDtZSrRGBY
iDwKtqvKcqZ+sfFAKVsCVJG6buN8mX/ZFbQPyq03i7F9DbsqLdN9m4r4bVnf7x7irSQ+H7gvQY++
aH5P39M7p65b0g0UhK/HTSGRwNOsxrdjThh57q1Tx/oZN2lT/6Cq5MrUPbdt3/5DVc4jTET1WBKW
cD6+UEGkMGkHTgoEKA7RaduAyC+6v/60cOPvFOnRLHVVHJ3OTiq8466OdNvBBDV419ACK6FiaOPt
v6uxhosEQ8SBsaDKNTEdizDS+Gi9v6GgNtVdK4oDGRf8qGzHqp+x05EHc664YxLRjyye5GRbFnOS
LtdWWT+2LjsWhZACWkzcyAxZis8HIkRTjxd4S6gps+KcmJzxdCV1uq9GUoS+C1urw3ZdPW+UK/Ut
4V5R85wBpmKaNNuq1eMsGVArLZFZ0h0KUwUuq7b1VaEZVCg9jSwwaXtCjeoeQbUGwCePCnybk+m3
eblmB5Ycaf52ZY6CNwGittf/iuCFES/d0SCroSOnt6C0WeNTW8ryuaAHX6b5kmDPL61AnPJkQfDU
XRTuScNWVp5SpyOPf3WWBzDrk1U9WFQDGqsrrfbAilulUJigo2KhWmPFIhCHRSnAkypqtM62EBq1
mbX+Xkn/7pSW7NnTKYHnnyiIgsSt8TE9b1fw1hnCx1rep5sOE02JhULqAY3yUk5sSYxPv8HHXEnN
zr3Y/4VqOgm/jATpVv7DrNjN+C6MXWyW7iT6GMogQG2ZAyrvrls/oNfbg+tcqI6gZ3RgU9Fq9ad2
0ZBA5XkLMk7fPiPo15xQHyHsc4qLaRzqLBfvCdMBTZi57rqgNJyPJanm6Iaow/aUsIU/eBKPlh9e
O0Gd1yKn47om2/gUNrU2/P5UZ1PwHRgDVhqfhljMM8AcBiw7r+t/IYhiUneRDdvv4LgEGOQDWJju
yhaHRPwi4sUqQsh5mSq9ZP1G18oOzj8RHYtVEn/ChtV5Qle6PDQsyZIXc58fFzTw8RMz7zk7EfNz
R64SMPkmvYLvZLZWEPBke/Auq8ZDJjBD5LP5/U12BaPL0KvKQo6NF+uTi5pbu5u5TKcHDBTbXJSH
lUFp9MGf6PkP6RzbHz9MB6z+OjOaQ5Ib2NvoDP/tzSMhYFkt5ggR5sZZeQONXiEy6TWA8xicAt1P
ZJdv0hugTCRc6ud/fHQTdRVLOPhDh1QQgrKeWbX3rjx8bYZCAu7KTe3H2lWwiC0irMGH/7vRCSID
5SgN4FTQDncmKMUOZmiXZ2ByBpRsJcLUEMd98TJ33rvA/QJP5QEvAGxKVLUJ8c/EN+xk4x06ufKM
XU7GyiX15jM2KwyIsve7prV+Lzw5sc/GlwgYzFTTI4JB+NkmSz0qMTmNGwQuiEnjO41Jc2wjSUks
PmCI1C70DM2P0RPKeCfT5FiYWKf+q/rDrEQoEegHQ0vV0FLJkXmPZf2K5zWSAk9s45dVbQwU6FCu
TCrqqFFfwBWq2ltgROq7Py9BaB+5yc+j824ZPqP3n9I0FmCRiJpyzWx5zAlxa5lVH2Xmtn8rmoNI
D4LOlTEMl45L9ef/6FoYgx+hJ081Fq5CEWD7aEkSbd2mvjmlY7F/ysB6wRhKtWgSlnMJFFQQvG+X
F1MPBnTo9tRxeJy3WzqFZYTynK68VM0hY6fNiVkxLr73e3ICTxY4VCNXZ045LOKvXP4tDIfx6vEl
5t/MVeQDFTymt8EFbZ1jhZhyX40h6ckieESgf0OBrO1SzibAjlU5GLdY9YVJG0ET0eQs4/2ZAabr
E3c8FXaAat/BAt1sFJBJZND3a3yj0bq1cGCJJBPzbAqX3oAwzHRfYqSJuq5gJ7dGyMWfDwtjW6e3
scXiWSEjfwK7RSlAnde+e81sK68r1Idd0IKwUGoVaKGq7U0voYaSK7lp5DvF35b3QNeGetWLLg8g
4RGlfekuyZFSo2OJO2uoGRi/HeQwsH6WrAl7dkRyvFEtpXtSYYHFqFh+2UG1PEojXaBBc3ju0puG
T/fW5ZSAuWrNBb9oA+UVXK258AAmqBp/0yAAx0NVVBek0ZwhbKm3jr0EDAnyPB8erUrhX2AQXirX
l1hyxSImNP9uCQPOF0pOweu1salU9ljS6s5uWvNhGGEHF+BCZvNf1tAtIvzN2g3l1J5CH4qNNpSL
nicO+4K3uafBgcqMBfFfsYunpe4t3T9BZmt33Vb3kZ8vv90vCGI6QXA9T58PPvjOg/JzkkuOBcJY
v+W/DNmlAZ6qEpHZJ71h+5Fi3Ni834G1MiMCVE3ym5FpZpsxEmT5ejmrw+ojP8bzsn54OrqY5ojg
umLgnM8BbhnLkwQfW8mENVtQkFfzpYeYFwh9XW8XTlzEFnkiMq/pv6iVnrpwkg8mX2tfZEJbAhRB
ge6c2mnuTPrdSl2p1dSZFgIQ3pgWU3TSA9OMO+0dvSa8M8+Ad5z4XTb2iMtggKctYTPNah91/j3C
M+1/aN5fC35sf/E6xjqx906paTyJpSAvNKyvJa4jomUbUKH0kTsAH5G4+C1AghrgkLR2dXmk8KFe
3PWLDcwDwurqNXJb5xtKEU6DvTmeJ32qE+YpqUHK8b6ojqKuDwRiIkEDoWzxuQNq/rKPEpECB0OX
rbfpm6OV9Lwn2rmpXL1GRpjXNAD/HmTSK08P6LonihDrohI8sjj6a5dQg0YgGoWQUjmTZk8wWZy4
44Fykt0BD5ogAamwjSQ2u2BCWUy4wR4bT6fGU1CEecgCjdHPnd0wzsmNYaLDfViMlO9O+r7Y7lgZ
1dQXsVU172KPeLvSZWeXiXIJZSOfGN/jMiS96J4pHyqDr9WaS2nc9JS8IQfqQLB+l4A+MzqpbsJM
griaW5zfcbOWHMBYnGawZRSZqYmBV/zEkMCakiGpW56W9mdjb1vXSXjV74to0A9lzEnIS/hrJ8Pl
1EFrshtnIANmUjX76GcknuuY3QtsYDQZJsptbjbWjT3oO6497dSwYj8KJEF9Qx8w/nl1WdcZfNKw
HHr+SPr4lGr+CC0WD1YGv+AEq6aLH/1WjyUdVXahstjvCxRi4Nlj+VgdrL19A8mnXlaP/J/O8UeX
XH+O/d4T3tEd6WZqtgTObedO1TgOqDGbWEJkxYInTN6PuDxXz5JYHBwPGHWnGcbB7jsmjG+jfYDj
0rDK3VZBXUnTy6DGy0iqlxXOD9h0k+67rUk97t2Ytz5Kwq+YNRQcJ/xl8ErxLB89w0vOzbmlafmW
4i2GaxEvGVY2gD6jA8UQWRCkGVHVXeYnycu1/Sdh6udNsxLb8P8rtNXpMC+5otRE5TGcHTbhbaWn
vrqM9dTS0eo5Z6j7RLnqqvyvy5Fog27Iql1U5vBNnciCI+lW2j/ItDrPGU1tYs0WAOf8mxadlMZa
p8Etp9zzWvVsT/3sjMViqweLvwiV7Q35yBAJJs4d2YWAYrOQauwTW8igHpWqBqIwzzEgu4TbaJrE
8hFT9LD+a7Vm3Ivx7ZT5AkwM4kuZixVwgImnRNqSGSZfnW5O5tcfPYOPn7jabaEDlfFk1uucNTGW
4qsyNH7jxj4fRr2i0rFqFw/JrQXh5o+p3lac5xYEXLiN2Mduh+ysKu+qINumoDmF97K3nfDOQ+ZV
cVJNh+9UCgDVt88FzsSXNSvDYkkTNbjxyBlOqjTzMOVR5QQWEb6kzXCEauf2TqNHCbNuPK55glwk
LoFx/d4rxavO/Tz8t2AmanYIK2DUWICPgUgGNo9Q94bwnq43dXuYcGk9qALcceol+Z6MAuWCzlbD
6dhKmswf8shGcmwHYc4CUXroXyOy0YO6cLgmeGwWEL2IshM+FGeA/qp7d8DLDBI6cFiczGK1iie4
eXPCXT08SdAubs1AZtVPd2DYZ68KKARzEpsr/EgUqxnCZ3dTYjxZyPtXhvma5PFHYLYkBnqqZ6NM
yYM3YHvfZEd20JpgKUuUZiBSc1E98wMe8CtyefiDpd96B8WDqyZ3Vhklvg+tWtXBV1rnJyWERxup
2K6P6e9z0O+LzhCqP1g7oWSoWXno5O7eMACwknTrA0q/LHDQEdCaJOOX2xoIn5kApus9GN4Flk3c
Kbg9hijHCpwIllyjR3YSPS6rvBV4q6d3H1v/xBOrwIhsmmP2CxQY/NGf6P31kQy4VY0O+BChNSkO
Z+oB0gtNqpRr3/QXdl0G/xl1fqL74FU0B4hINhyEiqywSoYwGx0pR4JOKYxU/i2m7LEbfBb92Ta3
e3xi847j6RDwcMs/uqV8LqbAa0rimJrAkXg52VtA3k1BsSkL+ZDRk33XW8PmrFUsxukXxaUJtZnq
3z9DWz7Q47qOlISlOLHNGjhQHPPrS8EmJDIhj2EZKRL+DfIYRnidhZp/C7aJt31CVdFuQRG2q/Ip
eX9kpmORcw29V995CCBI8al53Zw03uEksT+M6V3wc8+LhCmp/0jUlvAZXzqCZBJF8R1YSjiyt1hr
rGsllhwqM5mKqYWMx1+PiF84p5KDBEvk8hrCp2rZuLw0VZgn90Fnv3ZXZvS80xwGV65JhAocbBe9
aul4dvecBv9D388d0LX7hL5wOs0FB5MWamoSLKoN3QZ02KQJJ3b80krDaBnivv9IxZzrqd942vno
zigVKqbzbijY+fw0KQ9z4Y1PQZ0FFoSiYnkD3t+Qob0X22Gtk3oOveF7v75zGzC01xwqWxIoQmrw
kjA5EHVwUK8aBHTv0wfxei+2F+RGCgrazUtmqUBIVwiAMmymJduBIQiMh5DzFMD+f2D/KNU8ZnmM
0dYmaJZ2hpzhBE4FXXjP8EuS7QujYbEjLpyda7GpP3LznnJRTh9usjn8AR0SaPDsFHp0xiUL++B8
qoDTRg2eLaV2GKIjwBWnwqRLci4R3uFl01+gbKelOiY1hVSjKlSEE/4vBcMb1rwowXnO93bS3btY
+G0TpubNwBro7uYVDbQ51C0+pBG/9KbR4F2xwk7rVFvMVGRb3HRMQHyJYHjqAoLjrTXNqXVqxEow
zbecV/t2y99FfcBZ132AgOe9OJt4/AvhPkD1D0g5Ae0KQhT+yrb/Qx82Upe+xme2v+eJiIRTc/UC
/7Kt/lqvgzuktsknTQnwBjpBjqCcebim3C2HW3E3MK2K90F6eWYsELBDSR2KZear1aoetN2cGI75
dxe2keDKU1tObf9fSnEIXO4G3MB6biGGt1o+9H0GTzLpB5+bqtVHTE1r7L70WEI8qkk46VUikMCY
W3B2a6jo2k3VjoPaVMQ+BYzdIezlXWE8EDKFqxM/msxP0BEnwHxefnQPrGTUZaXiOqCJ1N0B7Zrt
0zHZKgsQaN8jZI8EARmuWrTh/l/Urk1DzidwQPoM0tQkgiFR7puZ6R6xRoO7aPAPLfvCpZNygK+u
lnF5LnmhaGWPR0eDmIb1U8WqLGRs3j0XHqPPDYy8C+kz9xMb5mE050SUqclz1wg+fIeellRkmXTo
cWagR/qb1bWQ/e4svnYJq17EStBjw/YJLuUFGycS/Shh/p026A33rPMoC0FRO1Kk1CwWstU17die
bm/OmkBpIcOtn9d6INpa39QJGUn5tInnqdyW5jZg6lbHWOx2DjcHnfoRL5kAMlHUuAdg21RxkHvv
nNuFGu44pOuD/knZ0CiLy8gbQXqdi/qUOFjoDaJ4hanYkrz0VwXVWZeD0VPIH74+vmGJprf0Nrjo
fOjGCtfJ66cn942JY7XrNbVZOF+QJn1N27JxPuCbKUK97uCBjK7FdNM0LWSEKIaqLFdS9oVZuxo3
jZI+idydiJWNcj2yoKxF4FOmH0OpggoceeLkEUhLveStxOXHvJBm1yTgNqwWKlkTM0/PH64gW2zG
1KS8Nynh4rqLwcawXyVDFbLTJRA2q6zEEyXj1TJ6cVchjh2n+AjEK64pU7CBuvWeJAwZ5z7u7uLV
7L0jL+HZB6KcqgTX8gmPnMwxDI5vTC5xO6v+WZipZ/ztFzRgVzlSR7Jk9EKNjobrODN5NKENpNiw
MK4dLCCGG4f9VhLkLJWGu83qrhUqeUK+HGXOPveQsNlBO97OwXFcVMQsCZQT2Sg0hICr8A+OzFcM
WtBw54XA1wMb01gFo23s7E8/zyDXVgKfMRXmfEez9oqYA2YbQesr8mZ+WeTqA3hDQwXgelfjYGK3
/4I6io55MS6U91MWaly0u0C2lL2+KsH/0pVL6JSTmIKtt8r3tpxhbFSmAa3c0Y5iN0oSZt89UhEs
KyY4BA68wTim4FAfurrdcdbjOGQzTLSWAUcql3OPj8/p+ETBtdBuPohjHABsOWiejhZFx+AfjeGV
nxwySA7IRi+kICV00zG6rYLjPwdjq7kv77f8LvOxI1yxWHfTyh/mpXqWU9g/OEO5tV3jee17pdwh
yrYJUs9DX7oIAXtJp+5R0DTCYUw5DPwkRufvkQKCdydLsZTUWNSJE5FzoocEmzYKv/+s9KRJ5XAU
Yf16QuXK+s1DZ67fn+KfnNrXibsrAJwNQw8fpKDh8Q5Y0GTSYYFc8HvmM0OPIN0KiftFuwoKx/mD
VKcYPltP6lcSDJ4frY2FVecPvibqyKeiwHwrdSzQB6hR4DXask2PA6JEbZzMJqX82NdCZ4Hc5u5V
sKv1Rj4KBHOIVFx6jugHL3lbag41defdtYAK7pb5jOaSacOe1Ed8p/AsrWwmqGnb8TK6qW1OZdBf
udzV/oB1jQcyE9zzIRzlHJ9IrRgRcWYXBABNt69+h5mpG2un++q58r1jdi1fUH/TTbMrRTKEMRqG
yFTbbj9qi3KxXHsSiaW8miA/mhpHy8uykTkUfXCvF6OxDtC4aN5R8qDl6eZl8SYUi04mu/JpnfD5
qw18jmEmT143YC41QpvJnwYOdz3ROtVe8oBJkUXgo1u7TbCRaKfLndwwCm7WJf1GdZEk07zmPOyZ
1yPRfLH718zs9QESm9DmP/riNVrF/UMSwtfU63+Eo8l0FQlQoN8Iz76J+v0N1lQc5weUktcy6ypd
VoN2CYNn8Mg/sGI1U7U7mTSIS29gB7FjOPpQ9FLUyKjJxzhLc1W/5h0xs4luq0H0nyV57XeQxUa0
Hptg9v29yA98vdA/aTSHwgYhYIbgHCXKbA7BIclPzI3AhZtUDw+VdhTFoSFdaLfXjRSEW/bRsKre
rSqeo/fL9/s+kAnUkn3EK9EFU4DFzcbWqQ8lRhl/S8tz5lMq4+4HN5c2tjc2IpOxY1w1pkj34ESQ
fKhUbKT+EMVWN9zar+7dcvfs6xBLIE6FAGgzYTowo7TvOC+hlVB9AmwhFWjeU3eId7iIb78xDeJn
cbCjbLnlx/YyEg8vtW/n7BzBaoodv603GR/rilr0i7ak3+bFI3OQNV13vA3i7wHSN32G6x1hC/pm
0ORw6+AzlwBQ6FfFK9In3Xr4idfDDFw4QLe0j6qf+GBREijymSsmHnXCJZiYLREs6cBCYV7+8FPg
WH6JCCI8ZrMAp5Dla0rpFEvA/rCTn0Wp4NTIH5kFhrQdIlpPdbcB0tUz+r86YSuv/R1C5mZfTIG6
IKYHt3YZECdX8mf6fED3+22jpAaCklPaFKxhf87ORD+zcDY48VUEpGEnTqzB101nG7UmsHW1JdgG
AAxqkL5Kdo4fWs6Yhs8IK29ouoACxrEV5VBkcvXal0K+yrq0NTdCAYDB/ZYzkTs8CtiwD19FRyeD
xuF9AlFhW85SUTztFS23FmIzR7LeSNrET79K+DCBxAaWVaiwXbOuFpU0ejcHZaO6g1a+/Uxk9oeY
Gxf+1GRJUferiU+9LoX2oHHx81qUnjtIxvueVhyndorAJn5MNLnxyMSVIRPSMn1YAMVFDjoNis0N
0VtngWUz4f4jfxX9H4MVAUgRNhK3WpPVAGhsdkjV/ULmYi+wZGMzijgjPlR9yZtn7pNLhKC4HzoI
SBxM1DrWlkYJTeGPibPFLL80yN1VXvDMe8jJTMUFgsD3HF5pvkX6TjVhpLWzLOcFbXD3bvA9q6bX
GObWTJe1RVZ6pp6jv0re1XTWsQHLA/mDTroHLli4nE55LDYF+1Ea4TLt++8qQzWtAmD1fmiF8zJR
eEBglyAbB9jsq99fILOpzjI2npDu5Y8v7XKaa6XqdWDA9M+jr42nUFr6/aydHvGjK6mxTifzEubG
kG8dSdsQqKMEJAJnumgKpLwy3yF7DMNuicBJMGrpr7MK4+PAwZlPDa0Ncn9eIctHYxxDptCulDf9
KhhP4YOpQ2m2glLNBYLGuGz2uL7uSbUqMIF8SHHI3Fn6OVxfz9KP5hKMHrz2Fr4JBoS1iS3rZ2FX
4Zx9M6/6UH78l0GzFekbabaJtl5pz9wb64Wirg8U33vceER7H32uZK7XggUFxz90XZ8A5L3KqrtL
q5VKzPBQt5C/Hq8EiCZVnjJ2ylIe+Unuu/kgOrIZNpXMDtuB2xogwmixYve6Lz+HAVFtpfFIp5bt
Ya6ITUKqogawAo/sGWczoWTTOee8kN2VP0Sbtoym7J+2s2xW6ye9clvShiZwoNRidKDfZYkEIqlv
wPf5PgCADbHn/1bkYPqAUl68XnYsFHtnWzkSYd/ApXxJXbM0Db/LiZerdznAdeiRNOmVvxZeVWXP
9Boydz7QPNlI2FJucE066itHDjkkfWKXkXNZ1y+0zzWITPAC+j6OsLgHxJmrq505ZCJT32IP2k4f
aSB5RGrVxiNCz9/AAXwCd+IitAHsTqLuNPHQYGW3jYSNxoK88Zx5Fqhym7L/cibesIYUMPwRaALV
x4M9W5FFl8Cl8ukR71EjUHov8sQ3IwwqXZkkOVuTONcsXcU72tByqw9LkCtl2T3WnHXpnLdc1j16
f3DUGJSUGmohz4HMzWKsiApg0z9hDkUdS/NTNtRLuRtZp4Wl2hmuIpkmc0eMCGxarXxkmSVzAK6c
dnmFWK0FHM5k67CTJZS6RddoWKFwRvfh9sU652FPGZBzxOtrpwp//peDDWHXYz2B5BCYQzIjCP0/
at9ZFKDyOdEo2qp5Pl4mm4vqjvWd8w5JDa3QBxoYDHKrQs7Dg5JlfOaHqwylnBQR/zCJPhdD1dHi
nlNtv/6ea78usGVs81zJz421iQxgarU/NmYSCsVOYpDZrEfn3plpq1Sg8uYiUG/jg1zqZERRe1xH
sM80zLpPuh+D7d8yS39JaedVdzN8p9B96zv9rfqGPw1mpcdI3JYgxtHM0EAYNHlcheXI9hodQqRf
LjFwREIfPj1yeG9JGP3wdu45t/mfrI3CV2sqHJr7eyB3QiD8w1gd4ZLfHiq1jZiPfMiYnyodIw3J
WDn9E8oCuWiGprGu3Fco2dlGL5mrtDALMboPQgdPbZRoMsrqKtBEOWufkFP5qKHEC6NwsLG727Hi
EHHge0yIJtIgIydTR1ENc07OPfdDy/iuxhGVCK8O16vVCoXUYibdd0nWRbIKUgnXHBZSvDE9DdUx
moBdOuBWcwoJJKpbUChQmN6KBEHMjzOVYk4U7DAUB0b2FX5LSRwdSY0eqhxTLTWagDcpTgs0Ahka
05jcoxF5e7Miygu65F3VzI1QGfvkg/FxlsoO7s8R8yGvdWHqAWlFyoE1lYzfOnqYk03pD52wCp1n
j6zGzpooe67a2lRPXL/anUDMezK9/skKMGvoJ7ZOchoCkM/YcHyrKU5gLMM+4ITfXXqQJJWOOghx
OnrWFqvJeuEDwxnIimkXFgHPyKaWstJ3z4rCDfoaJJPqiDI5QeTqwBUaZQ+4JVSMMMw+lUVSSisw
Qhy7OoV+jjEHgMz4M1xZr1jp+390/PaqE0l64a3YC3glCH40MSJ4mmmEyVKQunqG3ptYATXZurMW
9Lhb82Bt/SduKpbXt1BXwLAruiuslH816yJYaLPRan+jy8WkwYvTFXSxmKQtC/D2dI4ZrF68Nghg
f/aQVdui+qcKiu1xp9XhtmM1cf0MjiAo4FAE5MgzUPgxadQ19Bowklli0ZPrgIngzMkSoUvn7siH
CWtEu/8BaIL3hYD/31Y5eV9HDHx7ErUaFPzp9DGUhwb1S07R/nIIN0eejDLQCAEUYAGKkFWdQEK5
86+Ub9iuY8xXcO9obvL9nxUpoHvcETgJdGzSe0bRzNRb/o8UNS0RiZhBIBw6E1XRkDxXcZAv4zne
gmFQdqH4IJuGauWIilghGP73r4uO/tF5qsjLVSPaqZV0MA8F80SzK0FT7M8MuBp0Zb7hjWacKcBj
1TMz5jAacc5Onptf7ytQwxncltKnATmvZkFr/1uFrSquaQ9TQdO22dQmpJN12HuyB7sFt8IAUoSu
TVX315zcBMfAI7BuQtECDGVrTFy3o/YpIUfAJERf/UhrPP8zcHj2GoNd02GhiX09/rMHXi2WDNeQ
xiphoZhMhXJ/CYasr/iUv4DpLD0SfMq6kwilVWOyLy5tw2dwZ3Y1kSJtSqn+2av6kXeKLgLECtHc
0ZRMGrQSuE5HP8AI/S1zqt5ei8TmZXTVyLWBlqr/HNHgXmN9hPdpG6yMwI0RHM2NYiXwVZ6apgXj
rVMBEPLnkuGyLxG+potnid7kzvHwV6cMpVgIFTHv0gwXjAoLIWcCFTVZi6jdmN1nEZt/4Bzka/NT
MbJLG9nv/xeI1NDjRvLULdChn+hxntI9YK0HNQLODUgHuWc6Stky1DZnedxKPDX5h1KCQfFyLR3N
wuZTWj96OqR4egx3xgelCyAmFRj/UsOEPMtri7KBAOT+m7pDKV3DeCYUk/XSKgVNsMqDScOMxJIc
mMKbA5OvrLi9I4e43q51VRd1+8+6LBjA9LPGexgfU3HuQPV3Is1EKTNwM9OotDAoBPADVYioyrzt
MeOSBcsUNVeBmms0wi/MEKHVluhV/ffjlQYEndzZeYl2KuLUDbny8os9dtc4KhwDPDQTqaqIdcgk
GFAzypuNGlEX/JLj9ht/E7n2+dxP8lu8O1IMMR2hD3zu6feJ7MX+Fds98ojHTw2D6mZbHtofUskL
h7EmQFvXjMPmL2giIFXVSCYEorvrgQy0lYbBr0tChJ9hKNTh/BJeCMWdanByvzeT+WdI3bUiOpMN
S1IYqQHylrmkyVP6gdr0VyZJGMwGsFJU8bD6bm+yKGMVUimaIx9IPto9Ir7iDDOTDTbdMxKUQnd4
lB/c+YNOHlpm6/y8BPWWFOmeX/3LoAfxtF9c3vi2yLHIEgRCrZKXEpG0KYyXxjNGpC1mJxYem85F
6G6dSsG7hYhwilKkHecOB0h01jbWVmythcDH/wMCM9E+/pOBIk9RylIecI3gMm3STXnP2A60XlVk
+N/1VHqCQia1ADkoVfsluVYTlHBWzGRsl6uky0c16agKcRpr3PEoTsdN+5k7MAn4DKB6pkpMqYpb
ymrJV76q9P9TSbuu15vFIa5/f9qZHvgoIvrbhbwtbrM5sLSKFYu5b5Bhj5ovF48wTW3vEhydbG44
Xorv+8N4s8zPAsyHqVrpOYzFKCvlKnpqFkInEAWsGPuPVWd1hWWMjlswBrTHpzByggqi3vOlXt3u
KqgQFmjIKeAvHBWL8qQrF3yvN+ULKmxqP8Cd60Srm9MvfPG0U0W1Tkh2fFU2aeTuLecZJx0ufAWx
RsmCsiAKUUYY1pVoqqLmeIKEK76vyqO5HIuk0Q1JH4q2YI7b2tLr5L7BdpK0H5JZbICS741kASBB
2KDKlIWcIzYbADjQF2a0jFGv+NLNoNicX6MDBMbFfdrZ6h1H0q/zBwvjyfFG6u93T0l0/Pzv3ypO
hqSgsVWnPu/cPiz5FBtGffDy2Yrp10ZNZ3p/oWA3aAs3+6YMDNQ6xLyqkqqqQorNnDJbyUamCKFe
QZeE8ycuD/p2CHwG9+ZrbIzFXCiNqRxGOd0PAJ5Q4Lp8Fz8Y3UlWuowUlbW3+Rijlu15Iy0D7kJD
sSw6amRY1WzEb6WD0rmBzMtQ+N8nqAYva2YATyTzegWz/BV+geBLWkmTyI+9ZcL+a9Mfj8IDZ++7
ULcM9GwAt/h1RLIjJ9zeNI7ziMw7jY2dyyRQK5ZwzNCbZ65wlGBovOF6XqR6e2EqPFeTOYkF89Eh
2XcJT7NT7FUGi8tBMTteAhxqDMsZi9V7jZAzIC5VSg4ymFTXQ9UfqIVF65yEehHREl7WQIxoobE3
GlWIK43XMUHxfhU3Rd5VonUv1kPyg/PlHRG5zUONDLqrB0Q+hf42NeFL68hViVrmf0NOVUy0UTTj
Zk+fIMiW/khaFB6HhJ+hLvr+M3fd/+mz/Y6M9eJEPa3BkzBGuybIDj9i6zt6WFNBYayalh+NYX/l
Te+CXTnn5qkTgzW0dhf006xSBum0yKLxmNeJ6BBu/v4ji8Ff+ZnvI/QISo89OiVL8EH5cSJvTDYN
DOvYacGEyrLIDHZQd0SHZQSwe1yWuYcKvavu+/dJjr9WKCbwLjbdwagcB6PFL4Nk7Lil2jPAHKQQ
ZU3AikGI4Zob02NTQ1zG6gIasG5sANq5wFNXI3SuFz0olPj4hUJD1iXe5b+qipTucK03qURCrCpE
En5e4PvlZBjjijVocL5AsUL2ufm916elIKWFioDLTq5p/7LTfOnaFyjtYGWwCRuiCpGb8sRr+yDh
cicOXXF1mdGeYssU8zNsCWd4wM4ckjdrPxNavVTOl5fBTLBwQWZ+tOlgs06cwKZXa2dt5WhdmIdh
9OgF1EfI8vSWvo/iv65FL1NVN31HuJlAghe5QFY4iqRTmcEJYNuOkFKGs8zEnbb22VrRxtv1jGv3
/qNWjK2IgwiCwE+rvl7d9pFLfTcguFDKKLeRevAucffG4l7Oj/ALaXBtaz1KURa72markp9U9oIr
1vNsdTCiq5J8uvs2uHtQC2qFzOLr0RjK4mkoAI3mXzy3OhXceaepkNrJxLUkYcvxX6+SUakPMGdN
ePRvAENKW+7PKHzs9HDYk+rfgPLE40pPmmkkdlE5O5k12otf7MKk5tKOeEp1eig739cISwfGRWDc
lS51pJ+rd8r+dzgjcpbBK4HRZzS7vx2ZJK42YVwpCLNuGjnP8P0ktV0tGwmOtX+RQkCZwjlA81IL
c7GLfEMf6pdo4AK8UPC+FMUGJ+ColoGHdPX993a/em5xfAId0MkQRbo47w5k5duVHpI2Hzl5Qvbo
OsUc8z/BfzpATo6r3QV1yQlYFHcnNzPjbyHOWi6gIeLjg9rcrUiAtg7pzJDh6AClMthjs6XdEeSS
TZK+UVaU+GCR2IlqRGeg0pZK1fpmkQ0l353W1hkaQXIdWwJBk7TfruGLqYcZ4hk4WsyUmzUjXL6u
XSgqNTsdGdRpqUd8mMa3SjnggerzM8KpLiYAn66F9nLxaEgYTFCUcSkhgAlHU08TitX9A+o5Sqrd
JamqgiVW6IVtiT1VTnbkCY1n2DGd2Av4HNorTCp7WJDrwaEPx7rQXMg9i98M6Ifa1f5ilWKPfIRM
SA9EBKu6Iiie/9Otk3vCyHwVaEEj4o4ToJZKha1ps/DzNLh5kzh+jpYFceLxpBJ0NkMs1r4+cDGp
a6xSQt+a4cCAZL8zcPJRCcG7wZEK8cXLDIPQeHK8qiOBgVYVb+tVtVZAPmH7+lWd9Eg6njO/5543
NclkMDqypk3ioqW8F+YFmw0HsLxWIxk2zWZhkkSPTNiEEeoQyy7cgBa5TDYPdy+F6Ih2W56ZcNCQ
0MNzuPLiUoaLa1j3bnV41B4NR75RO1mjenrdfxggMgc36+edBtUE+31eCv1KZDSD9/tJUff3qy0p
4IwdUcZuiDgddDQk/8ja63a5fKI3L1kfPcjdZ9v2Emm3i0PGQUm6MtThDAmCKhiBL7qs0JovmoPu
1k0L/oUiD6Dy9gSAUjbOSlBCtKMIVzlzZ/P+3a/HDdAvN2icDvncSPN5wTFyxYJKD7fglZDIhVH9
mYeaHghqet+lbcG/iFRcQOlI0+hGaFa76oFobuDkZLi+kmJ8XWVLwDO1xAOmWlH/30gFWOBVw4NF
FSNroj+6zfR2DBP0/58/EMRHZB0JEvWPNOnQcr3vgc31Zl1eK6EH1vjvK97pzagKjeW4Gjed5Q/w
T+RQ1yw93TLs/kXPAI+0HyoKVyl91tCxLZTZmbcs24kPBRoNFqwe8dbAGUuz1aT+ZXlpWCid8lOv
VpCc5BiEIKy9+ZIK6sbzSqtdGFCYPZx3c3hPjoX9Q85CRH3y0p9FHKYLZ7NWWjGmb8uLRuU8KX8t
yS2rUWgmE0eW6EbztuHciHnkSc1PL7yYtHaEsBqSDaGeqv6m07oo3X1S5ctermGOQHRr5TZgvUxh
3UCSuNOZ1tD2rqiFnNA/3JyKJGGSd1WBm1y6LkIQqUbjqWzjUrXtTT54ZYnP3nEsooUkfo32UdjC
EI6hqn5QkobgkBG9Av9fmsQLDYz867LkHJAEZkBWUlD1KdNz8T2s1EtT1vklOVr0Q9czHTYcTuO9
3jUuy67q0uxIjcblBI6fndSmhSuLImexaIGNhsYDtUNwKYdf+ErhyM6wPWPQGr8o/5W1epi1fst8
PwBPE+WCTR9ACOQWZGl1/VXA74NBPROkpP6NnGNHCSoM0lX0PIVmmESyRBXMh3Rx63xddRqOxSOb
KIBAIUi8ugqYz4iuAeY14JaOzA4pBXjPHLF8mysFYwoAFGGOBVmNpQ2fx7SZjVq44bYiDfcSzoRT
fc4mWZYxt7CVWatfD/4Qz9+C/8YHNUNFlmu3aGuQw0X95MLTJCsIAxXIanKuyDfMIBwGzboPLv0Q
XGMniTt3bsd5Quh4gXvCF6K+Odx91ZfD1WzZ+deRSbg3S+r/OQaHBZ/AyS3nyny8DkkmZUnLIQw/
zHaEpdCHxKn3Ad0294d1vgRJyNtxUElXERXSAn7bTsTjdRlCzQ5zpfClHRJssmJee4aLUVr67EeU
bZY0tdEAvWgoqYuFViAo1/cKhxJfjTucU1/RBX4AcSuZs1oZcO0a/5fIRsi8g8+vTedqD74Ty+s8
oWt9p9PJ1IU008tQIRFNWn7RCwVtyp4p7EQM6hlbX3JrUQzJOLihFGqbrV7OGXIlUwH+ZyxE/U4T
0H4q55hMkQm/JqkdvnaHBNG6NpJixG62GEwKHTXtl5UXU5/CRvz1FcMGbEab/ghU0vyHR1dY0UFJ
Oxi7Y5S6ULPdnkzQu5UjCrGFxbvHktYki6zOJ/w/anUCoJ2hn3M+gZ1IrYYeZcMTuO/eAJMGBldx
Ont1yGiXZYpCdTJC0VeMx24qplMq+O21GOa/HUVHKxrz2Gi5tEDoX4JmwfnXNzdkoBcJutg2rqQ6
hQpoK2pTbtJRLFEv+uZQSbEysGeXayl18d+7KjrbXqqnendZpkix7qsBhTC88PHYclzxvpQig7dP
6Swq6d+or35CwnlfggavcF4l96bf+LFUE0TxUQshIYoddPKODlnXurim7/p1Mf+pVy76xM19EZtV
Uaz7JBYhjn196pXG4G0EshDzEkV+ZuH56+WiQbdpQU2+wGEUIl0rQqA1/hsxgvsYzS95eyG/MIig
0ZxYl7UPhNhQSDxw1DVMBP81nk4uZV1NV2cxAosWxkgwu+VtgTyPydToDoNSs0daLrty5vb/hiBF
oUUeQ2WeyV+OMOEkLiq79Ww4W+zyCMwz3MDCxu+LccSZV9EsJqHRm/7rhOUkh6FSpEH/yilgMmtf
GnLbHDPEswDZERTN+uaTCYHvbnkUxkKagB3nSvubjxc1N09q6NOBz+wkaqBrtrYutAKsLNbAuWTm
K2ok1FwXz9qgaxq69pwli1PQs9QiyG4LWu/yzntpgYLZFXvQ1WxWmcawxl7NtnCR1g7v5kS21cmE
Q7pI+ztgBwWVpZ4hKyElde1b0x5q1jy/iRZE5ccO9Ym7pu2KHBVvap6yKmQ5ld1bcVpBJ5uV6Boe
1G2ZbEEOgG9V97sGakyzdVCCB+q1jiJsD2tIW/LsUyjKpo0XaSiqs2WK2WIAjgfUwXFedjXLz7MA
qqiDQUE6P6CWKEV2bqKFVGA8tcR0+UElQ3EcxafQw9nyYf6Dox1P4zZjPSf7y+LT+cU8d3Wcfi3R
SuceYx2rRbSXcfIGGodxteIYPyi+8+U+vlQLX17XEW0jeCBpMXcRjz0+oAzB6sULo5hyWNGbj1EW
x11T4XXcRLNZ5ltVEHKL7i/S3xj1XISIyr4Djw2960nrHAt9OitKeQRu4Ve/rtKq7y9+Suz8AGF1
mxL3pZjF88vhFuLZEBhu9xjgbh1OUXNtFllKRmLgy75TLQu3/Sj783MXn/DN/Pd8YvznEHrTPQ+Q
XbghUjXmuj7PXzTMiWKvGuTl6tzedtgNs3yXIItdjqhZ709tHs5AMq5xW9zazNlrUA1/+SsMU92t
jTSVOUKIQNV9tKchSFZbKhVmcPlUTcx2FIvc14vPQLzEnrXi4h0VEfZp756nq6al9S7zS4ekMP4s
ENamg7ItlWXCjPfzIVlri7Nz2QV9i8ndd2teefMm2U86ktwG0RRCLXoCQCsTE2/8Yhog+CD16Mo6
G5dNoTLg5DYeIXHJlYRwie8LsBcwfXFuN2VXuXMIu28ZTgVzRAMKeN/7C7pEs+jSoAC0dCS9cziX
BOh3dxC+kLuXoZ8Nt++XNbnyqxpZx+UAqgxK55r+AV2JtHnG3qFKRY/JukCB317X2WxgIFv3JQjd
GD0L3Qog8oufF8dC4zBlcnEPalnFdxVDpfjXXEZ2dIo/1/kG7plqK0Ca3mkiJiZ5OyMf+zsYZwW5
fp1WBgqiBrS7lTxOOpxZSaLCvnnnJjb6hEAzB81063I/WN9VO6d3SyBOWc6ss/Pk756+9xKtJQdQ
HgGMzWvDEvr5xKPYRsQqohI1Y8Vjs/hGLDEbLhdiotkdlSi4+VOQqdmjpL0S/ASxUfohJjvvYdbM
vCHpFY0c+BDGU9hR3l7D/azJVbg1V2LZW+bmORGT6TiQE+3GPDkyM9CUVl6iQmnJqftqXjbGdeaT
WOKEYhjfUCUVAke+30216DZjMlTMPiNmNtoB8e2jKxnOc680Ie4dR1azQlTYx5ErSPQFcXffakdP
2k1m6H1WfIPpS6KPp93tKy2aargwT02k8PMLXhhN+VfYLzESqoRMXBntArmpMuFrfnmtsHvGPHaa
z6aMxvdhb1xaNqVpvKmkZx5zcznEQvwWgd3b0BPSg7AdScYleFcv0xEkWtBswzLMx7scvesz16WM
hU/xPDers6Y4hFxFNVRO9OlECBNrChEsz4CS5Gwu78oohot5AY3PXuCfGgo0KJMmaF7wWs99etuJ
5hRy6ripkVwdYZu92GtoTUfbZnwoOheGBshBmfB4fzpArJ2ti2DbMJkec1sIfaKny7MQDJafTjnF
yTgRyzBjWa4Yg9mkos2caxJlYnBqIC3I1keVGe5+tBgYmt5tFOZ/mUVYSKQMZXWvnS4v9tbTUzFk
37hoINN7ofJvE1pU+6jlPulMJctaG5h1V8DzGKZJ2wkrBXz7ZLGy14OL8tzNtPiZM6Wk4kD9rMR6
SN43r3d2Pq/CYoreYOkm9VCxAPClVf7a1ENAtXD/tVkU6Kht9UK408zHvoPwZG9UFmccErXq33oV
COvqkGc6PTAWDlgX3DtIDD3JqR2ecjp3rRlwhb8PN27sjFWCZ2AKXfOe8TZNZUsVB87AGavVQPPk
1ffbIUiBDZMZ0fiGFCywiAul8vWLqGCY/whLIKs35tdSTKGMfDtutOLHLT/Ak3JxVK+Qzv04sMUC
LlrpcPkCywXRFCoNkpqj8EyJFogI3Wy+7zi1GI6LLUq3tEskxkNuVnU75kC8cApS1MPcWzLxCy6B
/QZWRhynVmGUta9OAIrKLsvbwi3ykderF6JaHpzLRMjEsDPADi5N0LCp05MeGiD0w4Fq7V6cGgHW
V6dodwS0J1eMx9FdMb1qQHhUmwEJRsM2AeOuEJTRbVhuQe0z8wMj80GDEq43md36aiCH5UmQ4Nh9
0vJ1h4EMJE3Bk4QOPeM0KMYg1PLAfrko7Nw4qBmYAdxRwKcUixrxlh53KOxkkVw0V/bucdg0eLOh
tLENyQ6wDwVCdlQ/LrhSjDNdvNe5vn1iT3ShzJmAOlNYh5wFt5pk7zPBhoj/c/kpxJISStKWurw4
jSakBOQbLpkh/gwSonqtcfBes4NLTHNYX4P+Ch9uiS04ogo8fswHdF5PUE9nwngREkvemb8wP3tx
5Y2Uo1bySnGJuRZxYK7+YDaqGbXUWMPW7EIDLmqzQmZolYgmXGayKaiaG/PavnWW6HSwDP2hjOX6
mV3P7Ral5cqZaiz0sc7+U9RCAae+xVAjVZUyv49a05JaWxYVnDYfY5dG6UMguiaVjwqJdxfv/6/g
Cja9cAQ9uvGNlW3lIBI32DVgYnZWwIsM0Q5NkeB62kC8UoPPRK+Nl7THrLNb6AJJwfbr18TA3Lm1
qmnvA1ugPnpNuEEQz7Q5HtZ4tYfjzpPwpek490GS/p9ZnL6CatjUEXIS7JAZf/4gg3+TeB8tkTOS
3Xenfhndg+McJMWoDNFbd9KInYtlaeMogskzDyla34OwEIXLlcKFoxcu8UJT2oakd0Z/OWmXvhoJ
yROugXy68ve9ZKzCwUSSOPH1RihAsgnEks8wJ7hK+RhdY1+yXM9fBBsPbIe+VEsqbSCJ+xRguW6n
nfYOuWwsvkO0yjHNY+DJjrbeKaEeOf93oXYCNk07SV2aou0Z7OtibM/+zAsxKYcWeyzU1YjpvbcL
PqwvD3pPvNVw5m2uXKBtgscouzzMB4rqWcG6Ozuah+msN4ipdvrTQR2dgaPsNbck70ldz30ZVlmt
f2kWSPq3EcCFIPQ41P+PM/eU90Y/xFv2JAvmHojtiBgFEQoN5uCuCTEQjN511ciu8v6wVdsTU+Y5
la5yah4JvDXXRDOQf/m0NVxNISRtlJEpuVHDENkM4KW65EC6j/2vWV8g7SymM44vjKqKTBZJ+fLw
n2k0SbtxDpSVKHPqDJuCMesQE0D+ES+KF8+butSJGoQOuRyx+9PhZBHWE8E9OqvfJF9Q5a+RrvCb
hOfZbqafKNevbZbQ30rqmD+L5xbXWcuVt7VfD/CR01b44Wc5sGuE5WN3IZxSBZfZ3daSe6dHYluE
nSz0+q5bs9RaTb3wLIMfkVWO/D4EaicWcJZBnvv/QDXtcaYyT4YBVckc3/eG07QJQqA273hzFvdb
aGod72jSSeetwpUySVjnRlhKZuph8+qkCie2im+kObs3bIkM2WgfE4Yunl72KdTRd4VhBWc6lHIF
vUBKi9x3ShiCdePrsXsECXT7uma377D7+rDTot1m0mPmhL92zSlz3AevvsI5+XgwlCBbOJujZNna
wOtd1n2TIN9TCKTOhBp0LhJWuPJz6NGW1uIHrPqCz2sImObfcgnoecvbOlvjfJoaOwMURek9WgLY
5Xv0rdOufYkV4MIsLPeQsfxO8wmQHsC1Ed5g1/GKC+b19cue9T/pR+diEhnEi3rQwwlNgLvXBfxe
Z+Kav7dd0VQ8V4jOvTVpM+uxYtHzb797mhfdT89hAaeCbMoo2w85unLSeG/drvI95i0jy+8mes6L
hJD43tqaJTb7BmbqlurKLf4NnUT3c7nflXXdeu8YN6RwxG0HVUzUd7NCDJjt9YIgRcYcQ74s9n01
XO45gKtzsIITUMxel0Y1Bardld9g9v6DNyQam8ezaAe0WA1UixLD/YWvdzWw+17DwkZPFOCC2VE1
EXANQX8HfHPV5H3TD5KSF3vVAVW++KMPNLszNhmcdSN9HclJ5dnE/gSj4dJWZA+otyIupuNgwqcz
1y/1isKG8h0qQsTo+9enPMC6O9vFmNV8GUZ3OjoPQVc/ogfq55/tF4gjBaMtLFVmRRXb5wAswZuv
fcmT2wXvUkHbDRoT+lbMyiiJnSDkhzcr4iY5PV8B7PH+9wpPmrby0LImrX6h3RVjlPx74FmZ5Zjs
UOpASgNB1cpj/636lVyTmrCJGqjduEQxl7/Oig5NFXarP9R6jrU0ELl2bFYBWjomi7UBhYp04aLi
b8JAURnXgPFQ7Z4L5jspOfWFDeEduwwan8Q4bMweO8T0IhDjZkvOFPoyhxuwS6c6mMYLLvN9X2Ja
s1qYA6gcpgnC1d1UpWB0G6cTu1q6IHdcLAd3wQkv6Pi8ZbW261AZDfgPKD1pXLWNuFjetW/ghUiG
Z8dJV62kbiX3dXP9NBG6IHPiX9bn9lAsgHuJsEHvTKsw8ausOihFw6R79YIRk+iaoUA9d8z+dswF
880Bp4Sk1eeuD66ajNopogGVSQ10DxImh8aQZJNobssaCuXL+r5AoUwp5s4zRcIUIwZeBMLK5DU0
wIX3pvyhaTZLv50xyEDRXILW3Sm0KAjtOlcFCmyMh6sqDKGnU7rqiyfy8i6qC2eoxvffF109r1ee
BaVdyhNvl2hWmkzHUndKf4gJQ9sI/TYxMXRi7+FJeLPNBRLj+XsKQ35fN2jA6XV+ITyeOl32VBTK
Hi7vsDRec+JMkmP+0cJ4oyzfROH9WRQkF3thl+YzhL717vWyOT87jHNyyVOEvC1LsYDKDinuMQX6
whEfLzSMF1BFxsxfcCOUpJszDXZkOzJwIvICvOIyYfgSm3+v6HebJFzDNMyCTtPXzkDxl+7HFQ1W
6U259gz7zkN2pXJ7It/uwIP5MqihFSCAFPbV/YDRXEEkImxJ3dnWA4aUnuWCGLILVm6X/n3xhTtR
IpzBUQaM6qNqJhLIZy2YtWUQU6xXU7Ll9vE/5bNfUDl4gBqrDVPFfDgy48F6TnE4DPDcFmwn7ols
SntPyd/w/RsDDEljgh5v3Q6n0KhDDlYax/z7wWjqDXrYKQ67bbF70ozP2HuP0y2E68kZwX2jRgzF
FWNcSYew3/xWq58fYFFF1aEBpwj7OQEsmoV83XASyfSrRrRjKfSpO96ynHpn7nrL+8PeM1xbqtbY
28dlWPe2HsQ3Cq2CGBB1HfQu7p898B2NzXr+9NC0eI73sChigkY/3D0QYn5Qwq2BzXaQGesx9Mn4
XHrolwetijxz34sOo5Mz2fQFx/PvtCKBldhd2x/y/ilqBZVPJrbviVxDbYnH7fPOBgxpV0plt11S
oEj2qb/gZI/EH+hcQ15pkYSx9eNSsQizJP7oXUkjQEeHhG+BQnjyptg6NnuZFpupv7rOwI7et/DA
ss1Eg08g48F+Rk6iF5YyQLLe6MYRbI/Z11iBQsYgR9RRpGat+obMCA7E0OsvojNrOi4fIDN7BNTs
TPnBGPK0lGMEppthqkwXlfxRXDHOHftVMlVyzYJ7tJVNElfK13jO7E1/joVaSGa1CdgpWSSl4rbl
tTU4+orXq29kraM/AOi/zcZ72wCb/uKASlvb+50x565M0tsOnE19rHkQEN3SLLdiFHX6zdtGGapP
6sXsH1w4O9hUyHKzR3uzpfzEMsYIaDccNpC58o1RKRK6wm3II3kHsiHzFkx3yBmN6Shubi27KAiG
G7YhXxTochBhujbA9Q5PbMb1npmYn9405S5CWvlvPDQzL6d6Jpz1dNvqiO0XT2+ZoMgOUodFLJfn
v5jN1UVK3edB74WK9aA7Cm2LUbcz35uCwuMJC3PWD5zCzio+kfFVW8/SrdelJO0CiOfc4tSQ1VWC
eRHkKbZuoByO08DCRsAUDZOGC1yevUKM4RZWGzojcRWWGudA8zaEy31CZ1J01XhUljf7cBA55pyu
07Bv3HAjQoiJmCWl4E8V3tx5CBXQBOD+K9Irrtksai6C2Ce/xbOIuOnzhjjGP9s8YwIQlLGxJJaY
0LAviJjCUMgYN4UYkZHuHZM5dzHtWIjiZ9bIQxB+83fQZ4qU3RPlv/maS/7T1b3eS0iW4Dm6Pqfz
lBpMOBf+/RmALEISfgk+ZTnK35aB1xnshY8GtsQ3s14kjBKf+YpdpXNbbuv5ptMDR5tSksUB8yIo
QKSX3+LrfvGHFOLgYSWrqM1eZBB5jKI1IZQOQQxiszu/ZjoPEcfYCH26SkFVwhnSuMcCD+tS9qxT
SeRFbC6N7f5iRUkpw45muNH/A3VUPCGrTgbYtiwmQGa8VV2PD8QOWCwYRqNo3B4DFrnx//D5zbYa
jeyHzxzf/8EElmOFDX0vwqSRo+pwGSfxF7bm3B+lfyQJsEnaIcu4clABmnycEgWF3L60U/bWMxzQ
4UFoSlIkDqbQwDsra0+GhB4Iimcib82XboFWfDYohN31qkMWkKX0jidQSt0pMQ1R9yZaxj6x+0+w
KU36RT1t9qE8N2JAqB6rMTCaILs2RUElijXLTjcnj0OtpxDK+cJS2kZQn28552d3P4Q9iLWNx5ie
ZNajWnEwC8jAElbBjrbH3Y2Hp7Fwt5TeL30j6xfOdEuhjWQcGlMa+jXAD6HbnQHDzFVtRJ9J5cSN
Hn6LUwVph5WVLjXC2IsN4Jr7bzFO+gIEOxtLcGwGS7qqpG9kwHgNqU6V2IoLCHg6BV0Bkh+zTG2P
22n72NcqhBhX1xcj5Trgw9xL9QQFOwrgAtmPSoJVIc9ji/tC4AbgI9BfUWlLoteit3U+GoSO6kGY
l2X3vXjLgWEPzScxJH2h5DOEfuVLvSZ8BhI3GDZbCVl9DDBLRnqLvgQHVoZr3kKfHbN9nUY2867h
eaHZsEpLtoMssIx46E2batL4KNCVnW2AN8CkZcU3xoGJVm6qQgar/ni0JCYWCWzF3QOzzq9rm/cY
Pi2IwYUASVeBG6oGnysGcj+eJbhU0FH3q8GNgxFT+cxvkK+Uo3bwPrZ3dOyQc9Y/x2A+udC7iSA7
U7NJCsoOyySNa4gZRh6EfaexflRcZL2Ns58oLs1mm8OohrvNmDJB9pgbGpNI0CKBqDv6W6/QqX0n
P9jnrfzRAVcyC6hMUiCayfBL++Z7oT73OSJvK10/JYDGINV4xk7FQQDp82YKkj6a1Bee8O6jJGbk
sFutABYBOl0p2S1nYds5f8uvxt+g+7FN+5aVLBcrzqrM9XiOjzgOKCBbl1Ii8Vt5PqOFBMDNyzPG
75tM5HvDfwz/TWMtVCbPYUcQgPGejG/yP4+Z9S6ds1ofwfMXvs2cCttZY1Rp7nhlXFSje5duV5ie
T+OkW/JQgFvFFJ38YnlRVDOQDiiYdq7ajOl9fn2amwepZMW/IG9Mt2X2GSvArLhEaF6dWTuPQRiP
BtNXc9XkCHWd+xc2jt1r6elLICV8AfHSVewBsR1kvFq+If69Chn9WE4y4S/KkqQWpWA9QRpPhN2L
uIvFz8JH6zhpBg82/hloOV88qfF+ZKuSWIYWXGDUZk4/NUdKonjxg8LEK8szlaL6ZxDnkXBaJFpW
VAp4t+YaqU8b8LoGx5zFQjnQMCnUOgleXKgumQRIsBQBHcRk236V6PypPC3quZh7Ufo1UMzfJtwS
RXAbOHAzq4Jj3ok90XR8QLXdylh2+ZYE92AReq37EK0SDgi6XQPQ7O3O63BCiullOVK/CGYokk8i
8oAjjIZTd/SKqgyV9/HKQke4gU8OC1jQJLDN1OR8O4IA+F0fdjxqdCiyIOpvRij4P39ZrlmQ5bIA
aVygfpfQP3Fc6vCzZSJv6WGNrxY9mlfdi5QkjJqssnweFM65+E2rfGCTHicx48PFKzAgsEVnZpmx
y5jgzeLhyDWsK/beFb4/xZmy0ONXLLzP4vyHmnNkE59x+YUMR84CeqbLMgeYnPUSZa6VIjtBiXxz
O9Zx+8DP4gR+0kFxal904VYEN2VU/Kr+U6+BWm9zaeqgmR+Yy1npyVVICwUjVJFkg28qHikKsGr8
KO8DQA3MBcgo13ZVCvx2m4KCNDR493UN9ZIHFKVmLiNh/lUEf2EGZIWik1QbcpQhXb+kQRtkg9zZ
vnXaxQxZ2DfBVPtPBl02J/HRw04rQVGFt+F6/uNMIx8LS4J/yPHOHOjtJbh1mkMTHp6WBoaZN+G/
seyUmHnj6e9f8+EBZZaJTF5iRpEbQKBQde4TYJ5KEaEqwRvEdrRC6PUvpAq0UeEJQseI7zGy51/R
+V6rYo5Uig0XG0odKTmTapchxrSEKtRF0IgVrGyNjBfcoXJw5zbFXwKuL6ikJQkk7wRvxmlAuzwt
w+ykzJlk02Q6vCcklqKlZjoeaJUdoBebm+Lj1bjWMsLNP0ejONJNDnCEDSbtKPsEyJB11B33jlpI
HlFA7jXvL5j1h7gzHXAoPFbY1penhhzTVTbcvPk1tSSakicMdCAb89bRQD6P4dzkI8opW/UPxXNx
x3LLDUIjvm3sTffWwUiHhW8VNdctR5q0QAWFnfCcnYHqpLlLWv9npmDa+5i6Mx/GSMwM/fvjY1tA
qoanqadlYHpdvz2tY/j1oegXqU1ATHtc1ZtMzQtr2K7mb4b7tLaEbI4r0pC+IIW2/n5xa1dwqroO
dxk/9UJVdgOLw5qx700XVljuNlcibcaRMSPN9G8yms/aXvRr9fJ+VkJISIMO1bX8SpyI62Gyaedx
IUWk2Z0tSGWD52WL6BCs+w6td2oYBL7cCKi9Gkcd/NX3XNmN/9FRsUnewe8V5vcMJrq8GzCVWV/y
RTbPSi4J3n7EnoZG4HjTzsxWaipLleLuswlNuOT5l1AlQ92LuZmLQeuXi0+x+2ZiL/Ai1SBqLCZ2
iCrHuOuzPKMk+fOskFx9gwNDQJuuGNPwHi8bThVz0TkHNI5A3fjcFSOun9nuVz901cCzYiS8rUvz
+oM8/m0H/xCpWSbQnRzq0BPAYmtTpiQ1PiXyIHdLD1fiAgAAf3T4HP0yW0C0OSYyBY1Qs+o+Rfbp
3JJUJMxesu4X3Wmlc6q18MhWgmgzuHx8KY9xr39b5iWWbodE83zx4Fm3kSl64jDb1NTM6891c0iz
GAtkqwtxNbcLcgGgS0NQ8uh/4eNSyTy7QP8SDNSl45LWOKP9T/E/cBQjjKOvrtQ2mGq4j6MbZGGE
zzxeCw2QsXbSv72hruUw+55EOUYUioVX730F1zHm6TP86ELcHr4RtmgBViY0sCvSxoPd4AGtw6eF
uc/6lFpqMDC8AUwxmIF+oEGNkI+5fZCHnSJ+Y7U8QqtF2j8qZOJwCpOY1YOVNwxTytm2lBM+JNdR
FGO7e6riCAV7xHZnRTujhTHOMQinMk3BvGr2QK99M9AGeQ83cyYb1pU2Yw92sfrPLy+d6JyGSRdH
7nA5afO1aENpu+fkmJ9sg5CF2qAHhNd9VOHhINhIpCxHTm7hzr1YQE0Z0v+pp9VuDERhje2QBrpi
crBC14GHKbQmdkAU0UlmagI4AlcmhAYd4wClji36anVC7Hh2k4R4mLq9tzdcQcPmfsaFFLisXZDK
rGUWkN/uOI4wKH9dKzGSm96Jb4CEBiNhTLe9jEyg6Gu0HCyG/MNeGWI8SS9l30YKj8Yg732+sVv+
bbX3vTohmhUSbMTJlB0Rv5fKxKs/5nlP9+AvUBJszcAwOL+e9CfzNcsLoPO1hHYG7Allykaz1Te2
1s21RYymWJDMce7yZiMRoIAuZsDgrMnxyXpg9UpqM4ZKFNkWpotCfNMuoA2U+yoq8JFNkqBa+Ky5
5D6qPqB3LAkHHmjbGpvebAO4+bzt+i7rILdaRPEb80t6eepAp+TEy82nm6/MiF+P/OIuTALbU24O
o9NI9vT5xcDvrMnc7sg3zYyWurOnygJz0UlNqxF4+l6r3lMXWOS/jwWlb8E3+7od/4GBbN5s84ML
dnO1VUoQ5PxUd3az5lTx3r+W9V/x/AH+ubmfU0X+U69QTB+G1LkcIU4o0ZPSm6NnYR72+CKVB05i
m3eiwdJVOr1uFaGZKlw/vWmtzouN05JLGCAyV2DxeCNdMO5ZohvjJdKaPSF/CKM83BDJa8f70Jsk
etQFAW+aJAPDgeuuUhH8vljNu6nmgWc8XJ7Zd4On5VHZxIoK1EKEeUy3UvI0WZfNVhI2DNeVdOr/
OL0Py0F7xg5+YpuKVnFBUumJAfMrVegg7V2t3cIB64IlbAf197wZBl3nXij9hDnCNhth2qC7uTuJ
911NptbpmeF6dWLtm8Y0aFh8sP+zienf3MpalieBHczrb00wyGvmqN5Mo5s8UXTCg8FCDe6VMSZr
/xukiqZx3X7OAAPPeRjEoMG/SQlLMU7URNlYd9b5MH9QaVM9BpZL/dZr8+JID1gI+RdnH2U6fwh5
4Molbx5LKodait7OIzjSAtpgVIbHI1eUhUDnTxUTxWDO0kXNMQ25bCvpkXNIRxKghNvXjgKIFVhM
bK7d8xXg4dp69Nb2dGa3Rkq/U5xE4jDl943nANU6zLBmlQw+wbhPK07XqsphRrQ+AZwRNz1zfm2z
qqp2NM3Zk6Fg2nP0UisS7QKOkBW5QJ10KMGndD0v5QYhp3MsLrcOepSyhGu+Gd7T/sID674oM/ll
nWTlNNzPnuD4yw5y5wqyx0ZN32qHy0lVYMG7I+tBBZrLkiCaeU1S2fqQg7YjY2qVqo6YUUwx6NvS
pnAazjTL2TlWvfrKZ+3SSNC7KmEWQZidpsRucdpKVokAVJTo5+MJc50Br7qniZg0n57jeDb1wlB7
/4vRQiwXz9EZvPe/lDGIJYh/nuuet6JHJpyUesSTFPaQtXvZ17v0AXsvN0rJIwlFYfT4c5pdDcs5
1QezY6e/qsUrBUz+n6D9PN+gqO2gFnfW1/CDK6ZJQTEmgz2HDzWYz24Q1PJnAVd3MGWNfPAkl65v
ioBQB8RtxHaO5G9ESVX1MLGSYSVCFP3T4/QNPp5mZLdypsZ0Brpga34KVyfgwlG3rt4qnNlv21H6
CWPtx0CwdFZiJUAJndIoYnPHK0f+XDRgiWfPjgVU0M3cnJs/9ufH6SZz/beTE8huRPuQKGupf/2B
gfe9ZwxcBanSOzTZvlwV4kXrgs8JDZxG80V1EgX+Srnq4wAkuKyC67FP1xWyScQTfwuwkwo8u+OE
0eB9g+04Of19tdyzbwLDdL0aqAIDljN74Hwmi0r/NYtvZ4hlwM5Ekp26qnG7FndxepgZ5oRMGNv5
hsowPhtpVewMVLQZ8XNwXMl6uQrJ9orhFmVdxrMEtaFwz/oZtVkNxPOUOw5bUzmpbtgwLg1FAVRb
oFbZZYri/kzJOvhw7SLHOgqDtAfNzJIHQPm1t7rO8RpRM0QViazGxwiX5e0mK8S45HGKcVDF6BFh
0q28P4y6CPwI15RkRuTMbhy1Pi/XM66rlh+ZPgSEwveOXxRsRIqiccwmaYZ/TNXS3Zk1bux2QsTz
bMZX/ib4iqJgnV8igvgIkKsDcIomQEN5QTNBbYLvtyXzKfgfdbK1FSTJsDj0bMdUsqCMfsDqGXX4
1/Wko3rEXeIBiQubrpxDyGi+o0WrsaLUvNyEeqE08mH6DL8lUrajwnPdZAN/P5Kb/2tNDdTx2IPk
7+TPpl0syjtP7ayorWqpAHoWmFZlWgkRz6fDmDOnR6pWnmN5cssTnOyOlMp+Lp3Q4Txd3FVRvL3s
+V1gEd0pUsS0grBZ0VRZ+/GP2j3kgdrTNskpQ79qOhlNvYFxDm1LsShhHRefIxM8gZ1bIkGl0ZGc
sNbIfFn/elAAuYWsXJ6SnYR1owSVpJumCK9yWkDKLSvdm0ePxQgsCVKgSOa+WClLleixsxGyT3Cb
7mnuxJYfqo58v6vjiX2yZC6QvfJTPyvqLVP+c/YId6BZMG+Kvef9h29GNUBERXi3Chv+vqzxNb+a
uWIDYaKITll9sgAWj4lsB37lR6FkdVecgxlnDbxdn4wi2Jqn2gOyV0TklUE43lzkHjq8UabuMBG+
825QPd8KB8a/DOUSDwq3Vl2/3UbXI+uAozPV3Vw3+r2G13cR4t74ChwtPp5yFRcv+HC70mtGH6Qu
vRv3hTaMT0mN6FrvRPqbZ/GaIDPiSZnmfXjPFJQAvJJ9GOUHaHzBvdFlO/g6Xlly8bVkiSf8ioOS
Q5rJX8WvTdPfKnzHNznocYyX509QJfTVnM8mr9dvYsE4e3H6ZI1relw6Gp0NIYGqchMTcok02UpZ
icxVPW6ujzCrTAKGqWItib2uuLD1CA7aEW0VJiz3WeGM9toZSTE8lvuBIQ5PWPMkzj6HbFo02HZT
9ajWwG+5vdUybx07KRa4d5OS2EAKsmjrbQb06LT+yAlyd0nuWI4SNjmCEBy9QpZsf35hHasIY6bo
P0w3oIIgn4PDf3n8T5HFqljLDGv/n9kIL8XsOca2N/bOye4OZTGo5hPrx6UWaKjBUukPPGKKNtjG
02w+nRAW0bVYZmUK9kgz47HPtEexhzR14t9mg/WVHq8G2DS24CoLUhc12uCfG5ZRIhQLx33DlSyd
TzXOD7yx0RpDh6vQxBkf59YvLUtfMvslOQuG+keJ/q9rLNe2lEoMUqtJBAaUzqQN18YzkxXeG2Mn
ETuxOfk7NX1lx1cxMr+Yqew8+5WuC7cJqNm0IGG+RG2U0GfRvtrPs90mmW31WY/R4tLkMYZEqQSS
U6qrWmv8rYt5c6jirU1Ab7fjfdc5NIbH/cQuj8XUkXh9Tm94tKWB3PTTxN3sc0ejfAhOmUydnXw5
Ea2UwpqjK47/0h3TAdcVBb7lA2UqmJL9R1zgJeK4z8zH5iUfWFMkNSyK+0Mft4ei9vGl196k6Dl+
M0ndaXWD9xrD2wyFd4uiM5aI7orlHyZCDUU0lmNkOCAkh3EZCjAESu50Ade995strvu7/c4reCe+
uBM4Lll1uNsdHbfApE6hoVkR8GQH3lj6wJzFDqY+uqg8OWBeNVnq0lOnFcPk8Lh6y6DCsM1J83oi
CtQZ3UUfK23l/IeWTginNSCh+SyB6RQ0XF+HES+rV59pK/qeE3FjvRs1+XkRUf0UmbyS21XL6uud
rWmV8cLEnTiavHD4UXbFHFM7c5hr7Ry3QS9mfKR44Mhy6fEGlOIegF5TkucKF72Gq1GNXhX9JHi5
HCwBx0IFnDiPgvXg+EJiJqkh/RaoGI2hFKUdU4ptO+IkksthzhGpJThVGF9TFcurRkO0nlw5ZcKK
5DBorMZjZeRay2tJ0mWKggzJ6KINPnNRRakxeuD7Q9fPnFghls7gNvgzS0GcLQ8n43g0jleMEBi8
W5aDjVflLdipatCy42OjtYiNuXng7YYPlTdmQ1OFRFVPU9ME1skHppH1DO5EZCP9w2Rkh/duenO4
MubeiyHqQs3C91SxwYwxzeDW9Zkgs8q8/2iRAX7OB96StY8A2ghG0KS/oFSYpG2HJRcQHEEDun5M
1OtSXwzIsU/oEfdKe6WC9FBshwvM0CEym+tpskSXhMRRyvvJfebNxUCImFlTgMZ6Ng3UsEQZohoH
S2T65WFntStzoxWRZAixf6YW1QZwFgXO0oWTavwXmXlUUykkJkbWRczpOIwww7Nu2ms3oZSi4AIn
XK4UYUkpZQL7pX0/v8KLmsjOr8TI/hcEBTwHAuAOoSZ1IynX+6AHSFDfOt3GQSqRkGI2/WiDOJW+
eMMas/deltegj0JrSzJSWcB0R3ukhH5H+OWk/JHRgP6goGGQ0vyarhW//Fn86L2Sowa3qgqQWLUp
u1PMW/XRvKUNrfhBNJ1fKDqyvshueUBojmLurVwHTp+N80q+ex9bRwy/rnt7atgCoHl6x3xlyq1o
sK0FUJyNnQ9S/Bp0OTTNABszO6XYHLf2cPTJQWt6UgScEuGx3zDXVw2EtdSmnE0AsTFKTipDCFLD
38EBEStAT4UfEt0TV9Dj1wqxxJrHX2hJ2R6hpLM8pRS0rvBdxY+erTcWs2ed4L6cbzq1+UJEDOQx
op9HXg1Hg1419dMNp1wrYJlTWYJpcoAyiyFka/nUbWMz7dVXMg1UZDGZ4pkywfHQmSZuAT7wU/do
RumGsrHmfkY1j5Bq70dA2mSDwKpFpf6oES0EsFjkJH4MeH1fxX+27DaDTh5SsNrCj+ib/utOTnIk
u9rVBtVPphtZJ+95vFS1NIr9rNH1nzR03wCJ/7iVYaJwa3WkFAnsLiVDicps9U2MWQdhdnBbeO6h
/EbyB3zYALPRGAT/biFlh2g5dCYFU+Ko2nBxz6nxnjbLdCfsBvKhcbikkBWv8OogbJNouV+tDzxB
/nBtkzj6qwP2Uz/zwOagVmp0re/cq3gz9TZTT1Zryj24g+9DKQ37wFyYuXzv5dtMVF5Iq/RZkBhq
uVoPB5Kdb+bANetq4hMDRYE7z8AXPBAisG1VOrSataN51ry/1RVItB2w22VzJk38AGelDyfffr8j
AJoDNRHQw10H+728VjQy0ATfhP0HVhsbo5V/AShALdNsNPEwOI3x6kWVFleLBOKfTEmVf504X+/C
eq9sh/8dSUgZeNrfGHZkjpCSNnxrRSz9Cgy/MxfkBvZZy6MwNZPmTC19P1BuuoMtwg+xpWshnK0R
2uMWsruTxEOMnqnJarutd8EK2OIq/iD6DeRKTD6xKxZCrNnmq486ruLqOuRHgfD+ooUqEZlkcs3l
gqGVImsMHuza4zpMX4oNNLQohqN1qvZT91XjDxyY8a5G9YHfn3C1MgrJKDr8MxTTYbSBSjbfue5Y
KRpRNhJz76K9H7omXh3T9K38Oc3T/dBsHMOaOzURFtUA/CwzbLzDLnDpe+NDRB1dGD1IzNFBeKz8
UWsvuKghJIPeyD+y4q8/Yx/wmrzNThKBf3sgfVS332pgu9kTV1j5Sjhie1lmEf42dUJdz+Lo4XiE
nRUYkYOf1ub44SuXrT7f7Kq+2uH2+X6ZVp/AedZKqPt1+N4x4kBfFJ9eEzh1pk1wXs40hvY3Ij5o
ilklcvbqJ06QN+GZAIMPbGg8E3mAG6Qfw5yYplwWPxm9KbpmsZ6VZ78Q2twrRFZB3XRFJBgKR5gJ
6MPcJkD+RReSM7/PvdGTECF3XXAg2cwo8hhLDSWTaK/mYLmTGcWkYWCUSSwB4++lQCYPMCplF6/j
7Bh8/CHnBi95pqNwPB3MRS2pmwVHJchU6NO0rxtaV6Eq0E99qfHwytexqq6elYJNrDmPfqfuK/vd
mZiBmf+DPudZRzRT3e1bQ87vpyX5ffiFNe5ege4dk8yxz6L85x6u6UpBiaKUGVl1K52seF0h5eQm
P/FIDfR2elPTs1N92/T9y3mNYOWnzTYlhGSSTouyxPNGsXeTXB+Pynf4+SaEf19B3tBlcKKYPW9P
gwqYBTSazKchYX2+trHgmC97HBu5mdablCMB0Wt9X6eM3PgMEUOBeUDP2zOcOPMlvbkqy/SeY1Jc
9ANLNWX4rZ/sQDc0Rg7Sw//ikSgnvadVihslXrBKUpOwAnBpPsOOnA7GUWZUpa4FuJwkbUR1bGHP
joYfEhIGzjfUbrGo2H80zS2DkKHDaIxQIjNz4NsrT1vm8F33Dc0ynFZA6akE6Z9UFX+jEmhhElqE
ZPOqis0VTJTcyiC/5hEsA47mKpk3iQYXhO6/8pKIkl706+6hSwkTDAuBQGfBEVXIuXv7a+cnkchV
vUw+t+PFs7uLoq0iJ2ANxpO1VEgO/TPT5mIhTg+AYH6/sh6rZpfEH49dCpJhStfEo5jkiLK1Yewm
Whiwof/3c4fCXwxnMx4IsCeTsoYovFDZVdobptSi3ngXB3F9FCu97bKFtm4sUuRoPgXzUIgOPYqt
b8RrGIiw3DgD6gNDPrgqqThPlNunj7MuWW//L0Ef0Ed2DBiM2KA2UOFPP6kK/14LpNTjHrr2pldS
Vr5/Uf021R1t37xzJxsw+K+MHrG+VDTkntyz0anPD/X0XSi7PfNUyoP22EQYZ8Vc8EFGsO4nzdo/
x0+qyIscR4XWUY1AcN5x+vu9u4laH5iMhN4isRmnvKfZiyyWtOlOYlL+NR+PLOaP6wUChIncTHMw
gtW7Esyh0Pr/53zoW+kJPBucOer4uvUNUuErgM0bepFWXzcg6sth591L3BYUmDAluIzlsmRF3jug
v9iMr8vvSf/IDDEArq0IUVeM3YhGhpGuN6b9i8F5hdBj5rF74eb6S+O1bAz6Ot3P9rq5KHq7zH8k
SlJqCbnN4xYTJnCKixc6DtRSgMUaM03CC382BrBB8+xmJBNODvkiXm37wFZ06KVIOHLEtNIqEHSP
JFUhy5395FOGmxWluIZwWEO3bQ5lalbiDfZJRmXv8Vb3UrGlMYMWj5lIn6XVOhhrKt3ZOQo58Mfh
xEEHfr4g3KfvUdffObcrbyZjkQKUYGdFEnnVI18uffEpCmjpluBUVFORrCY4Kynn7Uk1eeqNNl2v
RUO//TZ3qrINUCE7dDEjL4sv5/HrV4uMSos/zpPTVGIh3Vi1rNJxy4fiirBg568AnSD45EcntTv9
lJdtmjvct6qfksBCXFe16fp9ZJzFRAVGRvt4NLG4PQdG5VAFALA9/x2Xs/vWSZX7E4K/yAuXg0wX
/+IjN+6nkhuagCqmQHWKv4kcPer0/hZm0x1pKPzT9jaZiFSFpNG1q6sncr8b0SJuCb8cCSnvMFEP
e6chCOa65XzNwsLbdxNez7n3diBlgvmBa23AR8g3b00hCliIyaVGjFHOHXw21WmkVg5Sx9L9WNz+
j0Xv1+TBFe47mLf1jjEDFPvNvF4qdl2v36UkfwC2J1G/QJkytne3voGZnh5I/ZFdS9xQFtUDK18k
AF1LBLDWXWFFwBFqKFzTl52h8EO2YRd8qYHN4ucnNTZwH76PQ+llw5VvflRJf1OFqtOiESClOueh
2sKYqxII1cukTaDPwBgi9jv4/7+0mYWQZe2/QzfoliEq5kzbDEr7oc8qNYivKhE/JD1I9Tu33r8+
raf6rl4UCONoU+QTZPYITZ77ydgGNFyacG6rtjEmzaRllBesza46XE4u0lRGex5UaXkJy7n8H/T5
cUhjZft3KnxmH5hBY9eZ1oYh1I83aBiAprLB74mLoQsEoXfRfQb8u44NsuCUjkzoUg+TtU+oKK4p
9N16aaUhpRKi52s0oiSnQbav61lMihol4BRxpLKYqwvagy1nJtxKM6VoPrjJUH+tpti1EUZM+/7e
4upJWY78x19dOGQ26ZvYuyG0wXBpnfhjQkX5/tvKq5vw1UTEI9jdELjdmsDEztkJQ1Ih7wxBP7qj
t4zrCWaZY0+EgVgD5ERA5b62NaXQ2PDHEa0INh7rQ1xJWwAloEyL1wVXu87j38T9IZNcKQ26cmNL
RHzuAbU+abGP6d6DOob2TJq1sqYsF/EYt0tURVhByz60GSloD7u1BNs4xzeniuxva3NLi3yklY77
iQfSvmFrwVACWTh5IlXiNzkr7hAYgrXmjnFT/wCQ/vMkHUDkX7KAZjvD88dgvli/Voro+lhQfoTJ
OuvESFL2BgyrEoaCQmfD/GphjzRiOUHy22i+s4Thcf2kBa4JidiavESCM+xyZBcqt2wA8lb+CzYB
hmVcLtlCY6kih6Qlebf9GMIZ7oQ7KFZPvQaTQDKhSJV8XytL1RR2g9e+UVpD2k1G8PVCVEOAG+6N
pPSOWH2RWaVd8Q2egNYCG0syiPR/ACAx9/+UbrDbu7ozPdtcb/I+bnD8PN/sfNxfEtyorFMMrS5c
MAo/LMfPNyzTFa3KV+4eKzz2he6Vvl2+veHpkG+CG1e2XDMhfQurxnmckZED+UdtYRyS25mRJ+WP
Ar/2gyFyLzilexv3YzKsTvWPDOweW2Jxs6f2Yd6xMJ3RjtqPtvk635T1cdTKHSPHtdhlrsDr4ERS
V/FWXG51mTsMBsdE9nrrAvv+RsP16FvTJFw17E+zzQhxMn2KN6fi8c/3kQVZc3+Tf1of1Bp80URt
HKmcEYeLQeUJK/wnrSR2tS92vtmx8qZWgpfqWAJ5M3CAQoA8X1OVUnT+nt7bPYiATIKSB80Pw7U6
zV6e7yh90pH/3D6z3D1nPvTWejkzOsQLTKrYaXaGjIP1nAlgoGBZWyQrXEVH8PhPImCNEQ/YbgO+
cE292SBK9bkjPPpWu48GZHAtYJEZ8n3+/fXaCW8pLs67YHHMYe0vQwBfQGe/zxkHz84aBOR7eqmd
Gayv7RFlqagmhaMn+NkvOJ71fMIy8XIv/eRh9HDuVF+aoOdsGMFwoCVNCq9JG928xrHCJ4Rlrja0
hh8gakJXDwICZVUJKMiXZQla+4eThsHF4PagfrFf9ojy9uQGehBkQp+rzbOzr72Nb7EPJHkzW/yB
Ik0D5TYwn+ATv1B5zbEbNZaExD6YCrlzQ3Wtze4wHIK49VP4l4+YNeDP/RCX+IOlm9pq/zmkogOu
djsMnEc3lbkGkKw+a8t5Emkgjh5HEdpBjM9IVO0f5iLv9efqrMtJE6PfbwNlTG6FtjWpzl38wAZg
cbLlJ/cejQfXsTPWttXCVE6mSYjj77iAWvRxy23BuUdao4q2MeICK4NlKSVZfaWQ16zJSFCJPpuz
GVtxegLhB955/AN7acOD864kNtkmJRcKqXRFYzKXd1Umaxr6CHvhJTgYkudlXwNQQY2F6MQLWxUO
KnoEipIpioh9prm/RzzjbHMyIZBtHwZMBNNwTdnFpXb8xG9PbGO4PLL7TqQSTKWJGyeQpCOU+dFf
YgcNEwyUJV5SZNCgOcLcDo9fiAfMF4es5+1E8Gva2vM3LPS2GlN+nnqfejWFwT9r4Ht7eP5e81GY
5ZqbmvvYmU7iD1itpTs0maf6CZaI2cXKru51vwd7CqVX5IrlPDT+zpTTV8ur7RK3ml0ExxoHkEEt
sMNu3gnI76iZxhC5Ogd8lsXprRYFBWLR5/4erxbyYFhuPqTKSdDgNFKb7iHTGySkSFeahx+1ZEtd
EJ7NOtqesxOegRvSUlKEW40bm8L3qg6atYefRo603Mljxrp9tNHHiAJyZaysMZE1FEacde+CpAv8
n/GrsZj76rvml5dTz8bivRgZwf2YgyGX7agDwFV0jvknhel/ZfZgWvpaZeDb8bmbUOFdctNdnr/Z
6mTnNvuMTuikF/JNbryA2zhRDOGZfmZKc8yJGouB4MotDYQ22qT1HX/QXklTLMGB7QU/V441fl/W
4TczJhXecIFBQGkhFOZ2C6xUF83UMS9bTleZ1C+wMbrhrnu8WIytNOU3rW7qiG0gY3hfBtTkkWsY
08nF74J74Xcjdbbz5MNDQxSd7uGpUnYRKjChnnyUh1/4+U/S7H1uKda04/GSKGAxmVwrjiAA5Bc5
q55ZIFeVwUq/CihEti0b7ccvBGcr6TkRWt2Z992B84VbwgxgrkrLSssereFcN6atMt6RExVK8kuW
dIW+DAb6CozVPO//AJGROhqIpphc6QUgBMK0jCLIFkFU8lNJ/Gd8asaJFHJ9s6H2B4uwRpzNIkNA
FLS1VhZfwRJFatZ9XRINf8ee0p87PLfw7kpGCISH0DLyXrT57fU3rRQ/7EPoXFG6gMWTYhnaPptk
n68bwL+hGH+Njmm9usqIuJn1hFRON9A5wsQPzw72AlV2RcYYLogsFDv2evG94Jvs9sb+Fhc/dD0p
eooAaCY8rpu2Pc0PQeTm9FX7+fIZMsD5figiU8IF37KpBlgKcHMb7oA+p7Q5Rm5DajlKl3jSnC2D
efSRuFRvt5NtG3pgI/sGkaxjQibxvN7gu89Y2mKEdni3Lxp1eOCF2Ii7tDFLfhyT+Ex0t1l93FeC
R9Rx45iL8defivBsHMdu5xi9GQNbFxfwz1ABH1VvgSb6bzRWZua59dlJGLWr8NuHUwi5vAX6eBd5
P3E0OOthciL2OgLcdpfAvhJFnJ1sAhwGKVMrRmTO8yU+wUsA8+oAThC9/9a7rgulPoxOmRBZrXxo
us99oHVGOj7d7RBBaen4PL5M6udvLyhAN+1as3hRHXTkj8R2PcNObWt2Aw/x5Yl3xbaCtslZgYDp
EW60K4utvrAjPSR+qtN6dLOJzHfdGyBdybTvpFqBqZ1AW22VxFtv2UE7XvtqrkwZj7Vo3aaAlXeH
XPE8Kc8QcXOlu3BJMWhqTTps1WPggaiwXK5vV72ot2j8QHum2AYfQPsBqtzlvCJkqI8wJ4s/+Jbr
XAgXpfORkD9CErV992lvTIg9gM4nQ41K4KSlGU0L3DDgKgg96VufYeI59A7/1MglDqkVG/cluN/E
gyAQ2gDbEKUrSSUe77f8Tnz4edj7C8Ao9KfMv0AexqIepj/7wYAKsplUHf7pJ949qAZ6Bw97qVhB
YhKueAZD/NMIT0zTdQ0Dp2cY2Mty08I0eSG/bp1oE92r6ZlDb7O/6wiPNWY6lyKsiLz2OSLltU9W
B5SmJpe74T0faRUSjE7UVhpJIZWhz31C2WEQiHR7CfXReEk+ltTdrUzJlgRqcP80by8UOcQRkhqv
KCPaiTOvX67ZUtI62V66g/w4TOib7PkM+HK+vNsY2zrR8eT6LU78zdBOG1D1FVeEB3EvvmYRYS6G
+/Ly1QuFd2luvyr1wuXVzzYR7C0N93GOtdp0+l13z9QMosekcV7BOjcdEBx2YhP0tPautThDt1Xx
hw+T19iBPVCKq90VDP9wyNiRTF6pRl367o1VHl1f1JTWcvMEqW+TK/Q+pSdXrdKuXMHJculp8/Tq
13xh+gYldYCdgNt4F9r015Cnz5FaE7371EHnKJqQXDlq6/mcqDg5ikM4B39iYzvyx6GYSx7ILgmj
5tXRQvG4qQ57qOriOF9m+4u4pKMmAYXfL+4C1jppIVp8tLG0wtuz6bvyJo7/76QB8KD+msI4PhHX
C3sbMyC1uLlYGswe49bAEowTT8Uwdd0oMLolOGdYO02FWbqS6WKdEZTBHXqvu5MVrKLEdh0UO/AH
9084ktsZHmha6Z64/A9DGpMXUx+19mhu4BSz5HHBRLIic3GU9TNX2CzpT6jFBFeYg4Ewbg4AtBzW
ztOffuMxiIXNRsxPbb7fyhzUAbIQWfUeP1dXbayGJ/Aat9n9VBpPmYzGgNlTckrR5xZJwXrlxq4B
jYZFBpyc5ExwiltF/8dJiTEFXhWyV60L+s6+2S1U3fJyGCwvq5dsK07+X3UtZtOLQRddM6ALvSMU
daZOhiN14mzTR0c1oZWtbyyo5bD0efneOu+jft4Sf2pdRURSF87IESJP6yJQVRn6if6GtLtNniq1
C7gLqWWe/dNxVrsN4g8eiUHsYsdVCLHQliB2OU5ogQCLgN8kAULgj6L/TX0kbxLHCHmczkYhPs7U
gdc3sMI9hJCucAFslFMUx2VhEYouMn0IIDt/yhZDpneZKExyCzF8hR0/p1KHh/uxrntWK9eEH7FU
NbXxnAIcbmJ0rE2ifXMIPWPiEyTbiQlBIaqzyKS0Hgm4m5gU5zEU5AzXwY9yrySsxuIEdaYW+yY3
YYYRhXmQaWma+SgjzYuz2GEYj0ncedeidsKWzaf7Fm8YzIK0aTMNmgEZMNyXVkv9UeHZrraTEB2S
QUIISZpHIYOA7aM6wGbOK7vy5MmJ0JEcFooJ2Dzk+p7t5XfNLGIiQNSKV7V9qPD35jw5q7Vo8OUD
0Uhe+d7/kn1i9D6mj/5F5L58uBbw79owP1eXQpP9EuIhPIPgiIoCC8b0Dn6j6CPKmEPuTcX9hADr
QmAR0YV/DNGnJWTtqAtwu0owvOvBR+nNCPf/lrLkzhD2ypK2V62Cjlj9ygKJJFEaucEDKdMdzMDW
IDaJ1GS+dwc9BwhhyzQU0vaZIx2BGlZ2OH0lgNwPuK/Sbb/AoXcn5OTj2/NW99d8xzgppi5nnhPm
1GiYSmZ6rTEQS6X8GNgTik+qEIc+XvcxEGoD5bb/iwXfu9BcVUlEFV48rHPc+NLhajY9st6TIQcD
kQcLOeiuwgGDJToHKWr1vdU3xsW4TJtTpkFVwuGJCqtbep+Y7pHeXQkVPD/N54+rUbjlGifcqjFh
PvbHOyecl4bEkcJJ2MDMHBICbtPQ4MrHX8LBLTYzfCpj/Afk5KpAnktxjq+Y4BW/foF+LJomhlmA
YmmVhIdxLi704kK7RSPFSp75PfX6iBtwgnG2lUcSxBQnRJCdJn4cc8UtsdmXCg8SM8/EhYJWtbV3
aU8LKqNm/T3lAVtukdGXxRI3oicmazyF9PN7EQe1u/KvdF8r/dmUh1/h4r0b4SrW1QWeysPshF1q
88aI7f4qJAq4BGcGUaZenFoVrX3tipXErT0AXXeDJq/8bzTU0tw9PKBKaYRq/bDHHO5KPm53VZEV
PhQy8isEV6ugpxE06KwJ/72d0TaTBHJ06jGxHCEH7Sx3F3adxZ6GtzVG86NjBZEuhLHupKdvJOpl
xDsM/Ft0EPHBJZUrQzNyjR+zmymT+0P3pbox2b/BzXT/rhmAYomNmDDKs2Yw+IymnXRpikOQB2qw
HrRfTIq807zHKQ1YSPJ3r2A7pTDhi/F6NDucLBBdjzlGdVbwzwhyqWoma7YcMTHecI84riU9e9M8
zdFQGLMRrsWfsGAT4bicudaReutvwUI5xLWs9vc7Nswozn4ZpUdUclGi58v5QmoBtFZgaa3StmBH
8R1NMQTEVrZ7POxOb2Zq8IPiCJiWy9QfZqupFrhF1BaKGtp4CD0wu0CIMJX6rclmD0VNs8mGUzxG
n4vQ9ohhKhWSP2FTESaTcc3g4OVnFIxQJpMIisVG2/koS/eG6PavVSifAnBdyS415GQsOwcB3s6X
F25IUa0MCQf2kZIqAv4/Q2nF9d07mb/0yeS3Pe+ps2Bs0E+FwTiHDpFI1Uy9KuPvGeQrNcSxOlfL
w7YUANbJYCMEC47R2L0x+AVlixNL0OkLx/4w5yI4zt02eKwCoBGBwG7wS8IH9nFrnBrG0gtaVrGB
71OxfQzeLKvEmQ1HovheyexSZ/OG8TBTIAFRlIqyGrKLsGLHhjs6IiBkNoxV+1FTwEgMSSRo857k
48BV0XsCGtRREgMs5xBjK9BAWG6HMObd6kAFizKpmQwG9aiejKKajHNsAyeXfBmolEZprq9VMOQ+
qi3l4966aKUwrvuZqkt6l8tuA32Qu16+JK94aGbgVKy0MMwlpyfpNRWL2sK0RdXD2XjLrQ7o7+0f
N3J9eFoGWTYRe+l2DbgFp6eNvvJOuYVWMC3s9+1pobjWkqj+VtfdkOkej/T2y/WtRa8cMB73mfHu
nVvIZDisND/TUelseX8mC4Y49XvhRbXiS/6cfYyLzWNTfyy7UxYQrvfKQcEywZecSc8AhtnfyFF/
VDY7qvisQRZzDoeSc8s4SCBBd++tK9lOezXartC7IALIsMRP29BJtaLsEJV9TBPQAyjUqsPqsmZI
yPtklxTu+r6bwNRiqpQfLSPRZyqUbCIPMO9G926gKLvKRgmQ/IImzDZsFoSXvIRkt7yys9swnyOM
m2TU2xEh005QVghHwBMj8+42XFXussrvVAf+tvLiezKW/4iPKVtuiufGc7Oe+UO13B1kKjl8FZE5
DDc3Z4pP4S/bUz5UkySmmXhbTe0kmXvbGSDNjlqFJCM8UFS8XHBtkLTnR8uoIP6MF81vQG+MHYxA
uewCh+F8eMEH8Kf5MSgtfDo9WmlR93vXyVeI8I+m9ojucdmUqDBtGXx3j3BUHEsRmboZciDPo8VX
wuy2Dn9c17ZPfS8XewrLhuzuoyqhbvQ5uaQl4KYskZTEnWur+7edR/kDw5Np1M8dlyeDkL7VWsNp
CA51GiiPq1QDEMQzjIOdPiDp1mGb7K+bpV7N1EtSrAX3PJ+QvYcM0bRV0imr9uQni4LsD8TPx1PK
s1Ib8J9u9aRK7Rjt7XZbLZc3DUInbkOVb6j+Z8hpHJB2CuW8gLEv1z7H3x8LMTgT2G7nsQPRJeBX
R4bX1VqyicDnMN25LgG2Gt6cilrvOAE0N2gmC0RiARnSWljYJplxTPNk0JuImJv5RJKEzVhRfP6j
iROz0Tvr3gdEqMwDLxUpZRxpidQlcYYBS5qpBrzkdBvu33M2H7L460LvUT8gxdIimeCmGHDZuylE
egeutOJ0vHjc1CjyQK/znpzILY4nqVWFOz/1C2Pk6rYHPn1SZJ1D8Y7p5ZqVw4PugOjSf8oCBYm7
TdoZpTE5tLzcQfC8L3HvFITO7PKqkeuhf7Kpk+f8K9nEoWMBZrv48nnBHLAI+4nPxb9RBlqk7aZB
2M/IfNC3mPERAXlkybB/xDxo7fROiqjCObm8cn6xu5YSWerJ2zDfs6ZluhBH5mp/mGsNqwrWP6CD
7syWdIF7W72glnL2gVLIOiaa9Aiy0SmdtOEj1EIQYYT8hWKXRVQJmvJaBc3OyBuW2YGZOH0WjEb7
9ewwZI52tkzRr6++qx9N8A25SuBoNdsxV4sXUeNRNroLZSWMA08JajAQYWjfCZeUIn/0XclF4H1G
D+R89D6idPn1WUaNIs/suP3YDb6iVrRXxf3ySg8+P3aLD70jkFCO1y+pYAZtMK2NFc6FJEpXoLAL
zKy8z63oJHmxcL6oM76ORFVfB3McqBOnrHT8AbXwDmpCc+4kgwgUvSU1F39HvCy3kQ/ixaShFLEl
PnZ+BN08l26DZnA7nBjuZqrt4tcnliaeX5sk7DiyJFjMgQ2pZ40jizvjR3UOe904ThdRFAf569uT
Z+sio13nzab1mVLy+jb2z8wf5lqFGZaCptabRxK3vGfY8Egg6k2Y/mAJ3zHoS5v7Mpl8A/Y+4TFc
FcEAK/Zrm62cIdcC0B0F+qn0Q9nlTlw+JzdSzEXX7DvTlXecsiLt4FNgvLpObveBBWQIwsJHXNfg
YDKbAgJphF+sS9YfGuLKvHDah3/frpnJfTfeRwzmat1lKuHx7/OX1paDMPMlmPxf4fvG8zpTO0bs
yC2fKoAbYvBScMR2SMTzLpmm4B+xunjX93rCjvce7jPLkPwoW3ufPRmFaajlMrcwcgeMaHeMOmhx
xeN1zAba5n6h+jBYo102JThDq7rlktYti6fA0MSLFhp5JdLfy316IlZvm8XIU5J0IGHUafPxhaPQ
V4mV+prTEsiaxLvTPuX1G/zUjGyYBCW8f2akP1gNot9nqWFsOKQ7WUfG+uSeNZ5cQLT92AEXJJPs
ctDF5W5sHCvNbCiXQEn0hNbQ64T4mApZlNlZoi6G2Mf7W4Jtm3L0ERM0krHolVFodyjOX5YJXd/O
odSHX6F070yw5B+B8gfRwOv7IGVNLZCxnW3ZZhdsL0Vu6pOLzf6l3ULpRQ6GkLwb8/zjTm7AY+2v
TWbmxhL+VBv9JRPKHyeoj3rhTTjWXZgE78dzrcQu2uVeiR1RBkUxx/DwocWC8j3oXeWBWpdj8iDm
8sfmGkU4JyH0IpyHIpuxDwMoMeFfT6cIJfKfAAVKHt1ZCGVAHXTmEj+bdjw/3PM5gNWHsZGnJtd6
n9IAWPKytGzzjDJ8zdzY+mG5FpkILoyspm0UILuZXdH9zv9si7pJQhSyklSM7YD8jkLglkm6Rm6W
u+dT0dcUqzWnkr4asiZimQWByM1N+/1Y/tc1OL5MXscaH6OFLFTJksd6wq+pwtKBgn3BwunqQj0n
2oI9DrHIoHXvrn5hGFwL+yNmHKj2sIb32HI3CSnmtiYirGMlLttvDWpOtiEmsQ64T9QE4s48uqs8
5XcrvG0UK69psOdpJ6UuQ/D1AduMj0lmZTEgOD1eOs09vULSZYeDieMCAtbMSsduY9JAoE2JMo/M
Gbmy7pHywKVltsXOKTxpKu2Dh2r/SE1TWFFkM/qxf7AKLyvDkdd4Knovx2di1y2Pt5bWqStfM3kc
WzjAMJFTW+CQAhLrSYSA4ZEWvLoM4QRj4oINThvwrn2yBu+gzJeyKoQyF+AqZo5m9UDEgli1pIJ6
42vz+bXFSqLjZP3IIMt2Euy2/f+CyEZA56G9SwjAcOtT3/YLIHmMWpLHvDhg9oYCN9n7pK2IcHdc
A4fYBfpM3fqAUHxSmgVWMuR4PYKK83cogbN94ygh0w/tdyYNjS3LlYXtX1LdXYeOy1ZvjVGzxA1X
nOWcchZzbBN9NaQvziyck8fNtdTC//qYZPN1g5f2tQ8ANjlFG7Ekawx6inTJWsNeNO01fXD5rSlj
yXWwa8puX7epnc4STB2jly0Pl8YZLMo0QECW2J8IHRcslCqknWeHxYVVSRxrm+3OEVr0H0kenFPM
CymSPdc/8m7EK2hD1/4nR1qVCPkAI8Ein/4QQbnh9KPh64HGB+N5t168sGQbAAh5a1YGAxU6J2Bg
98tjk2EW0MYz8u3qg9qf7HUYSB+cSZ0WBzQk1KdKyd5a1tN1Ow6CBmI0FBFS8qWqkSl6uYwLD7pe
+oox/T7vCCZGu0nBS77cl7XO1y6Mf0ddixqm3nYLA+/w/OvvLahJkF91fhGZhHujJOWgXuCmWrLz
fWIF3EyRb5RvxDo8z7DB358vx3r02LH3bJgT3f1xLKpwovEOFWaiTeXz4GpKkVAMpQPZvDHGAkD5
r25i0KV1pro9lgoBi3M1BExdAqOoBJJUBd736+haX8JjH36LHMNXaslrBOhKPnXMPsPPqiwZNkZz
GimrPNy8RbyHJ3fidUHSt1HsKdRHcX1LtPmyXjIwavW6wriWX6PoTLMUbM0Pf4dU7gMqpCZ99aLv
Juq4s3UiwQOGMC1acAQD/ZdpYevsVZcB0jOADAxGZEVSqHg5dXRm+oEmD2EXVmLBsBCyBKB3PFwf
MXDGl0GTyxvEi1jinCu7UYolxxm4cPt1TheqWjXtPL3HRDWWXIxj+d20JB006Lr6Zmv9UDyB+tGr
qTNjDdRmKbml0wnJfq0ONEqg1G+m044NOkJnJjkZrk57norXTqUHWstEuckuoJ/1VnBkpu95JpsM
DmJ+tbYqLtYLtmy0vDHog3wkA+JkMKtsyYlnK164dXMFr6WbtbA+4cE8w/rb6iMxr+/pq2b+e976
LpM6UwJ0Hut6mMIdSxeJ4bMnsjQTtKxcSpUyPzc5P3ecE6OyOIx369zAojGPHGUdKAgTpNKYBowE
KOM+fKYxVZGioxzg0107S6P4STm4RAn2dONnFsz8gLGsXLhl10dKjqcOtqMGZNedvK14n7qL13Sg
cGynyu5pt442vxZ/MSsCea1UBKm2IqfKx4y9FBPj0fqQSMPS0w+YWjIZ32CxFsIeeQm6QJUlsalV
+uNRgcV1TG6/tZ7MGGGsE6XMwaSAlkgZAjBN/cOGd+t4huFvEjIiN2Y+bmhWDNYoAnKj/o0ulOoo
v61YuUNFUU9PksuFl/cHCUwBuLcV9uPPBeUkZ4biumEeNI3yGj4LqhwVbDjzrmGjRpwZI7+jEkJg
j675N9wGlj6hqg9h273MhBKlxK5QgwyP+51Fg/FuM8WOETaQygkfEOcrOHjakJtpdmCt+fCScHBL
VoHzkezYfPNEvAjowXEPGGrrdjo1/3KLpJinH/X34NIAeLAd5jIsKFIgyM5LQFrTxntJcUXSagIC
+h5UZIZDJVVA+O6A8shQ2p6T4PEVf+Sp0f6YJF0BIoNG+D+zd44A967g0+aALDe1UyzYA3YAFVW/
OYDHdOfRq1GJ7vfnCJHXrp7FJm9xWSzGXL4yM9U9q+tWWHpP+YbjkY/z4aiLdiDt2OEC7SEMKIZo
b52k8pT/vi3IIXxjYpuAlnHbq7oOpyhMp9FvSptxejgQdw9N4+KL4BHDwYLlRLvRTXnAfAeQEb2Q
5ghMY1oug/f9y5CB7bmaVd8VF8wfRLhiE7OKHGVq9D9Yf7XmGVScUFlTbXhmsMB85i2Z2pK+wtuI
VfySH0AqQZQ78Xjxee+oegbXMWrczZzRKfEeyjqRCyC9gX8lhYTNzJkgqH1BUDiKpdPfZyY76YmU
Z+GYgvcUdRkzpbTZ4MzLSa3XSN1FuzNGz6mO8PZw0ZmPPnVPy1btfHyTeSLaxglGW/h0WJcGh4de
2+6MLQ+Wbi+Zd8l+BhaExibn29WhFPo/jYStZNh0w89cU+ExO1XLjMjWgAcyvY9NsiUjBiXew+Zc
VN/J7Cw+sclUKAiGiX4TVYfujCGT+RgVLMf8e2mml9lh1XhlOkB+ziSJTGPwbqgQMosPXWEhbcwG
48+P6Zr6XuCPxC1doF7+Bg3SyowS4noEOSK+LR7xdajb/dHEfZX7W3mYfkLNDuxsP0+j4SBM3CXT
DDYC58FIivL62KNzh2MpnpAYrf4mtH89NtDknNvqS85vQhecvgNYBrhAU4GQWEIl9YObo0GPWG1O
I6QizKfkQzjW+O812jCQyCCzbhJUDI0aGl4yo15I3CCRXZzSPqN0VRs1/8dzjCG7ASaG7DmxepYJ
xui81iOGAuFMuBdGqeDxwRFG77xhvapI2udJgZzoJ2xa9Lz9uGRDrs7wuTnFXrIdAcq66WSsHmUQ
ySf2MBC8ElV0IlwkPSPeFZ+CyG17fxvBrGfcn0UwS0V8anDS1+Bqp1t6ncOt5BZb8V/q10HMT5ft
qqo2oqLiP2JXkBOgMhEsX/IzEjzkRdEzCgGxbmTFMuufAL7fnNsEDG+6hivl7Q+q5ygzvdny1AlX
HG7swuXKKdaN9TwIIqrm/Qq4++yCbenXlVgCptvAm0/EwHBJUl+hyqlmjjO+dY16b1ztZfLOWnZt
KNVSMrXhmrm0y4BoYPRfYi6rIY8DZzrtW7JygoNMeQt2Ge1ZRe0OuKMKRyFWz4A1m56wWpjtVKmz
uEUD0/bqFPIkvXw5PT8tUMV8zTZn9AtfiLUW4MD4yHBYhmtYCKXQ/f/Xa+8CoRui+UWcR9PaHbSm
Hmj7CMlVZqLgdJgnj0joiXEqYaZGgN9dGCE2F/nXF3Y0YC6r2ps4v4wB1b2jlIEtFK3PQBBDHS3C
lXP2So8epC2bmQArDden8OYvht3Vec+GClUrpPtG3AtwNopn4awbOfqlBiXnI/fFhsomGdoWG78K
pT+tpfcsNVjrx4Su/6rEnLiN3vBTyMFj0jlMrbuYXpuMeZRsA7dbSS6eVJHJvX+VWkRSYU4SWHsF
ZNzYUQ5sO7eiYv+IX69/wzSGh3sSPV/RJX+KdyJkdhxCZHj3zwZVph4bryEgCXfwUhTaebwCchu9
2R2nTN/LcxyfQrpjYrkfYeMbQ2G77qXu+yHMwMfyVPrSh+ZiYMnzvwCzFxB+50kwjd4KriJVq5rG
FmFdvqKeiUljic1Q5YJ4Fht5vm+QH642IRitAQYbWOeYWesuSI/3YQM65hIFRKWcfvAIo9x7L+Mt
Lu7Qmb8GLWVN3NTsa+iOAgg8rkT9BOF20ZnAp37gy1MgqUrfW+1iVqv+3vcwkunvJroesBt0F1yt
5wSQJGCyMUp4ql9XiMbyN3Ca7vKEgnbZvIdTxKOGpi6p88BrfT6u1HEBK+KG/9ERdXD1xABCv7no
n8rjKPHRQNdiYuk0M4W2aV6qUS6f6wh5C+U6lAWwaCzx8268rZQBMEFVZd3vdfMbeyD3chqkUEHJ
GNC6Ah3rcYZXn9AGtWPeYeZd0xx+kddcwGciu6VnIdjogYZtLlZtjcvbcKiLFcmLJ5osy/OTZhfV
KlFUwV8nEgzIDmYQaboVgq8Nou5KrXEG4ZhKXAo8uLE4k+zxu9RI4e/WzVV7DO03tGA7n5hINoza
GQF0WPsoeQeMf0lFozxezEg5Q0T2sC9xELB+C+jh+B9q4IPIAN++LTCenCuONQ0pXvMbNbSSxzUL
Ds6wh5YOlMJrZPh0VBdYD8MkN0F/VNCz2NBAwTS9PuypvPCgKG6RD3VsvyMcm44iqqNGTAmGKg8E
Qtvu8LNDJ8tnB4hhCXfrAKjzfIckVYpsgJDbutOGdWIychOFR9qkDEpIDiAmB0D8hxSabR55orpZ
yecu0XDofoAsgzTXsUgj4WfeVOC8S6OGvbRMzvAA58j0I+L5/iKFZ2wNa8nsSMc4dsbnETNeV7OD
rrciFAdbRlckHFsdbwh77SZ0CUD1NnU4bmw8K+3YWPXcDdjUepuYXEfI1xZyczhlJorz2u/Hucaf
2ZOLOrb3Gfun++DHmJY+fd/1QP5QTcFYjjCLV5p9cDSwOjRdsUgAgb9bVDS0DO3ltGXYmNxbLWCK
WFeTWweVtvUKdZ2wDYOBf3Z9et6yDCmjANiKAw0XaB31Fa0+9LFhdLniigm4gNcZdVMcUi4O+6x1
xUQWBQCflCVsjHR23hMjnBqssOghSCo3XB4kaO2FiDsupEiYpVlbgZcSPxV50EhvaYChVcr9TxXu
8FKRp38ntzWbc48BlHRHi9yYxCrFVGEWdzfdy5XONJhg3jaTb2S3FnkZLTzAxwFapU87wr4EP2yk
b2dCuMfqL7rWJjnzft4EL+4FNkU7U1F8ZM67vjaz56g7PcA1+4tE0KmdnByMtakUDKp8q3oledAw
ku+60WKgqLhB+ViVsIeOeqiZ4FNKFni8mkQ8Arw840Bkf0uIEc4mFr6uaeSZk6ecPIksAafXc1Kc
Q/9HACoCJxawzZjB1vfTA4tsBxdxItCv9dWpU+KSCu2Z9GSK1Pk6aUwrAyUY0y8if4PrURM/oeG/
FWK8eQCZNekxjHUn1epTOw75jqFnNLiCmae4xOJwqXtzlUXMCpCuBm3L8J2tMtwAlQ0pARMVEqfL
6+m0Irkv+6qZ/yvemtz2xTAc/tG92TnNh58OwU+BR25hmvYsVVLI3LDVCkcAN5uYbSDHaVlyiwRV
9g9KCvfnQRjidE8LXs4bv/9Xr2ztSsD7BIDoLDbatSJ8Kx7Ijk/WrQoyNXPM6dco0/Dx9DSt2rpk
Krhr7fkFTWVGsGupPnuTlICv/C37/7Suiuw2Q1a3crFIZhpXgogLgnVvYkAE145EFdKFLiZNdjel
1Dbk4GL4RBE1Rf8pDnURTSjl0Lt7fEdxCbGp9n3O1nUHd4C9nRYaMBRfgloVFGVxDg1njqf7r0De
p3Rc2J4N9BMzie7L6kAfIGXCwYC7V2QcSqYj6tVYchWcPv4SE5gZYEnvUiurx2jpDbfLpaeYKiqh
obatXY5fCqR3LXSbUuCrNY/wXSaamLplepTQx0GwHOiT8l7Te6Kvey2Js8jG0QLXJwjYoKpRuXyn
PaZTnzY2ZMx7Wm4g/o2tsBAjq4tXvngwy0/8T0ePXM0V8AMMeh/3ncZieYtIa0+9Q1EgX0izuLO9
VKN9BqJNM8r8kr0VDIsxxkGUpJZv/vpza4xwUw6xFpjthg4Vz7IEjGCS/uAGlHVTjgty1UETVm5u
nTTrDf6Ry4NAfqLOrKUFGvvewlKpFVp6dk+XE3C4u3dZreuKMdwd5mH5hJdLHZlQ/6eWnc5xv/fs
SpXrKxzs2fjY5CyeS8TAJlaG1XiVcfvlmBJRf0kW2Hh4rDP5GuGkljvCB25eRY80DgqW0WVl1qsU
0wVIdOPbPC4mdt1zp6KBEX0wzZrqpJKex4+kkx2XlIY/Xx9VSyiwN+5K1qjm+cZhV8v1dYhjp87w
hU+On/iyr4S7tK9iVsVFv3IsD3GGbV3WHJssZlcd2JOXZIgwkCKPhnYN0C0WJ7NgCjhPxeFVdlSM
BDNP4AtLXDqbjK6SyAsycN0DUa6anyeUhwuSA3Q/6Q/OawKRDNgjVsYzfboyD5GWjqs4/HmRmUtB
XqL8JmMRWWtfGeaDolyVRm6uSk+gKRxpU9NX+1BF2pamYNEHRn6OAhdRtKqUF9Cv7+s+zXRMVy4y
ivHQ8Nq8IdXSvBP29xrfgLai++1lTrGyhU8+u94QYks3jKQ0Tpk/0wndGNJ0vlMvVXoUqkWlIc5J
hQ/2WPptnkft5HdpJcpQWdeOf9aNeFB2TRpmATCGlI9HWD2Q1d/Hk3xwixnVjx0rnbVDBejKQfLk
5k/YkiFNQ7qTtherETsUtfk0NbQdK28Oh2D219jAFa4nGK+C62frgd77XfRVIH515p3KM+z6r6lQ
k+EwonUcl0FfqQWx2O1DnT9O+01mocEqQkRNu4HohIrDvh9mjwNs0++ZWP3Jts8mZ6XUd6dAgbLt
IxjrGdzuQSW9qOvYI+HpAL2J/XhCsiClXsyO7dWC6JfPO8cc4TsqLU3DTTiBeCnFguIkfkyNFIAd
ALjj6hlMsZXdiA2BvirHxHT3UCo8OcsQVMJrldcguEQm0czEGvwl1G+p0TL2vLuHD1dMJW+2vdJf
zq9Gb76QqfUg+sm7UUqvIm/MYHgxX7MRRoHGMOxL8R4UB4cmMDorpNarjV1LTplDD0hWZg7L+Oyh
gpOVzEyMb4RMWDpcB7o0ZknLCrnTzc8+ZeX/g0nzwARkQpz60jio6DOb8LsmSl9UToKnDnx2M6pY
gpUbE2Bb2gk5pgWn5kAi/sS4pJftuWkWsd0iQIOKIwF9jlzhdQ/KwKnojQis32pTGqFfhZUbd7DH
djnusvydZouN7xOxvCpQaUquXV3M+bnIt2MqGBGZ4ngznaozdnS/VHLEl03FFjHSidOWKXQEfmBI
Ka98LxNQc8cZtG4oKpBJ0TMUjKueZZXV6HWogNyHQAebKuyOU4puSHMbiTpkmh02TEyaddHSgg8W
AgyuwzAqTpJb0MMd4o3JnPWBv9VVlzE0ErkrIcyWzoGvhECP44jkNvktvTPFjVVgji4t6fEKJ9bD
d8A17cTdmDZwczMHd4hoiUc5XPczGcXRuvyIuGvTV0ujpGwOzoz68mxM3vT3cj9zjwe6gda2loJq
O9sPRuL8lmfHs1FhVJbyWuDUInR6tYcj27mKlNoc8GfmRp853gAO4we/GsgMmEohGEMapNU4h715
cKh7GVzkkwA6BctJnTHl4hFZWGK/SBxXCsdz9CDHoKFlPtz7IDOa5+fJmDCf+taE0nNyY4kqaSit
v96/w7pW9Dnkar1AzGDEiWBIKOcPfYWxdAMTuKei7m3gG1I1L687VOQDFf18LsuBz+WxpFMfWMfv
St+hbeik6tiuSKjUf+CAZNsPmp2vHsQzu4TRCWCNiQqF8xvKl8ddXprGspV4Mxy3YJzgWLKXDpx3
ldbDLRbzg6tg0itUQDeUhQN6SsPllsGYLfHOCE2jMqvo81XHdLK03pAde1k6uTuJ0WVnXl0A3Hs4
CpGZUNka5CTKelspjV+0ByBAhTrMsxPL4DoOS9kj5Sj71N8QQfY0syR0PCOO+yktDmPSujKrck2O
gh2jJq4L99CB58yhu0UBQBCEfbDp3ZIH4G4cvokDZqXR9f8lZ78ryAyi4kAXP1VfnA0BhECbxH9P
uMKMd5P7DEkkl79Bb/bTEcZki5JsV2RVZvNQtzOZTi9AaNhyvcO7Pwb7JJ3J3rTetsoCFDM6PAKC
CmvzPOnCrC7HF1Gh4XuTnWAjHnmJEIrYgZ0GknqD89eTRFqyh3+Rr+lQjNs5jzm4QQGy5G7SmGyd
quET3UFwRHTdOYoQ5PHOS8m7OJ/MmMRoP+wA4XBLvDeADaVUgFU3Sm7s3G9m3zcfHa4UrMsN+Ez2
2dWVP4NIfcI/n4YSTK0S13WkJR1xje+nNT+lOJ9au+wsXYC/9m5E/LSu0pqJAr2h2AH2UeeV1Quc
UtgtRyC3vK7SngR1tvF9kS5mI9YD1Cdoronxkf/T6HfC//m+iFMJ3+sXjh4KTvWAeGxDcudpUOBm
wVuYCEvplgtce0551LMX+/jzUSD/xWFzIre/Yy6L9/h9llaHLa2GJ9MFEYr65TA3OGRcSsuXoH10
032iMn//1Vw2sPrQb3aWdJTqSRY1Xc/NTOq5MWf3Q+X9nsrEKuQsCL5++T/4bKvqmqB6zKz9IRQb
M9pzid53Kt3gB8EcLfEjzxEWHjnKZakVeynpJ05/HrB14vm8jtZMj7co6JTlorVoRl2Q9PFWqoyD
6xr/e6ekoh9d+L4prY0fHQ6J6Rv9IjcGt94ICX0nb8+i4231J9AkPE4jdaBZcqW5fK1LCN0iQ2BM
1GGV+/MSt0jVVQtPSwg3UDLCvzF9FjWyS7pmM3MMmQqsDZTH0XTtrTnGflMRX4wE9nb7YlIH6cpA
Ijencjk4Uw5fRoBGoYBM4YcxQihP7Vh4cYzrtRtY+IcwjQ0lk3KOKyrazrKhT5ajZSK2h1AmPyhM
tVQwWKBWW1rIdAoSvl1eju5UXVtthmY/ZhhraI8fDA7F6snVrh3llxUSuBx1Ce9Tk5F5PQxbDhj6
URRxxPNe8zU6URoaGfHVhdAyqRaS1rc6VHHeGs2ilsxDSfqrmMOvwDdZCtAKtwEuEwv1wWQ5/AqB
wAY4mthMjx52vVq1HW2UMu8jj0v2ak43vKZOpWidVJapYUq5r0ty1DeXbKnJAeg40Ru/kxaxrdOr
3JbNAlLuNPQYmA1KsQ8edzOl4cruuWVbMJFgfSLd0y3XMos9QdVr6G3ClmPTKlLMeXhmi3E5KWbJ
FZcMejd1Vv+Em9DNC8omy5xbjDHFvnF5fwMdWBHozuMr/l9ioJTS18/THYfexi4VedqjXMdBHNQW
4K4M+dXywbboTmSsG8tNDtDqIqyj3TseVNxvjuXBwACw9sFr1AEDoxF45kzgbpx+NvfO8bOfw0Xu
s3X5novM0c1EbRpzViuBsswQpPgUYl+G+iQFInpqzjFggsMCB/fkupMyU/Yh5mSSEfwtEX5NI6dd
msBk+SYWAI8hoe6Qjg0UIh8dwZ9zBQhNjwWM4r7gRwwFC0Nb6ZXkCnU6cPaGEJka+fkx7y+uPU4k
kCr8vI1afZpWKT3Xn8/UE/1C5fh+IGY4KL0XJuo+2eT+F7igApDuzFrEPagbffhNyrrgYZlvBE6m
tc0l+LmmHpmrzxgSfVZ4y/ChDFq3gsYUfRnIYv1eBbAQLgGn3DGKQ0Lv1rOmK7qxtAIamaqV+hUg
RVmkhCL+2JQSv5AcgXrAfNH0e5CSrm5qML4+7HqiHxF1LkZseqoz8GuGtLP3hCv0SVKBeKgWjKjS
3sogc6dA6GfWh8kZjH9bULv0+gMPezPS42MCK6uBF++s6F8EabZnMKZ9FSPBWw//Gv9aKSOOpv5T
Z2pWLp1YPrahR5QqixhYekGaWDj+q2Eti9DHX9BCFJUCVVjBaCMZROdgl/pBObpd+BP6fZ8QUPX5
VstmzTlRgwMabybM1KoDPOoZZsRzqluyWYpFKFOJ/YM6R917h+jH+HQuwEHMUmQchHsvtzSe1sh7
XrXmdYaCuTDIAZ+hYcQ7gBSUNnxtIEXvtSaenSj++0fkJzvsFP37mV44/I9lDbKzUUFC6g1VVC1g
4t1UMe7MuJToJwiR5TDD9DCn54aqnIBa3Lu77mXFiLyCj5RtCyuZqrR38SDD2+yEL+h04vy5E6xx
i2I6CVBko16jyNBwySDHSUsFupKLIbAxCQVNeophhqqDfu6USSXmlK5oNVmM7eOzYSvaiySbG/mJ
nnYvUc1SAjzcvf2YDP+6y4qJxyYfHF0A/T+676CQeCwPy4i0eho7P1eqyYGfKyUkHTC/NWRp33Ap
WssPaHGALu76R2vKPYjUPsNu+4eODw+2Qml7BagtvvvCbEYQA41fEBnbYWkbrxZCmvieyi0xvfkp
wFrE/09W8fZAV0IYmvMBUIOAb6BTUXlj9pdAQuGLxsHQmX+8gbAYLp4zNRjAzzvgxQgdVAvgsiHq
bIFFzd+658T1xDJ6nDPUGTIsoemOWI66nqixP25dj6wjosBcKgsw/Za8qq42fKw0HcWs/aiwTkz/
RWl8uyFCHUbYcab5MyyNqgQPKDZs+jhhpRYxPCeCxzjppGGZopI5hFJ3TDoDfz4aNRczpYE6mCPE
GcxtUD5bcftw65pMP3VpCJSG7/tGe1AyZaIU3f+nfeAP1q6fUUoNUhSZyhvGSsKtv1Pw6w3sMGNR
F0iT8FQWFkcfHYmUf6TW1tlzI1IO8O5F+WNpv/FptwCuG1S1InUVu+d/W6am+TihlWEkZvjfBl/w
WvFpQ8fU2RNfUvrWqxYlEctT4BTJDwGp2zJpkGcEDysJ2asZSaanXREWP2PD6fnuh0eOoJn9nD1d
AoCyIR8dQRGZWvC1kypTgt0MqFjMiM3fL4kzCYOMqZjJYgGhLYanQsFWhffXHtj4OfHWxXrxAV1g
20jrPfpLkeU6UNK8WSmGgV8hMgnrvhvDxRqxIllO662oS4npn4rHictVDXCyGCRPRnB8Mvcdm5BK
szpITcztofdnk2xhHYOVHnuqDk3aiRtpQ7B2e1NUUBBbB98LA7qVzFo7lIjmDHk67C2YRE45zXuc
xcMs69uc+pH/nGI2/jKqJ2W9B3792BpWxixMc2544zYYJpB04Yv9fzwDXotszyI9NBpE5bO1pWHN
bUJuYxC31lpD2DGtoYM4CX8lur6dnXig14zNfam5qkoiEqyAIOejC5pFoIYnJeOtg/fBzF30Qpbs
dsGVs3Vcr1/UhJGZciYf+3wRvePP2+vaq5c9HlpVjyQTcZSFJWhEnBMPcYU41IEAsZrWjyZf6kkK
jnCi88yRTOAVUF0kEkI4opLK/2S/dZpBsZOABhGLbtNagzQIjkb8xqgpIQmjOrReqcAQ160slIaC
JgZ3He1Hj1y3cIgU+YcTW3/dm4+blix0eqLv6rPo7AaTzOAMQP2CVa0UOZRxAfM/RC0cycClb/oc
Haww4XJkX1V5EVMxFaNORbno/NrphMBpMSfo5RUvjR8W2vPdx9PllzFT7nEWOEC6etMIAIrSrnGW
+PZC8OWEgvvsUVHAiXv+jm4163gfLCdt0EZN3wWk5TCLsR8vV8EsNcGZFXNbphDpYxOPDc4uzx7y
W0rFEUVVdHbvyELcCw98BZS0FgzKwY0XqzfIIzP6XKJOWIxxRKbIoKFHKnlJD3juENGk0wKlYq2o
Fi8z76bXRQH5D9dkiIsJ7Cj2z7R0jzSQxBCmCsFo0AAlPT8XwZMDt2vMaio0bE7gsYmFeZhkDcR5
TXEhahQxkpckou+UiYWj3ouBpC/sIsnFLeMI5BmMwOWl1c7u6/QXq9Sku7LCUf2s9BQFoG8mXwkX
rPQyO4cogynbvv5iMC4OqchpQ2ilNr2iorspztBMyNErU07LCnfZ3d8n4AroMuMG7nlm5wBaIp4B
UserqaapTDmC/PZjyIjZUSICJsGiv0dPCronMvKMSvCM5rzJqvhrn7eSDN3/zM1uFrgYJEzKHAqW
EEWy7dfv1BQsWqHbEpzXJtu5Cp/zt2JJIcj3+UFbQZ2+QeU76FmL+xX2kCuekXkfce+LOI8pa+wC
nFvrqlTm+L/wkaPj4j8uURk70oCi45N1Ht/qtHBlxwXF1r/J6tP2UXDv1x4ZQlmakKQhgA1Ix8Jv
9yz/1IcLoprl2NO0pE2Fy0bIRR7I73uiK0XA7+zs9mKZTdHGzefqdzpmYy+kJii3uvRtEm+8SALB
npEhS95rkCaWxU7nhm3KkTAryXnWEu67I5Z9nmGTp3RJ7Dn8nYp+GCIH2D3Dhrx0If8P/vPdy/cn
0md9VIjeSa1GjI6t/rgd6+EO6Wd90TLuVcm5bc50bv2B2GLPPZLBESyOqLVowLTOgsdnRR6h7MZY
E1V6p3tdUpWBksUCuiJo9pHjOzUcueIhiBmHAUHWJpKzXBBAayY5sjKvS4lFqHeg5oGZo6PgCLrM
0sfq8hwbqTTg5vZgU0OMmSBYu4YVtjN2HeCbiMuwnAUX8bt0r1kBG0vd/zQa7ax2Bb+KPKm8YmRs
rxneTa2QnVqpNa71OTxkoXwCM6KdrK3ToRbTZ5u6FvJVBaBKTzx3S9iZvnzCLRAM/+Ru9bE0LDXy
j+Nes/U3aI7gyKYtYYL7QH5JAsWAp5/lxbftXjHybpo6ibTgAj1vgdWZUvMMDx+7PerU7Pi90Q+y
lctDEVNQPqdgLeM/NvjkeRZbtDxajKiGY3za2NX/JN0VirBv6UZN6maojWlsH1xc2BTjyoq36+IH
MbxD0E5E4em78olrrf5Ar7sbuDrP4oYrAL62DjYbmt3soFMEi79boOFUGL92kuup0adFkcW3r9Tp
1/0T8qQ3DD5xeRH/Xy9f0vOSclJwMLw5azWAhEJw5+xdDmiuw+CK8oHy927N6/s2XHMrusGGzNTk
e6bhJMWZUP/KkGWLDoUE3pPSOhZbI/3YE12lu7ixiDFWme69fTQra35X7IuWXZ4myZBUvFRqIi3E
tqE9Ab4Ar74cMH20yPX33ZmzURrHFNI9Xr8CHLKkNxK/xXnsQEueBjjNm7ESRd+3JqA95RJjkWlx
4Sn7YAngvl4LJY2G0dAgAzwvgG8BPRQ8nHZhCwuxPuEpNApDaFZiQMU7dSD2NkwS7HXUJ2g+ruXD
hWWqsediov8B86GPckn9Mgdv8fD7LJ5solbMEnE0/9DeGAYF4ehsG21BFJMYdCmBNXt/vdmS9s0B
E0BflLteSx7kiXwY9eo+2p9BsjEKgvKAux66bhKT4MGHPpPGm9enk06iAgVhwIKLPhAbS0v6hzvs
bqHadFMw8VXjP3tEqg8mSitekpLTYuUOL/0Pz+c6ypwQsm0fsp6o9P8o4VS/aAoG7eb+Df2dGITn
ukBmEYhqk2/igfE4OM/PAxdkv1sdvQYxseK9X/O7ONIRGwK4pMx8WXZbrqwcybNAzM/OVsdXqnLB
zJ85FmxO/WA/qOdJWPqQFR70uG7vOvAlObkHRNtDT8j/9VQw3Vmv5NazLJEcQXbXY3c8xgflehCg
JEPGMh1osKSrRq4QWEgAxXJDsPAeTfl8i5osxLS9uy8PKIVRs+zklGQpw3X3OFXzaFo8kiIoXmlc
h3XsaE8EDW1OW+ThgRY+nlcAF7h4fuOMuG5cPnxWqPoRpchOx7XXk1B7byxljET5eocjDvDu/z4D
7uyHV8rX70v3i6dl0mL8YexaGOGhQ3m2P62e43gaBgMUdO6sBSVGK9+YL6MX+GWFO7c/VZvnM5Lf
hQIMdL8y+IZxUFNuPs1zEwsct/CeUjx0jL9mGJxUbACtw2vgdk/PUYHMNPS6pBunnsJrcsooAlY4
tiTeD6DSiBdUMAFZL8EiU3CYdoKqAWBxpsCOMi38vNIO+ZE2dZu7nhdO7aFDDrDDGcF1yJGV38JT
+o1F2i+tl85bxJy9NkNfZhyaXcFkmr6JTIXPt2O+qJAByQnSkYj5OkMLR7u9Iu2etNkgPHousrhF
gYWEyprDqbvP7MMYuiufLX/npOBFyy9ZzWdh1PLSzN5PMoqrWIsuoT4aUJ7VuVjuWJq5fxEZExLr
5CIGH1ulNd4UTNLjtN6g+gbA8q4asfDuyRuOTFggD5CRhRHip7DH15g4qxBzcr9j0RBS/buGPtbH
rlLlQgyjclBZfgJeZlB2D0HWLaF/s4nLkWG9/n0lWzr9sA1f3S2NJpNKbuccARzNg5ICBigVOupQ
ubYNLcdL8I01K3H35MIl9cO3IP4eDvvDt6yysJck6ZBH3V/LZDg36nopw23IzJGGbFQJe8Wb7KCM
0aZq45SC4el9loinI6WIZZvT9Jl8gBqGunvFc+q9cTmomKwR3n3g2k08NoX6pTbqDtmN61Piu27t
J4EBw2+Oz3IhFQVP0eVH+L+lLlibiR0x8MhQnMQUuuUvW59o6JmTXSy0ailK22WQyCIVQF3kEyOw
1snPkHdYtY9xJAX//9CNlsop7ONGw/PinDvvqNWexaX4xoN/2ccFSJDp16ClbP9CKSOg42QaQnRD
DJGsCcTLaD3Gi+lPgd3m2p4BPifFnyQImmDW1zOnKjutQ05moCDGFBDUiTfxkdIkj3it/vklxEhT
niCiRXAnoOc0F+tFKzkrADPWdKcQyFwOLAAUw4NpDNJPD3ISypVyD7fe/Sua29y72jfslpt/KhoC
G3cTQQtzvP/dg93GngNL9kSY+CLrqrd7dnmbdFXxCeEdXQQftLm9av0PaStrnddjTpOqY3dzkkGB
vX+s0K5xsZb+du0hoTvSYBiZQYZO9YPhgOYf9I/b5uyOAH9+YTRG+FOh+6UiFcefbkf4juk8Jatj
ubEdiMzz4vRUHMawWEJqPWa/HIubX04lsEWTkWHHNMyHRC4JjGs65/GnKAfT+s2RuX7VnhGv9fg6
Zzv4e0RhEQp2/lT7lvIBYGBEEF1mF8UwRQMHiITuajLdkB6hLZLkCoErq1ENAWYNvcd6w0ozg+Fw
gsbwnQQ/rjH0m8RElNeefHC5q9ve6KUTIZU7jFyQKncwAoPRz6d90b4UgJxmMVhgd6fZXA2ja1q4
AdWHfMReDZ+ZzoEda7wkLC5Y7KEH9iVqD3QNeuoSD3+S4hq/984kVT+IkW+WfU5g/mX1zT3xpChx
v2v7AA/qeazOcnae9gc6qVNWkZh58IMPt2SpcVlOj7L1+9EmporvLbU+yhcyToRQNhLyvsKsZyhP
Kh8mPPr4TYHv8Tk7sRd/+tU/xWv0+E0DDitE3NCn5sutxXZPr9a+KAlr2zlT6sR9HDXtIYQqHefO
v3xz5I3qHsBn3koW3BuE3LfFPqkX34r9eNI+tMClurTWD1lvpSOump2oJw/lC0CoTHjO33AqRh8l
BXG1FrHAdloPeFTWEVTEKOhrpY+HUdzHMoHlTcBD6aH9o2O4lmxvBYTN8174ZKfVDrZMSReEzv5L
/oKPck1hcVt42KhE2jfg+SIZOYDNEeYyEg+6CXZJobNCv2dVyNlmsHeucMtc+4CBImbWFDD61crW
FGZ/C+mzr/+SpiuHdJfaNma0zH0RXgwTsfureYT/am8VkEpS33z0iOEXi3C35bf130vZMayafj6N
Hww7ipoCtwcFXix3LpvegfK0Vni0VTHS0hJOLwvmTgGgeaP5X1eU+vXh+tErTBOmg0iZAN2Ibnz+
AP/Vb/LUpP7lq5UYv5kJfA0KmrkBFYzNjw8yopGIjYyAQMJYDDyEJNkk3ilvxvoE/RgvD9S9ezd7
p5RqcBjnmvQjdoDjpuuseXgv3pYcpBtumXy7C80LTFA68yGC4K3fyeePEethNKkyo/Osc88WQeuO
Q7bsqatCazzymoknYI3ibw9R2qo+HWWYEnWlxPXGfccqutB1BAuRDFoTX7OtavZ4UAQb0/s2AFrt
2jjDYRzRW4H71DsBLrVLT4XKQa1JNdbcR71RUp3PTTGtTiydCOwyqaSdn9Qsa5frvpVKDZXVZF9I
y7BmucuOEatHUeGWq9E1FhDD9c9s+Qz3p3u76l/vgf0BtwJaVPrslgF/0QlMn0ouj27Xdb9JYz/J
MNw5hmjTnM5p3WgPcSZvnVtiUeg2CVLSmJDCKiEAM8oibb/bnfO+qrTY0zCSUMEKQorp9c28C9oL
Um6TlsC7euajoNlI7DpEvRDwo23yDgLTAAzroVcVUDzO2+/k1DhzA8XOd90vx2zxQyRT7DBqLuqa
S9pZAWymvrkro8MfoyqnGY9D775O7+CX4J/q4/jBs7sbSZ3hVVJE8paVMbjIeZPdp1ZOpTaCfkHb
taVyZrmXVO59Cm6Ua2/vH8r2G2FyKJ6Ygj4I8DwlMTZTsedw/rm3i4/rb+z9Hr4JKsaLW7JdOQ7S
ErCht4l4/1lIk3hZ8/vVbssLIsvOw7LW6lfbzbfzleZz3IQHFtJlze3ouTcNcHY1BcA5dYtLmG8I
ZtIvcqoiV5rFhWI0T5HvoNGYw6FvEPfY/5wU+VmucsrhNyL1OTU9P03RwL5Cv8cKGgZHOLytXNL2
z6q8zIgW0sG7gkJ58QPvKh3dA08DeoPy87RRqXJyWR0hNEM5a9wJAjQGjVuB9MctvRqHDotV0S8Z
gJhzZdZ8/s7vPDcUxhCJxjuIAMAfiy8n5JYevXGIy2L79YZm2D8kD8KNFfNk6sTWkC8nSWIU1j+5
NfobY19Eu7JnjJG+QhIGLHPZ992oy9xNn4rKziPctNvcG8CJdWmYBuAG4Vltu+jUzDrUg9xPT5s7
mJ4tU14AOTIM+v2NqMCO6VbmYDx/wAl9bG6QZWCpiMw3NjrcQcVdri2CVgitMHjdKdKL+Dh2L7dI
2NtSUiC2Xw21ELaQb5dXcYcPD8c3VmEPGcc/7/Tx3+EWe8EqFP04cws7+A1arrftyBVnTjdpg/15
px6cxyjB16Y5iFlFiFQl4W9Ip7oqianSp+81tu9beVP/JK9AgVPO6H27fZl/orXXdAI+jCDmkxGI
RA6j3OiQbTxtQ86WETrtKYweHiCn4KVWeSbxbbcInHy0o7rYvVtlLAf000sgM3AO5S/JVCgi/vl6
as2t9zGrXNH6BXy/ZE2pdUZ/0SPXtiS6hp3YSTQk3OibZ3baDpZggxi1+uehz6lHBZdpBA9IudlK
fsVfza/NTPoZUS2Kf9V5RvaDeG+pqknWdRaxBx5bQdTB2BAdQdDMZU9Sm1uyx1kKmyMsPTOi8Wbs
fpR1+uoJEgZAftH1aBF6/KKCjp5WZXLdA0l+kUOFl2Jp3tB1R/r2Qg6rfLErRU6er+/gGReblWfg
eo9BhclupTF12Onxfqb5PRlwB+qg3JxSbHoLpfiei4VcpvyLsLgovTP7auIZPDRCdt8AmlegpzI3
tNkukdHErmgnUJG4y4uSxFxr4e//+ScYBYWgqktreADPwTIXUJN67rHqcy2Y3BSARIdkj0a5AVwg
hxCqltEE0g1eKQ3vh6kr/XGtfEm+PZi/nQ1S+OWLpAyEGwtWz9PpF0ybUbEbwBuFOheOnwz5E1KS
iAqTfG7JYjDPab4b8jZ1VJrMIFMPvpfxChI8Iq1oSK5djnzyzQ45ASvmcqRdOpqjJQ3maeoLPMNM
K3G1/Nw+/ATnKccnKibbvSbMjx6nJacpKjmRdgT3fmfFD8ZNtPi76Z6EEyQL6ZVaEA2isNmSsNJ4
4dGA1mDUYSyAm+6hIy0Dm8LtCv1bX5t78lhlpFOWigx7vDk/ojamTg34PKtNSPisjPUT/6CD7sw4
bytWVMt6BPDwvEol9TonGTQrZvTpWHOVfKyUX4QiEprM9/qZGmApGs7ehGsdKezXFVdpfsF1fjHp
7E+T7OXgYDhvyT113tA7NML6IBQiFJZZNmvBI5WmU5fACGR4CN9xH48LfBJOkHvZC4yOZ8pglXN0
gcVite2quvmtbVrPG7Z2eivZEMtNp7H+BMqbBLk4xBvPk+XZGeX3loMHQhZL0LBClIU4FN3m18gb
terpw1+9eCAWa1PzllcQ0+dvvput0hKgWgYn0/rDT/vQywKZHJb3LYU9E9BYLNIZRUAmrOlynoj5
mQ3WUJW10IO/QbfdppT3TPju7EO6trClKAFrh3zx6LhkfMoMscwRBxDDMSpW47mojETUteoDaX/h
KJ8OfVWGNuG70DqcS0u3u4fNLF+XEHNEVty6d8i3kkukW/8rweUH8/Rk8knJOyPh3EnbSyaaL6Y9
xHqfKfBHSQkDy2L1ddssub9ogaHus+6lrszFFCU0MP/x5N5AnvoeglNftGmuHe9bYwl/8ZbvK9wE
LPFcJiIkZjlDZG8npy9KhkRhCdVU5UKQpMsC+yQ16iyo/RN8yT+9Yh58nupQ2hOk7CL6D8PQPWoP
YPCWrdLeYPhgt0vii4Kdlf4hBzSMKGm1GleYmP4MgWmwUkY2BRvraU4fHv8NHdjoVualQH8Rcnyw
9yEVmGmRmU2LzHSp2fXAJEW5ow8ua8v2F6yIsQ9jSmFz45X0FXQx34/1sXG0K9kP/l+rdbSsom7a
nJIQuAyxlJfMg87BdpiYa1JxBIX3d2dVf0r6DkUpCXamhCHxwRMf0zd4+X1r54gyoOthX76W95L2
4tL0JvTaht9kFkZLe6k39WqNU30u5ENd23abMe50V42+RdEZQueFLEGFaymOzD4K4F8EM3ag6BqN
wU3dnYEA+ueR20nga6cFDH+ORbCKviEATP/mV7hLR+emTAc5PwQEvCEspA1feaK05bsm5PrAdYUJ
h4Wjr02iRXyhTw1ecBSFecjcqRVEh6XGzVBk1FfckcO+Cl2QvFC8HVJEyTwQ2MKMskGVjxsDPEby
OJAU7OzoclUZ5/49uQOOoJ03PUZpxuAocXNkjoZI1c/w2rgrPYnO7YahRq7ggKCOmXf06EM4YGfF
jXhh2nKsJcy5etW79R0bUb/ssZNbd7wIff0Px3TlPicEnRD5n3tyYRTAYBkl9Nc/xfEs524aqykA
E2P2M8F5YcADrHu8jpSa4YwXT6Cd0rP1WJkAWUIWcXZKyKxCUMhkPv8KIc/p/sHPMrwA0ZNtvFz/
VHI/PZEOL/I3tmS51G6fsn6SLtOs3jwzJ9kEIHSEUcDm7CDzrlYgO37DFiImgqVprjGQYTSPQSAk
ghMKlz5EX4InTX88nvt8wA7UD2Yk2tNEhBwL4QPSdmoxN4Tl+0I4DFX8uLA/fciPPXN5S16T92iV
X2H45/k8HsWMlvYtyF+zYRA6HEW8NE5/Q1aG7OykYfIaPzU+aqZFp2lBhAi2AkjdCrX7pOirWP22
OAjCOhgiMMYtRcS2vKV2ocBmSNxyc02MJa3ghkGvGTeRE1JZ+H9lt9pRn+/CJpkGJsbS3tXuBGQa
Suj+PNh5GqBYMB+PaK8GK9OwQ7oRZp6YuCpWrwkU8N3NH+nSlUsCIiuuQF0WbUvevVMISIDjdsQ4
zizFLr3lTFUYlXg1leEOM7iw2pJ2FnA+aRSzx+DTtIIDDXNB9tIBnhakK8abnEiwpXOTbh86MQZ2
5OCtdxunoSxElfDuaYAWi0P7iAWtQOub7IPXvtQn0vQVSFkvOhqpBLW4OlVfYOXl21S9m+EtcZVV
Oj74aKA9YyKlDMmbLLfcIkGp+0sBtMvOZuNMi9LhJUqGGd3axpa3CdjqO4Uo2BYX6HTPG/b37aJY
vw62LGC+DUQxy+Af7IDCnWx56gS3qmL9EbLdfB5g7nXDbA013POfoTtZ4bepEjktL0MKiPUlwPSZ
Hiyq1GNC9aAzbKeAlQujXesjxhWO4ZpsRoNHY86wMpLbcOt/of3LTP6776i/YqOWmfl+a86TWcON
FbQNcORSdnT0g84ehWD1gnf2uDkGYIUdA7yV4toKFQMLtLUZmjcjoBfsqWFJ/FBCHz3hHkPp3AKc
FckD5GE+VK57IoxoyCspiPL/emgwUGnmZjhvSphvZoLNKZnYrC3IGu2BuYUnw4AWqV4AMvcupK1c
p2Nx7fZ/Ru4QeesUAiS7i2grtwi82KOpQyL/Ti/2a/OJONtd5Hspa4hOXLzctmL6eV18ZmcZgnN4
13gwSq0FH4wwEOdRnnCnp9SyhJhhq7+x6c2pjAapeZDJxz0Ut513ZJWoHyQQSVW9qM18mlUOJoVE
QS7buQJVcMHg9t19cbERzqWPKMYk4dR8If4jIqjgexgcqk8cTQECUFD2szh0x1UzP92wcP9YKM2S
v7Ms8X3vPehIajXAbTEv2M7VR/ywYPNZhthCghmgX9oKWXjSXsGfPwnN7qkep2PqkO5I2dfQEh48
ThdoIJaQCrl5rBlC0sPxfmbQk40w90C5P7jSk1hYKvLykDZiZ82/fotqdAZgLM0JytXjz84xMh0W
FBZsQhujhhnx3dwBMqTUEd0dsbBdUakkFahX/918Yt0+tAyHjFyWW4MMy00OFsAvtGR0Mjq7H9/6
NpfQVJ2D/ZWdSysGCS1eIgLuFzR/7kuX6XftgyUlM910YStVZqiViyEvVKI6TfIGa9Sk1geGjDwB
a2vm3xbb5aPqR74pMBmhKQFUtYOQJGIkcca54QRPBvp3rALutbnwmkhytWJ+L44sS532SKzwBB/F
KTsoWx8z5h3IRj4ajJ3BDkJH45fZQn48qRnDbKTBLRHfA1nJxW8dIDrbcs7Uo5Euo3vC64P+9BiB
2bfHbeiFWs0NG9YXnKbzIYGNhLudg2KZ5+srFaPlJHVIWOxtU7VJHJHnaJMaqY+MCLS66uoQsian
iyinEVH/SCJnk4g7OZJg2CI2W1dhghcOB55OGYN4hhxwTyI+UQ4iZF8UOswuf7fMnDQUWZfjuONe
SVrLspmsayl0AbTGwxFVDjNz55gaU7I7jU3u1UPFpOFiM2wIy5hUVzJuljxCWGkXubomtdC8Wle2
AGBBQGIVByYJK0TV6uWIii16NDxShyPI6qos9Hyuakt4XZQacTDpQWbi3ROfY8P/T5bPsF0M/zH5
eeSsgBNsfpncBPeLd5vFRD+yXuN1WaCJZjwQapQUmk+XAWNt7v6R2INc328MTVM6IJe+I3osMCuO
JLmCwDzmVZ7q4M6Co2fuxi/I3byN9yZC2YOFaG6t7NYCpKyxeCA5fLBya8AxMKsTt1Ch+JTC5Kt2
pBVMBr4yAGZmltrK33YSWbgWrfn2YRyqHbsa9g18vqHJCEYw+fKBRVQnPNoKz/cIe1s9GI4lFB/S
oNlw0VtcYXy+6QykLBJ94u7KNlCFpsMB1V+vhFh/ldtueNVoL7fD3h0rjgjLwdy5v8NJLUXrQJgi
z/gHcdSA81kPjgl5mXLCnOf07XgcFkoWY1F5K/plu/3RuPoqSPFLU+xugZjkq5E33uLfbu/gE9sK
2D60U8d2mmGEoF6gOun+k87wZ4XMp2BxTAGwhhFC6PJzlTk6nOmIILURQHImjg6KiuuEiJqfc8SV
aGU8EeXb2yHoH63PChiz2ISkM5qzMZgFVPyYf5Id0lm75dq34HKmoB0/IlPefhitq5oscgFImJF8
IdTDb988BRNtCNRpNF44TI8xih3ND2Xhcns7uAT3mik8hdK+qooBLpI2+SLUPAUBLa8nJwcy/oyB
BEOGWNDwFp0a0UlE0QiCibL4ai1PuccjhG5vhpK2eIevbSPRWgn8s92LvMy16wtqJVJO89iXFfUj
/i1EAf1aC3fDcOVShUby6N3bfOAgRLMSvDYf5iwveGE08JYcz7G/MGztQ8boFw2b98eeXheQRmJv
hYUZ9VnCIpeTFX51DmzsJU/NPhP4LeuOp1ht14QJ4oENJTT2ZiufVX9YKoXc48lnnt6Q03U4PP+7
7eKiJ9k4kPyOOnZB3S7dWbA0U+sj+9pwSxg7P3UDwVuPZhGioNFZeGzgcC1lA/Pywec1k5liyIpg
OAGfNimZyKbi/dGQbM6kZdtRU4BR2bGWIMZy1VGuIR1jAULz4ASoCdb5h9o2LrSPiOElSmHLtLeq
R+Zs42Ww41BczGiaUhr0y0SpwjpLdFsxXEUFPeAIjy1zrYbcZx6zKYpbulonCsO2EEe4Zy+7OptK
DU6TTQC/ooajC3P82sKmmB6L1Jkx20dIdBo8F03rpUxOD360ynOGxv1oPA8+oD1qpyHilwHKGtsR
yOR1hAYYjRB5cIN3+0w8g8G44eBzKhPvlsvs+WOVqpP9K7V+jW2+MwNqbAFvDs0itAs6tNkCuENK
iM3BJLomAuQtKoGxj3PuRSZ+kLVAReCKfQoCJmHa5jFu5iS9Ob/W2nuUgJUplatkdZ6UGc7FRmPs
V02NsxgMqu2sEGNj4/2mXzw3yYqjxDTVA/5WDNC7MJ6oHsVDC3I2/helTfu/kJE/mYoPzlN+uRXc
5MqfzRUI/dttw4jRdLZKsPql1KYOc6Sy/IP6LjlSFXiJ2wrXiTsi3a2aPOSmqGUe3S5ZcLsHhod9
aSiCV/uU3rpVtoBuCfTWSq+vRqU9yUtqwnny3NQIBGa9h8yKYNpKHC3U5GqpyAnNUfgA7EaYJoR3
eKsAb2J3c3Cv8hQMCPu4xom31GQZKf2pKZ5a4CiIsu9gZZYYRTGF5LJgYwCy78q8gUXREebr59Ah
Ra0x5rCQOR2HJbehNf8IGZS2p4yFGFNKT3o+jvdy/ihoq3EUItbQ/InEZ0FKr1dEaDizg1O+xdBG
ely1GESZ8plpx8Ar0RfqYbjPgOxTTSaD/L2JGTQPjGB8E0aGmGWjHB4cfizB6ecMty5SmA0bg9HQ
riODwH5pckrMXpQKO+AMRd6zkeFj5N0evzUpTj1fvE5z2VNHHF0jO4jjg+JGhT8pSB3zMwe6R7D+
tI8WlA2bqCjTt9r3SeVNrqpW39jlGiFVnPNa2QCrfuckr1FGBkjiE8WPoed+dNVLBUUS9HXtutch
Lex4eSl6iP0SGM7EYbMk2YbPh47LGuirwDypNOgOPmSrmahyk3sMrPcbLqGYG35IvPQ4A92PkLKt
ZHJBs59As0LHQ15SpOL9bcFyx4Yitiv1PIvtxAUQ9HpsKBeJ8EFs6zfMuMOSoxFt8w76ZfpV1eLz
qVpbSD5RJpuCXC34WYTXYIxTwQ8ZWFR4Z57o65ZiZcI47IT7eV+BFVNb7OxnT6k6r0IKpvAoa/IK
ifY1uq25kn3lJWG1kT8HojwldUEdibtBNmzYGUgQnIEu3IudB/PulIY4iw69ORuXJGr1OOwp9wZW
oxi3YoH5Ul/bVWh9yABiHGHcxA4x4j30fUsMrYcHL1udhYHEIoHruWW15o5obGbOkY9piIlo18vK
gnR6/WiUUUKO0VTgFBTg+ZkEMoNVXaqql1bsKfnoH3qSZWkhxN90Whg4yQ80ME6Gv+CI5rK81M5g
OdZbwa8qBv1LHSU4RIjZ30vNYh7IxI3PYRd0sIl04ymoHaSWeTTMiB8RLYGfBUyGIamFq6JsPWhJ
Vxccuf9dS19e5DVRfKJC/LC436Y1ROeBKOhDv/h5QjXG/sKNx2AdMbPVIyhaLtn04gr6euHifgM+
YmZ18S/33Y+KTe4oDhsK4afd0GQ3dXFaTo3RcwZo6i3HMFt3ulw9FPWGpJgaMBO5fhJ/PqrLXtFt
dCz/EXy8KXTUSvsjG/p1OGxNOMBMJEjFFpzYgl9Th/GC+fsXOSwnphCODgZIjR+hEHnzwzpuf3aS
DRTRPlt4aPfcLivHSI2s/i7Jp89jBr/MqjjPcaMQu7kPITns7bv9xfnPC+MOjwsDCbsESnDt66Sd
sp94hGWxpKYTLvXbiMi8W0oV7bAmZCJlK/miG3Q7Ag9OVxjwmZyCJynGflvsIdO7hNb5ZP7IYJ02
TEQN4GcrNAmHzkAosHwErHQTNZcxnKGzAmGkSc195bGwg1/+9UAbmLePe02l+NZWj8xgKO57irtI
VcNI8LtYev0evCEzkKZi/SPgT21LR/IeLpIyY4r3anfVigSp77E6ncLvz1qwt+eGxOxY9qdLl2uQ
b1oR4Q+KOD2uWy6uFY0v4/CdDIP+myPMXDWOglvJT4Y/W1k7woM6DsDUdcaahrtmyJH15dQA63Or
SC/h5dpAQWrmhibgzmiE6qZThcTcl+7ZoNigUeO5/Hvsaz+vYtxqZFTN72TZXrmgkEY3+vZEERnW
pqvvvdf4ds2T+jTZjhdPACD8UM36YYlKW9yJEynW0pMKMnltYeBUd4qbjyD+80z54HYJEb9Xz3w+
7XqYqS4uUPsCjqurWwZuUkDQjQ/c9IkUKvQga7Mzw56s6HwWWB7RK0u5UHs40k4aQQJ1wJYL8VnK
sC/9kNWsf0UMpbOHH24ZHJlSVWXurUetyUkipH/OJ+6gaRHCbMyTzBm5FPvvnTHadKKmZV+3xLkq
hnwWbNKG/dbQ9Y+bDeI75TviG9nSGmbtHhLeoTfHzGykk94CKEwEAiqfm6biFiTRVPMLG2wBrS8d
JeKIDR5U8SK1tAB6Rret1M91CrguoblS7ORJCzBF7OPhtst5xHDJNgQHjPcVULqlRgayGpN0/h6t
+lTxSJyPuYV7xHUV/IvH3LVmV69jmOTv35ZKm2Q0o/tFUb2taZk3o7LWAPdza7L2Z8gOKj4J7H3x
3tCsG/MAVYns3vyfNREPZwd6uXazKvPaVTE6WpkfcwRCdskgIgtM+vHft7epSJp95rrp8An8jpfz
yYbSVVsbPO5yetZDF+zMMbZwxH1CVVZ783bT9p+MJhWfQJHuSIu/KUVNQwlJ7lU8nmV13Y2nnAN2
AXCGXb7z9exvllQNalxPzw2/gsF/0WfFr0keQD7vI4TXIQ6JNMPvhjNJydR+3rMt+oYIu3FXJq0f
Zxkv4d4IKsSD1fKGRr9oW57LeS4OW2y9afczekohh5NwHpyoxbdMyXlCJoAF7Ysl064qHm887ehU
wgH3w5CbY/CPll7uMMlyY0/3Pr3LyYFl2hmUVwg397n1YsgkpGls0+6td67ei/J7DyXhvo56W17M
LQeowEyVYnSSG3RKlUYOQA2RCKESGt+lQ92fef6GSAYLFkiLmTmaBP/Eklnapfx1uBW7YMCr8BwW
mF/4tiQbo6C+V5GNK3InGAsgChalEYri+NSZmzBFSN589LovI/b37spU4aFFcKJ+ILvbnfk/QZ8u
7dupKZ51KxD36UMyN+83Kh0akTcovxZwa+ADTkEjah4rXur1r8CgmuLy26KRIJurwrAWngNcMQKm
jwNsibTZHYXesIJTgiPKwbBNFtPf1WkeDoucZr8KK3eTiRXiSK5LVyrynbUoQFUd90nBhjCaeIZc
+Q9ZD+jLeK5gkMoKRhqTOLMfxwfaoYb6ZHufXezzSIE7K3aZ+SdpUXMlxbytLDrkVLvuF2EvKM7H
JrJecETO+VTEwr9ADXPj3x7lNvbfWhsP1h0T1fEG15/m/bgIqfdsEvVrjliGgpDJzXF69TCOrlkl
Wtod+OwLycWgV+xetYY7JHiyf+gXviJd3v438kwBpXI4uvKjTxHcm7eDM6aQ4r+0macURlnw23lu
Bu+m25dPCNClZ6B7iGatTdFeDU1HhpNZILZS0+ll1eMLHgCb+mqX3l5edAMmJqCeCi7PUNKZtLGe
phOIkov1Zr1PEm1970u/rLOrSsE99n6EtPkD2OghWKymQ96/rWjvag8PRS2MFEfuP63vaYLVIgmR
okFEcJmWXitRnk+wlemmQyhDdDWi/Aq5Aazk3Nha1N/lI0qoQW9XUWtS820r+7iRpGiosWzvhlls
t3WfqQLp/S1SO4RjKycHs+QGelztN4lNCL26TiBFyOzxgLXCUoPnflIru7LyKbc5L5BFN01lzOMh
Z0Z+SIhrO9bDJSLcEeQhO15rNxKuZB7eTo7l806o80FOxBN3FHi9js/ePED14LohK0zdTUPMWvgf
mBPhS6X0aMV3rFk5+oxUndjTH+HAudjTWFM1cbg0TCnKvv3p4bqOBEsc0rZXUAFk5xyzoiSoMkqp
OIqPZe6hH+a3ixVdIqZAN5T6I8sVx4HvBrLKs7bZPKJmIfMR8KZ+PtZI0qnmTdiwnK+9Ubp/vuxR
D8VdkzvX0V3NWLuMBCrdEe2aAfTRaA5psYtY+ljlPW/XgBd2DErOL+u7ZDlfJYU7N92BqTKk+fdw
qZYnOL7Uht0GT/DopHKlogvXd4Bh0avKNPbOw7ODsShUuhgrRp1NPp9VV6Ecd3m1cEnn7vDRCj4I
hSKqSMAXuse2Tma/1O1HA7K60iDDBjkHA2WWi19k0M6BwhfGksMQHqhODqro3f+3DXrQ/6pXZf/e
yj7qxnvtb9F63SkYmnkLR7EAFJGarsDEi9MblJBsf0kSdowU/R6Sjz3sN3SEAR/+6fBtbdJnutBA
XHjyA5LYshCvBCFh+y+SD7+4s7e4SxBrpRyh0ET1xDJD/TBTVkRCszOlJW1KQnocSu0126iz/LDd
x0pJBLKed2JVp6NvoDjKlRW6EJrYKxHNkR20WfKb5SwodRITNLSNjCiRigNGqdchIOJpBj3+wf1x
lfwF2mpr/41OSyRcniOuTLyZfYi5lnKxi0eUJaYXQhRckb+8YRPCrHmdgvGOxKaugvZwFzR62Cjc
mK7M68TmPaKtPraWpuWTqT0LI+RQVP8jlgYREtJ0M0ID663u3dRA07eysAqOs406dbothnkfurYq
EPRar5wOd6HcOdfnwrWBC0hTanV6cgaEdwGEqyR5hkMW2amMgRwxjmQQUDiduF5syCG2yNlJY1Jc
K0VeSUH0rWWK85YR/pb4Fq4wLGlAE/Jed4J5EvatrjwNl9QtaEPChUcmsdIl+DMyEtc26OdugCrw
UnVDc3OSbqCgQJpzA/fEX7JgELokToQqKIHWxqXasrBa7GYbcSYqMIb9+X6XV8UeDRKfw1lXgD0A
Ujm2Dna60m9ki3HlzD7ulJXXhiaVdtt+f25wnQkRtLYteyOSmDXqq8bB+X2CXFjtidzHb5Rap5cg
ax5zutBaa1NqIHOwYpl/3Fy+coJviBH5dIWjy5dL7XJpvpnQ5JyoCIGXKPK2NqVHTJuON0oreHk/
hdOVo5opthpPKB/3corlU5y67t2O90N0LoVPdO0YyMQ7fOHgazDpaOoSRR6LfWTEq8g1mZLrkLLo
9lhHcCMi98ncJonnYEhaVDcc9QXHsIReYSqPN6NVrWOWbLWmkh1OJSqK90dN/I9CUXYc+e5st3gy
9Nto0OMf7ZW3dEQzUZN19yo/hYJn/BiYN8FEywn/CjgQCcBADe6Xgz0hL/TFK3w6DDuWkF+0/FDV
G93Dkm6Td85Mfo7KrQFXbRaq5pRX10W7GZC0RLo8g7ANLqridUv1xBJpEbDMWllsJl9UuB4yDj6E
5m/Qx65QrwAhicxzl3/6VZD9553N1uhFglcb4rBpnG8vWdw/O1ExD2Fh6fDbmVfz1A9SVVEQa7Oj
C7I4TuVuevxfJpQcGgLEw3/xM1CAAJXd9V/rDuZRdLg4/azzon4ECGdfo0xd+VEzxrEzNDyxTu0J
jbNB5g5DjMBEoAkq2XDe3O7pxcxXw57ltzzGEmHfqGUdnbG2qa5NnmabjITyr4QA1U+WwXBDEBkB
1sOhiln+gg0iAgOJX4ym/EBxsYI5Nt4V1OWIdcnvuBLlxRdAl6cHL9wkjW9l6meC9aqLPUmS6gnf
GKa1lMMq89gIJHcEJ3XUIbG9onLFARbM3iX9xSmQfIgsoegyRh4sjx/xowh2jraMuC/4TgG62Ye6
Bq62UVQo1eBsyXR0i4wHJStkg5eJeNfuLrjKIGim2jJRhgCQU0OBUOQhnAy/grdLHZhkv2LORa9T
Fy5Wyg19/Qy1kXuGhlxD+qYG0g0+PiJkDHKCNYXQAyxNDDP25XC/99mnd2nc5AnC/EH8WQ8M3W4L
QlTeVyMxM9dV340u0MZmQ9wPGl/9fXgVu24/iqytczPik1ZaDAE8YgKt2P3fhILt56PeZgDyBj0T
Yce4ULpxeJFeqU9fxPJ5mfSRHCTk5DxIG9F8q8pDMKS4fBPlOeJmMU6nyVe6evr7aolKRzFou4SB
1tTlhc6zEkcdPAky47hvbsyYYQbL//JlenWwDGiEr2mT+GOiFpWuGXE0hZEjZ05abkjx6Iyf42Mj
Vk0FjjgnFRdHigFFgRByIE4cAzBSnNJH8THlesu6LrVETgOyTteXlxA1gGwlEqdJgAEysJGArZbF
RJyF1fair85ZIGu/THc7WM83sMxYBsdXwfKbK8ZW+B7Bl88+jZhKzLEiFtSzXHMjoJZhLJe7AvWf
0gKJzvT2CxAGQo6/OGq9fsXCr9mbulT2R6QFuKu2SFGVuEG1gaQ1EBsdjb2SHAt+2gIkHmX5HQN0
d/rFCRe2HRr0arEITHjHSZh3XtQywGLro4zJUGF2Hw9XSzIy/oRmSdf9jbe6sRNjYVZaPVZrezQR
pvTkpXbxmqZvyzcjW1ecb+kziUJxTK6NVtm1cjavwePpbcnb8ZaODCfvzHoKDEe1hf2nV1KjaXJ0
cCREOAwGpqxGBCkA4eBgg3Zlwm5wVcfYpT3vY4EMIo3i/y+QG7M/ubPmKx96OahhM8abwF7eYbw7
MNJige8o25TaUl8ICWUHge3uHfYkuFsWdXBf8hK5M0O/jG1iw6t6VnzpO8Td5wtUUwvHoLIp8gPL
o1lKnijyOPHK93rF+353cygQDrZHJYoq+cLl2lQA83LtySP0gbo+TXg0TNQ2XmcB4bTzAQ3zk7sA
eaPRBpL+Enx9tAQA7HHsh/QOA1AASqW2Cz/oCsCy57WTern3Yh41b7uIQxH3SgjCkX43XIcoAJE3
czpArusw30LZ82ZSjwbo5QDrhQSy38Y/8LCB6XQO5vfB+JKPWpItKUd/Bg7Dw+ojSL6O1q8M2TVp
J0fMIXBP47MNVpD+B/4AviR1+ISw7i2OZSFSvlAPGfQgC72W6cNfaPqvmC8D208ptXjKuCuTtn02
glpdThbmR7CMcYFTydIIhs+2bEpDPglou5LKhUfSbgJripJN9Qp4zeO/Q0dzj8lBTUxHXuTmhWGj
8H3Sesin9aepkhWxwNEoz4NSWP/rjK9+QDuho1NEyMW1SAihIEh3G6XvSqfnBQTJboWreyhZ9vOs
CuF5uYCruhXbz33YQIjtTZnPi7mXiPHswdx9chlhUXChWLjSss/CHtcLHzqkXUfb8NtI/seDZ8rz
mzThwDzuLge3vI8OMzpSw5CunNPglLYrp+aDybFtoROYEadHcEp8l53oHjjJZo3tw1BRNR7cG7Kh
c6lznEdTBR4IcQUVsio58d/XILqACoflvz2LdUI8/KY9PsWJo+A6xb0D47VhK6skiMpoTwVFZxea
qfDg24G5fFOq8Ro6bje4op9TgSICSfMOh6XFJ/Syn8sHvlU9gSBjPdfKevl6rxRR627vBS9YdErD
6Z1oAXi1b17yg1CvvaFDy5qjHO9lVKpIwlZZEaTLK1pLv0ePmTqJqqnc4Ydus7PLA/JdvY/uwQF3
R5PgelS406Rn1+DuuIlRx/AxL/BCQsLNH52r2CaN7eV6DgMBQvIp7M0YwCPtLohV4rP8xe9U0tAh
5Bmct4OiL62FijZOM6LzWo53zd2JwNTMXZH/3kswkAB0hO6I7Q6h7Kpgr9THVBiIZ2lkYFdRHkEK
iMk8fw2n/7njngFH5zQLOp29HG9t4cBDpFIsqyZXh/WpG5gofJGpZk2gbUbKVKuvV7xEPj2R0iog
jUe86Lb45V0kQv5J/q9FMURwh5A5VGWuwjbSHBGe+vTeZvrVoz6AF/OfXQnZUFCRgAUG57tq5Qli
O9bWH7VLr0TIcfQPJnN915A71HbNj3NZEYWmoolo2tlHjrBTWQJWz64UkjFnDHz9CKSu0ZQG1nM+
Pr31P5mn14+KrlP2CBnvrpEBaVSBOEy+/lElokJChKacWCOe6DIQPZ9FSShH4LdPFn92WYusLyZR
CD/S70FVUpynFSd2a1XCb/aQ/2spHnFo7vUk/DCOrUDVaPb+yibmEGzzh4cmoSFp+6HUH17QMbku
hMnhxIe8LB0EaOh8mfKUFlqxtlz1P+v0KQmbCPx8FQ9owRQI4PsfsBTayxypCZSp9My0nxMdZ5aA
HI8lO/opjggZUt9QEPIioP6gQSnzKbCsw6VHbvA5syOrQbTUw8Zc3e3rnfNLy+skjpGVMtPLDToR
n+nYibXSzFVVmD//G55zuPpZk+xciXcqSSXr+3hHrdkOfsRtFZbFQpJAyjs2JvKJEpMDMFx8LeD6
zYCChNMU+P7ccPR0zEf/3Du2S9SLYfZak4rURE4TtmDaaP0fqeMMBVbqq3MbzcVtphyHUjFy5Sh6
iauzEfGLN2eqZlP7UA0LkXg8LO89Zeae3KGlWKWcq/1g9mdRAFsLzBPMlqPJ9w4jTnmbGE4uBzgz
k2uOEe6KZLkiSmUN6HAUCw1i0u75TcuTzhtCFnG+una7dRh3guWwDY9r2/VDOpC7wsLTf4c82QtZ
ezHLhZBCMb9AAYTYHTk0FQPOxzD5XxoM2YvrfsvnEcsksr7J55E6D022lXq948otxyJ61TQrk2Q4
EwkIIl0f781m4kn5nVALNZOazv7RuxxUN/NiABxuMSgH3SpdqD8WczSEtKd0IzkpVOxO2v6skO0v
TEfg5CtS2Pkb40OYWpb4ADTYQsGAQ70tvFg5Nwq9ZjqOlBd/UmIawbTua9q6jdUUroBHL+uo/Rh5
8bdeH1XrgwTxbTkDY44vY0WWKZk/7AJwZvG4DByr5AIBfPYZZ4I1wAupfbgp/m84mqwLPMApBbkl
wlaA9U5tbKUdrz6XoAWZCPSkdwaExWirqElO8OPRjXR1AS26InIr+Zog98Pkft1kZLm+VP0OvDh9
kFFA4savSAQ79QHHNMRhgTCg+0Kc0h0x6txkotCTXJob/lHq7pXwDWtzApLF5fn1Q+J8px7LQ9x4
hXXhS52NHztExC/Gvn+7uHJreMP6/jXu8fLKLaAc1td74Tpxi3JFNinWTh3hZwF2Lavcsbsf0jsS
I+A4nfH7ZHL5yWiy+8HSxz6XlL75KzqjY4zirv3UqutkkA9ZCKi38CmwqE2kfBHOLDOQ0enc6/9t
zIXx/x6iAfUsXnJV2SSYEGf5JrHkTUr0OJ3ID9q1wN4U5UwnZTpH+0CFE1A89qCu5/spuUjtTo0z
J7QZmAfv36iZW1JKia8VMXyEj9ephP9vlgMWQI7+g0Iod7xLWodwNO9qjawlGQvIaxFeOtScM10/
6q52H/lCuglQxcNbdihw6b61Fd+eYqClx8gfLlL2HTVWEvw31HMqAYCmWwJtbQowjSsukuGHuGEO
L0Yz+tH9ooJxe9mxqSSggmeqtSKvsbHHFaLwS44sDY/sP+sghAvyeKc24o/umzFDFIj/APp9a1M/
Adf6Tk6nSYm0il/Fh5Y3mrHW9uUL+GFQ2tsyzW7r3rUsb2VApDK8bcK+9G9jgWLW/fIOBk+RWEOk
xZYXxnGuaBZEFej+TpKjfsk9GK3sGOKIxd+2naDjSRJUr/wzAv4juVyA7lBb7VEcVSBjy/d/z/Wm
SdvCgehZDN+gLNa2H/97W4AXqP1KiIbNPUZdl2NJOw+OiHgFZCiDkQvhIGR1xqah4ueQ+veeglNR
x2HjMwp6UilhVRDk2AuyTeowHexqtZ193qRltawKZV2dTjWDGPB54QhX3GxVfJThAvbGSU5x6oBP
2890UAgHFVfTC+jAdAMp2fhw2qN1mhcvA+WHzZPM0f4YV7UOa8uF0V+mHii74zMi4WmHIc+tVh1b
EbNcyrtVFa+0+GorF1E9H8MytSdivkiP6U0JsaRlfKuEW34qctmKZpmgAPR67LY/3f2Patp1Fdbm
uxrXhIoZzwmHPuEaJ4+jgQEikGwtv0gHuNIJ+gmGnUOW7vVMKs91t4gwjDU/DWCssZLkhqlimruG
KVF708UF6sfyHnfVfXcJYQXbqOh+yn0u2cuBoDimd/t1j4G1KZysi2Uvz1ar4BNxoJboEOL/BFiH
vuXZnvMWG7nhfmwr/5F2uX4h1WMOIGOJkEeCkwTxxvm8KHKjRijtAPtgbDDWZxa61EsqGri32EBl
x7N//y4JlVCjRw7xB3e8EDVGBFHlH1fbT3Bgy2s90mNezAhcKgLpi0TsUyPUoFd/oQdIGekhwyxg
t3mfpqNB/3vrn7jV88N+5dT9cSKUIW8iQfTuuhH5eyV+u8zK/ukHctciX99y2NdNwl5C8SbMAB/K
2X5gwNCJtG9b4/k3DwOHRnfNrpkQ4aY0VcDE/nti+Vid64i24ipPEBR3mH6AjLBSBpyP/Ck9PjlK
TKlINVFi8V/82Mrsw1bmOUS8b3ySOOAJNxXhmziLWFaKBCykgEJ76IIf+WxR0QPAfIXBXob5sLS+
qydswKIlxprXymtxl36EQLfv2JNj7T3QzLbjFsZFC4vU5KaYMhT/6C+7M2pMsnxZ6Obc8wq4zO8e
JF6ZG66DXZNrdvU/cBP+wsz7tUbEzYpPX1vBhWJEHmbG99ry9vB00LCV1NMaULRHWk/9HSr/RQaZ
vl5BXuOZDEdPk9tf7b6Vp09iMtlEVHgKUmTK4FD6K7UA/AXBYyMVUkzDnLpXbMjbxcmnKDDzG6dD
PLB6j+N7cd1Q1uoB3p14ucMLV45lgJ1L50J0q6wg22714NOBEtYEdKiPMKb1qp3vy7KCNkIh5FLb
GVzK5WTV73q41PyhVHp4XcwEfgWu6xB5HEIkmCgKsKzol55OmYf0m02Q5ttZyet0s9u3jEV2nik0
ByfvW+29mINVIkXBTLDysFBvrNHllkXWQUWhYzdgBDbvW/3qtha8Md6NIBsyKK+mheE+YhP4cdWO
04W5C/q5FopWfr6j/3/3GbCX+QeGMs6uBROl+Z3wT7dG2CSrFr8dWeXcmfpUPG98cG5yR6lkD71E
9jFScYhQ6w7GXHwLiuQ0AlQyq/8IbemhU/I0YZzjQ62eJSxy2nob4T9hJyWRudK+cpzM5BUnhNxw
T2gZsVds80XtcazzDfqYTx4Cth80Hte3gyprNsfCQeRW3RyXybqBEtf3cXMNW3gkGQzTLv0oE7yO
PU0DxT+y1MJyJZXuXDpNKV8mj8Y+YyRA5Sa8NitW0XBmoTDbdtbHW4iUmRD5soPOjxB+mS0aZAx0
6vZmFeFTFUkBK+E+UjnZLTThxZZ1IAB2c6dfEkLdJ3nLKWYoHS3wL7gL0+nGi538hs6N/maSx6I+
OZqVGTx82ntvBeBB6EgOj7zWVjHjypyDMQpGtLBVG3hfyoovmYJHgcZyPsHoSIoidJFN/rTJbga+
Vscv5muPfl+IfNvCNhv0NO1Dz7WXVg+mVKMbG2hFv3WFj6N7twf1zEikO/hjLdM2TMN+242EGdYW
OBSkV4T/LXgtmOKk+gm0tDkP06Rxc7jqluZYgbuYSlHoDtRVfStD10+801pBkRcW2qTE3OoaGxg2
ncz6547rqHbRnmrREfcbiSP/lFgXCVw4RKZM3iHEsUPkwdKHAq+CYRcCAC3BInCBmKAIGFejGJMw
W9fYKFHQLNQ7kcbW1yZi+UDAsYCaNJU13wULnA93j50mBTGLKCG/UJtVum8NKDSO0krlpEMmVpxi
k08zVV1IxoFfFvMxbL4UjdcB14qpWfrJD7JGWjwpNFxEf3eBdEnctUO/AG/rxILemhJmWqAVryd6
UNzw/efOCRSXRy+kthlYqf5Zf+yKhDua+5ZYEdu83SfRTwu1mtBLbmE7K4L294Zfhk2sH+i+xYoy
Wr9arb7K75VksXNEmrb9TuJkOnCzo0mpCgFcRKVmo8qC1QZz1oIrDY7iuPuhY9YSUTrF4O1Hw2Zq
jyBCHnTM0zTsYbmXe0xbukkFZm71JOFPS1M85pe11OQgUe7Y/kVaid2peG/c8ejp+Il/mkPVOTKg
U/5jGZnQvroMUcEVGAjhbkMxrfrdGgcUzRJZWb/WdMKe7MQ7n5dZLhhx7d3VtJHUc0GPzrwJhu+e
Kt+Kwk48rNi3BaW1dBCkwNs3L/IzZb5bXizX/7At0LJBORDrpNgL6TtH8t/gnP45J38FoyOVkrjS
PSfbr2HYkjaxeUcOHqfUwnpw4md0QFIoLRjOWTM44LBBANNIL8lBhW4dS0igUQVNOGMZS4qwynDj
OHSAftdD01q9IEu/zwugxuFoGY9KzzqrV8OZAl5i7nVDb2h7JZ3cCVec+EvpAFxMYbgCZ5vjQNuK
0QET40lWgjsQykTS9CPDf0Bg/mwiCUlDA3eFJ3r7YkxtsM9/P9erCFplwatvZN2YONHXricz6BBB
uT/AvkuVFK9E4Nteh4SPlt0iYgHSEG2noSnfrADKSPgRCvUZLzb6OdJ+kqgf/fNIyH0AByVSsKN/
PiQdNItwsvleXLa9LvmLDL1xZ8FaB3XEdePWYMKWK06hq+vS1LRj2sMfHb8uEPP3CqjqirTMM9qF
7Gm3BbW43WWMsGBR7I3N8flsRpVcWknwbkA56mrwwMyUYlkjmo+RjLlvQj8kibPp8EkZRVX2uDkH
8me8Ce5ccKXc/TPDpzvA8G2pKrNb/yG8mtbBxalwf+eA36HfNClsRZh5NcX8Mls7LgH+nBbM9Tbs
4I3vPAw84LaJwcTT5yp9IlVMnfV3E5sJasDgnW6wzn2eBiiw9IkAa7mvH+b3i6AnPor22b2eu9Ym
Jnlqu3AMTBQtSmbDCuqTl1bF8+AlVX+JuwEIQEnZ6uLmOuc5lZgdfBgpfEeaGtvwc41G1EPM4RCS
HabO6d3Nf1IYjUIGAYC5UC/Cx6cVRSZ3h/7EUTCkfy+4cpI/R5G6TDKCNSs94/XtAkhJmcvioun7
lxaHWG2Qui0O6LoSqWwb25FFiDAx1so8BV81Tax8Ui0NaBtTvwS2/aBd4gZ2AXv0u5crObEPNeN1
5bsOKDUL18iLNkLxabfsQ1lP8KMC/2sYrTZpj9+h3RtE1Pbe+Ohfq3oiGzNYH6bYGYCQtJqnEkcR
h63Wew5XpVxRG2eW6wT/kTiMiiqGkta5cagxJhRQ+ZVlc3C38aN+VCm9cSyqYqvsWXi/AmCj1sDR
o9x0t7BWxsiKIPJdlSefAUg25XxcZdgopzYzDUZm1L9ojmlBMbzI++ar0jfcUOCT6tcphzZ7QgC2
loXqkBLuIeiy+YboMMscKwR4B4aWPdOHmiF6eR3zpVWPb1P4tmaMihwhLQA226MJRsAJXxkqsJch
cz3K3d/mE0P+wR5pIU9FJQnGzKphecXq2oYHDF8hP/4xLR6sQWrA5LPuls5u0MDq1/y6fMBVcCpb
FsoN1Z3N6EDensxTrHJFQjw9s1e5/d/bW76Hi9548ll7+8TfHiBn6RcRrMgN/YdpfrfRnL0+L9gO
j4OPDeguH9IxaSN78TwiDw8UxND7/1DybsZVzsKsmRVIPH33PO6lzy0ucKMgvi28s95pha41YCLK
V5SSr2IRYnGc52jEtePWnYzOJkrcPVwg+7fo9mcdvb0BSJ4kqN51HDnMn+Z7qwokuUMwYow5dz3O
JAy5o0IwCx86HRWydCowIuzpJ/jVqj+lVgHvf1aDGnjy/ef48N7k/oeocGoCwUVztjlotqernfIA
VO9mSQ3j/WbTIEfM+5Oi4chU8oxBRz65Tma3hjbQZb9tIG9xOLS1YNMugANnNeB5PnORYNHDh4h6
d1YQvsXEmVLyg/7ANiN1yXLve7TsKy5RBvA9Arg7/43IFHNOc1tGPmt1VcOKcDZfFHrgxt7TFn34
001vNe+TymbjTEP9188Jjk/8pVF0dvAEaHIX1B1O2t2ub85gy1gViPaDvk1m21pSsA4YqxeIfF0W
Euxo5LfULeB1NucGSX8lqlVDeKuZr1I5IHd6v3PSBdZQ3wh3Ag38OcHHuqTSmAm0GGvJs8bQt6a4
h5YsNrQ/Z6O70C4+A7DTLzqY+BoeZtsIZoZBvocVXYuehLXWGKNycFTpTh5m3M5rpcFcf5qFBVyq
MWwdteYTyA/U2H7R5AoyETHTEdzgVLErbQymKjy1/+aNu/HYT4hZOjpznVSkmgOgvTz+8kwN3Xji
ofeHLb7hJTQF0fPXmRBMdEZBV90ujd72VjlVknJn5FgAhH642lmVZ/TzO5nrpo1fkJcSCYz2L2js
N5K+ATOgA3XGbP1CtBFgMvR2KFhFg/sOd8E3/KwO+FmGsj6pQsr/g6C7SezlkDAl+hn+gDR1ryvR
FhqP2KUoLCvjCwU1cm0nZRXJSnUU0FJ8xwmK0SvlNl8x93a6Z8VhQdCisJtSLaZ2gwjmwE/lAA0Z
nxFd2z5JirWKlCLR42anaJUmhbBkAFhohyJs1ZB3Ug0d2mYW4klp8716lnB9qEhh2BCgGLvhDG6N
4kxIIh++KYMwAdB/SDydCw/jqv8V/oOWPmus9E217J4yNhfx+778frFVUmUnx94vu0d2q0QiBi7x
grG9BxeloPBn2PEbNUpG8rgmxz5AgrnTQDxad8m9isjybXc/bhjjvJYfYWBkFvghZ4jdkWaihERO
K+sTP6DADmtRx7pTH8snD7XojmILA0Ev6Tj7QZgUixylhvCLRniKf8/U7zUkqmSJgj1CVQxCTQQU
rBgkjxbW4IZtxOZvuLD2iNF+T3fS38t6m9mU2oMNqlZJOAKUddTdX2ZuN3HTijJLCZfc5Uti80U1
TwGEdgQ8N46YM3HQy0q2VGWfIhoW0wSNsaKolOtT4UOIvKTB0AliCCGvl1NLyN700rkcymRcshbG
U8pPQpLUv/povxBt0mYVnHr8Q5PCojj5f/uW41b3OmblMuCOJhbduBG8mlVAXQuSRJ4GC3hfZNXa
BFylPLe7tAaejSt6KWR8biubeTOZloi2KKMbzjuzUEJVd2/MzidbOkyy7OMUJEJrDI3In2ipM8oM
fZv+Ht0odAGB6K36zKHVPuH0lQL7MsC6eKmXdd1SCPj+r+ftgvIvzuz819WapxIsU2wdYsESfDs3
0GN84XtgwiyZx8ptkLtPooyD6HehiqME14IWQKu0ZZ/jApIoKhMBcHHhWT/C4qGycGL9VsxsdqTD
OoQpk5+9Bkanc5q5tzcy4bnr+BFrWjEBlntuSoHhQ/Ww2WhvZuK5zP2Pf2IENHdEzOpSAT41IJAg
8uHh2kWF04ZTCO31L6VaInAeGstrMLZN8QIQFLKbSqQmeXaUaMpPS+k11DkvENM8unZR45Fc7oDG
tAYlHvUEAbXloPCj1AtvfLXkpCJKZ8spw9S+T2NnWZNUxTfo6Zrd0NqkPkeQL+NNLrxIjBjQTZAg
ue5zAAt5R/1ZTz8EX44GhrLjzTNfYsIOik9vKEaPGReFWLpYkxz/B3SaK8rsg5fcFqGjuGZtpMYk
56sm30MSLelKCdiytKECURoxz3tnrU07QbXeu6huD8fQOumziEryWbHWske8M982d85dtvGyleGc
LCXMaljq1mNmVUhQqQm28pCs9FFEMqum2w6b3xknu6foQWxBEY/fN1pIGqdq0K0gkthJWfMy4K79
tWj3W3fd3jRjr+vsyaHuuZKLOpyNWjOK9NKWHUlSDnmkWC3Zb3HRb6tvYmYcMPfjiNk2Jynhi42x
U1hRltL2zdSxFx4/E1MP8EScoLSqBd0SCbLp8n9hpoqjaGx1EAawiyX9QSxzFQNY3Ke5vic3Oqjz
p69u7xKRu3BxhI40AX0ydiDPyvznxk1C+nBaSx/AUGc1w1bk6/zBUuDIWfuWkPuwfYaWpttOynZ9
JzGNCOonD31KoYc49danRnlMkf0j/i3RJGH0mo408cIHEfvmBB+xfsfh+Op37C6F9guRh+u1JVQk
zzgyrQ2x2l6yI8GtoHd+Tm8Ln3vy2o/qka/k6JNh7EzV/6j7G8WAkwTn/t6VC2U6tu+a8kr/zQ0g
hanizCcT14lShb7JhiQ9oRu2GMFW0lcYvpCGFhbGP9jNatdfUalOeOHGV+liHvwf7I1eCZej0x0c
wANZgH0EQE1S6FKf0jqqZUOFcL0S7yKUIzqWWulVDqy0/H589flrw4kJPzIJJbSlA+ulQ29M5uS2
id/dttzz0HLmCvzcGiYydpJqFeuRB0OEu7j0Bow1nQcFRGbCu7pBqD0bD4JJgKsNiznpSFNWecpo
ULRMh33sD4zUBYbjEQ9ymKb4+D0MWbVYpIlkv4UvCeUJBhA+st/EbO765zvZ2aUOV5Phy2R9kIn6
xtHloY7Z72mfcfFZbkHSdzbpA1QqlHuTkwmWUmcLrOYmqeFqySqoumLqeV86MnOsXitjcM1jbf/u
Vxm13CaH4h7suqXXrew/IQk/uA3TFBt1ORIirIWuPeaa4P0XUspFD8IQAWZ97IGchV3znkgoTtRg
lUND8ZmIFSM9Z1XIUOwlGUHRRYgapV2OHwHOfdpXPcUqOaxXFX3h1tXvpzihtaKjZsAizjmwC5+9
TlKihLTMxY5Py4nJSWfEPaNqw9EyunHfq8hwPUklt8TQY3O83QIDAVCBOhimyG2ZmOad/awWTzRh
L4IEmKWkngCXkaX2pXT0NyBiPA5gIjfuu/EiH8AsXpjC+OMw9a2WU17MeIsXaG15OdxX9kz4bJl2
GQY4yb8zKrP0tZXZn5oL6Ree0Ero6GumONZpiBULyG5I4Xn2XoOICTYPD5bs5ogx+X7MoOYCr5AC
0pmLQrNHkFbUC4IVxi1lWOhFUBeYrIduRNOJlyrrCCib4alXoQmyhQ5QOhTxN/kXfXJh48u3GXBA
D5/UU565j3LlAMwnm2Lg7xlp/QHMEvKwFU+QfTy3wQCE+txV7r6z0epTGdSjf97Vworol7DXobwf
cGiOBlSbMWVTo67vCpqb6i0rukvy5KhYwcUeTgX6uSUEVvsoy0xcSB71z0FSsCoyWqjhSFbhFW8q
MK1d9rEEjcRViRHZIwKI8I2e0bIGfCO8lM7krDmkYRXRCVaWay+JVau2SAL5B8QzYuqXW89GeoEN
jLNis2zODR2XdpLdJgDjpP2cnwvjUNgec8ss1fm3NoxEsM23xm9R5/j9h56LmXtBOJIFhtSboItg
vPj2bdh+eCxN0BF5dCg6iLF1Mm5CuGz6mZ8lddsHudUIQgsKYnOCi1A4tfUHpbCv+dUUDr8NZ8Po
2RsIwfBv6mcpjGbq3/1bXBZVNcw4FGDJQStl/PDIV+sHuk3SdA27D7+pU13srQBlaBNiH0Gq7Eo5
vcUCcQWkdR38KzcqANiJIH1GzVyo1k6pWN3go9SfefaZvQOvoeLwaoHIEpJ54n8+1Ij1w/361jan
6pdxtLKNxR2+ZnGh9oPqn4SWn2ZAtIEb9siAmD8Dd2pe3VzLwgw9cQxVD8iTOCsR1P9rs2lcxvJN
dzC0N5UOhcz0atEtgBQl2cb1s9cnnju0XrSImqVxRMI46AMypNCxbexC158fRN/k/r50ySiT8LBw
B10an2UqvA619AhKe5Fn30Rb7bkUA6ZNnQYiHoyb7neYJ012ARTSOA1muLnmF08EQVUj0FIV9jQI
eL6s5l3qw+SmhtcPkn9dbct7ug7Sf07UHwusk8bS4rfpQcXxSf5ia5xji1YAAJf95CLhmPySDSEf
CrwKHuYO+NafCj9vSJG9vZVh6XoeAtjC5e2QYNM8HrKN1BSOLiD/udvCp6xKLiwrvqNgaSGI4FxV
6vvtMwIi+2PFQjqZ805r1aq1BMCRLmRttHg6ygmnCTHMHH2SCsGF5DQ5ZEQVYCV0dZt5PZ1HhDYm
bnvKOuEyvYnODgssxybT9b1SvT+vp0IKAfDgZ1afqh4aV8eRuAS0ZJsCK7qU1verWfSCIJjcj+Nk
HG8MFacZ0xgyu+t2nKCnkCMx336RWr7IVhcuSYC3hs0niG555aHrlQM+QlGAmAzczHZROMv/dD0H
9eBrFnGrCNrFH/tG2CioePowop4E8TU00l2fLxg2dSaSvU6RONsp/blq2XcpR3Gjn2VTZvqM3B7P
+VsMd8MGaDRhC2Tm4eQyUlARXpT78e05WZ+H0Cb45PRm6jl+bgIFsoOSfsi+mktSs1zYeJjBbyrw
741IUHTxIR8SQuwpZg6aWkxtYA/Z6LF0jHYrNo5XpP72PvOMwep/8U2nxAVLfz7hERJLP9i/ANsx
k7bzoanXeCgmk3jbz9WA7zKmmlQdoRYA3hft3x66aJZ2KsE0VPapgk+IsillvBGfoPOCs5HYMbWN
LecrTsiwcE6gytcO52vxkBkAG1nWo1RIElzpEHzowv3l6hcBylItAJtriH8jSVvqQQ6N+T2Cowz1
AQJqQKY62Suk2W4k0MGYSJjEUFPHFVOaWze3iY76jpl6JbFtU8YXB5TrvsClEn4SHDiKZNOyqutT
pg8pRPqPIZ3xx39e9mcEDLl617DidpbrlxZlqTd9My1YW5pXy+y21ndvl9Z4CwQlyXVudrkaisQc
kucD6m6SC42ckvo0v/CKIDK2cNu5i2O7K0VndgWfrz70kH46w+1tyIG9f8WYwarfjh233JqA4iM7
50oYuAcpjoW6O+wY4+4cQ8XrHSsv7B989MUCJysmFk5oug6lgZB3f2nNIIETAcDlbZTA78xMwMhX
qP3PM4wvvBU4lMKPKUzC/sfCP35XaHnhrn7Fd81v8ndZtKzFgeFTDf3Red+n0GoKhkDYxnEg6YZ/
0N1vtIbJ3idr3LlCRkbO3QxYs2/alogz0jTZxuOyPfN03GZHUTlQ/cTYE3dcg/Y+OofQ68ydE997
gqhj/AjV8MAst+zRQiUKHnthI8NpPm9OF9Yi5WjCA2tivzW/yv/zmQeMGHvnR6FJ701e7nooTdbT
Gc2sVOTlkw0/RTBOJN3+zofh2gmn5e1ZtmZZBq3bg3OzOlBYy4ITwMgaV3awC0t14rIsQH3XK8/I
5IWOD9dDb/9m4DFOSm71gxUF6/1Ayd5Aosx5MS8gZuLk1vPUfMi7hnbaKNC7TmP9vBFgiuameCOu
+6uyCijBe1FA+ij4JJbfiGOfL8hsOgEJTiHwPiAuCPbP6kFAPx8tcAaV4/GU5PTZBq8ZFskiUOvb
flVQxuAlhIwV0FF9Styu3t1TCOPlDzfY7o9qTPkXXBDsa1NLOw+zMhVms0iz5NZbp4txIMQtjWT/
URfuSJxrtJXL6yPUj1oRhvM3Sofkc04jZR7SHXfLu+jRnZvplub/dms/hLc4LNuSP6v0D3FrrkY+
roHD+xJ+w33M7y2Ai3WzztAMIDOk4eotb79TE1wmJFZdYEYd+H3XfJ7CJ+otUeVlZr/ZKQFbG3M4
nNsz8Eqiux9wru9mBmbxCKzKFJt/F0IOZNHLDVBL4E3Bz7f2BPeAuc6VE8c7eK/KJ3v+vySDyYYV
tLh2MR2NqMT2tTywXDXmhYUqM6HBzgzXmeCaSTIPjsr+Kx3iQzscd2C8FHRDNVcWoL0Sw8C/y7o3
sa7lH2lU+TyRHKDipSDkzbmjd+vQjzf7daIdb3jC2Hz7fs1Q5/00aD6GHSHroSarZyQD7d7oozsL
7toP7j7LX3iITbbOQQKqHry+SLML3KPQWMQsh7XsMYec/5xbx0EfezKkEeVDk+clKbW5nUbF2bnk
NF5BHmhLUitDxKr2ZkjPr2AY9jHLGUePp7UQUCW1SIyjIGS0y2jMQkW9ykTlvEQJfD/nosf6sAaz
/VYGfP0KC/s5VGvokJZVveg0V+PYYVqVqrywTGlGGRJ3vD2D09uM0BCEhQ0xXPTZ060Go5uuTpVN
Yt6zMZX5SUKBPkepA47m2k5BbCFB7x0SmC0/V/O+a7uFWpeB3g+VRT4tGDbYh/KmXo4Ti8K0zJ1w
xKV/8ckj+/RhkED9gyR1jDIdXXuJiDkvElKZJ4Jt8dBI1C1RLMgYWRNXoGDBhs1Y+KIU0S6brynQ
nyoM7xEK3TM40IeLLP1vRssmxNoXhwkediRTbRdMIbJ6BHFLvZh0JtnTS9/nzG3bxE63k74b41BS
LidAEymrTyiQCK0U+3Uv+d+JbblDcO1o9xsaqx9LBcpjXBR6wWL6m2fGl+6Ib9xgqxyCGpNKJmmc
8xUG0RFJphOvKcAn2h6hTME7o5554CCXborCe1c6IhEACrFgYC2cwA0xX05HKmxGCni9qEHxhcYs
uhypKk/vMRZZfMPYymIeV+t+lnIac6NaCgaKZ+tUVKMioCUNA3YBzMmYyP/abnl8OJfP06i8xw3O
hqpfLLKmspEHBWQ8Lsk/AbHd67UL6hB12mS/BGHDbwlF9SvRxo4xLYiWrQ2tLfPfC5TIExmS4pDM
bJCpGBmCdrsZDnTIexEl5rv5pL5OgEfWn4czMkJSR/Kz9h5BQM9u6l+XJ6+dOy/tCIpqizAEWV9g
NH51iU2eZA1B/wExV89wBW6bFjwFkDGM97f+LfD5IhKNiuYuSsKJDr2FIV7CePNd0rvKQasJ2F46
oic74eZsjoLIXeD3tRSMoLvfYoLWEYhS9OMBAsdMbwnZrZmcARB8yLBsNhpRMdv+pQXwQ3sjA1tu
0kLG+v3MigdRlK18/+4DNxqJkPmFi57Xq5gI2HE31n1pulXb6v7yHPxTXTKptUbGtbPoHxCdnOfZ
DQo7npiRbrcEh1Abdxa8gHVPTe8tq1PyUwM3TKEbKidZfUFpyMtkYtWpa4INmBF45EaF2VTKRTBU
NNqbs/4WEu/m7CIK9K0sl7H0hF3ZFUwzsevpB7Ps6actCVznmE0AvvF0fCh4XDmerbkEkuXj7GnL
48/PvQ9qkadR7ZqvvVJvp/6JYzMUw9rvnEWVzZSWITuWvc93PQ9oN45EKvoZFUWc9W8JgLWfYRiV
CYMjlhGlPbjHWiIJrP2ix4wx9XJSORdSTNViA1k2MSdnOxJt0tpH86Qp7mA0UvbSdCJHtwdEcG0b
kanAFpxqivlYtRtdP7bh+BJqxEV1libxsdkz/iY1BYw+qZkSe9mKrdtFTq0SpUwhp1t+bzXYuHyJ
wS/NfQr8tVhxitNfwdqtz1nIEbz2zLAW6zw6DthbTRNPOgeyZPzCXPGhOt2BClwinqOympvSWcKs
6kpGH8P/gDChIJbz7pAiFKQweQYCRYbgYTMhJBRtby6vX5v85dte6QcDZgN0/T1OWJ5YVvWTjND7
aNZMiU1i445Omwr4SNIaWjarLP5mv30BZUBnFfw+2fpTDZ1KGLRdCXITFsopbWE9XtdYG7S2UUx1
rqd5kNlRN8efFXzJ6I6U9qN4DX20uo+jzg2tFOpW99A39migqzIfgf5yAtJ3YTDC42dTqRq2A8Xx
bN61Jw9rNZJyNrJhLYZCarHvWhhVFhZdMGWeLsmHuoR99YFXMAJp5fhnmcRsaj3HLKipeinGnfct
Tps/SqcBhqc8c9yy1wa3OmKJfLo0sFXPTjoo56teAF0m7h92ujQq3CEuKR2bAzi94gSRpiqgZUmT
5E7tZPIMOJKqyO986g1eDUW1JSrLbjpH9SYgoapi6p1DBR8bffxIMi8f36mVz7QtqFL5u5OHPgWB
vEQipaWnM/WEnnBKYEVHvs7I8hiSAtTsC82WRK8LSIxUXU1fuu9SAU1vjMOxKtzKe1XHIpOSfM8C
nZSKs59U+agm6RkYTwOQxoME4taA7gxGD2xjf5NytCOxGJq3gkGnfcbTGKUPZiYsgKfNY4Kq2+19
5TXYLCsfScTRRK12VqMhqM8Cy0W481FkqrBCl+t7h6X1JYF2fdPB3nOP1RHzBoAXzxNV5bDaf+NI
WvlGKTQSvrTq2fQXvSfaLqSa6z53hJYQbp3Hfjuqavs8hrDo3k0gRMjG0ZGExpSL5pfTYLydR43U
Re/IcngS0nb29tHSBdIW4tu0LC6PEGG4fO1lp3EGqOEnhV3V1brIhdnotHhKQXgh3NBUY0s1o5Sh
gd/PI7mkw68f34fTP7wZUVLfVUvb+XTSNi63ikMyLbbUjZCxbS54G2LLHt5T8XMItmH6GzV16xEX
msRP7QQs8I4dUpbxhQNpoiFNeFD+t+wmHA8N2WP3Tq7RlaPFSEyX8NY78scUg2mnVyAJ3k/2Rcwb
CStOIakA8b4NHZACCwJEK2u+JWqV64XW64l6NKiUN/ARCIVBHaz74jnf8N+RZbIRHHNJhhDRzUXU
/oYZPpQ5wn4PcT+NXdajGdzOe/muLKtgofeAHwnrPIv52DJfKkGxhmc81v6FWlinIvyBltFFbUDo
tzoZrkBT/+Sw419cWjsjvDZCCmjhQQcNjvOA8QpfvPPMviyRgaBZaibpuYB3c0CpbsytbFId4+lt
xzZ6qiE0SKQob0uUg8e+ZCguvnEsF6dBbrV66K7pf7LNnlmu0riaxxWQ1QKj1/UhjKwmD1zATt06
90QQKCNBN9OIAj4JwVer29dxBdcZvhpVCW6l4Br4E9Ey8EouxNyF1vVwWhnIY8AWGV+5AdlS35WN
r6MqbXacR03pdwY7fC0jhyPcvYy6CDix15tBWH3SU2fgzQEGFnZyuRf3jcIcNyk9e8S+zlzmyf9u
OneiaQu0sL3jPgo7yNYokMp5uI813vOxP7sso6NC0/Yn2g0oIX39t4TNYMEuzkWdy180K1T9S+u0
88sykeRx3PUtlZjOmD5iPjA/2jCOcsiTzy6vz3lXvYkm4+nXSzVGlgQPENQCGXJxy56lRTIjJXbs
0S5DmM0cbdPSFda6qe/xl5yYwFPwyMPINf5EkJskStUUORZT9lesE9Pa7hehSpdbHPKRinIcYam7
i28WUuBBE5/smmfV8tWAbMyjA3q05lY+kSLwsulIkMYVxqoJvUwcpiU3JklWthcUI/aZRGtVXyFB
QHqVYdhKt8N8nHWiM/Zm7jpeS/O6HLKvpdb0xTcDLXwHOb5h/aL0734yg15uc9uETcL5EcV7Pe1+
wf/ACyKBe2+rbq3/XmD5SlWB0SMKsTuPdBJumGR+OBPrl1D0MDiO4E1XRvm6lSI/6pOBEU7BObbm
D0uLLFBVnAxd/XdO7Ym0RoEU6yIMfnvCoKoQRxsTf5LITo32zFY5yO6/nZQGZiShQkZWdzJ56uuY
Z+X7MOzLBwZWsLnCzS4mY1TdfyAuVE43ScwebRhTQLhrpR0S8yjkRRREfZzhrlnjpp6cu9OmMnGW
EMPAUWMVbP503xcby/IOlFeBi4ftcVNdt6s7qKIBAGBSqGyzNxW7kk+unkA5gwbcyWZM7c10qMWB
tz91uZNflaw6mg579QystPLTSye4u0ABgEH0YSQDFGga8fISr2LNrPWHGYCn4kXpOD6bQqFGdP44
MJ86kKGnuKocPc6ifxRadFn+C3Jal/4wYLFzeg1bIxDTRjFssXTTZvadSKK2UjIgVnhrmD6UEImK
VybLNmp975+khXAx9W6aZm/bUVpLMPtLp80Wd9AF1wx2+c7NK5wPfceSJbE2AOsbMvG44G7EeKyc
50GCr5cPcb5jn9m3ofidUwXh5TkhM4jobG+HBeXWSz43EfxvaSzlYECdWP+xvmnZ9l1bwovcYm4t
IAp7qJiHXqdKc6TwuZdbxqXbtfPDYYFI5cGDgpU3Rg+eGbUqC9IDQVZBjUdzx1JcxuKNcXIFy9xW
xLzx2C4BW01rMXKuUu0g6bk/dMTGQRnuHqyngpPg80e666sfqNmEEjCsLEDavD8C8txAO6JpIGZ+
zWMMJM1GMsMrKaPIq0NL1i9JYDQcuRgh324+TTDmN0JUq4TzSiP4EQTnyUQtZxiuRwiNRdoXaZzi
5qwJXsPC7cCn8uJrwwCY6OKhfTillh1AxPFdB4qDMGbsnY8+K5atX77wZETOZ+qnrSBq7fIbNr6m
1H5GC02SMPXKu888OFwbQ8sGNYHh0vba5PEXuzEDQm68txik6zamkI3fbbLeFr5t4nNRjDKwf8Be
5m4MA4NbUeHDOJdpa4YI0wHabj/RMKSYQnIrmZQnRi9BsFQUAM/31+aiQ/l1Qb5TdYx2lq3O+fHg
F9ibM/KMPW7FvN1HKF7f8B53QehUXHSKvS2gb0uuUgUG/UKbdZrAuiUjNITYA4HjxA5ZWSgb0rvQ
yP8X0EAv4xXoqwhZbCkMtZfg5Du7tjzK0gyQ8Ca+s+cNTCnzCVf2anezy7oMyAnYAu/rrfOFAOLu
aDbzxnfbxtYFBopu78WBo0gDG5Wl+bPn2TLZpebGU34Ha/5vXINGaqk5gA/f6ohIRlNnhmq/2BbC
93Sumz5wOvRWhr0UUPxq90GrgnRoKscN1tYciPRFvhumkM7nKIOVMhfwmZU/jA5CBHm3VfhdDi+n
d7XBoqEx2vwklYShCbKgukm9whTbr4jWcPcaCQ4C2UKxQuJW3W9DqqGVdIqjEgedvmfka4KGG8YL
AG8+d/rwzVhut21rBFngKAom/Hi3zMIT3nrGBKhU3cbwyrnxLmvEqStS1r0fULGoZXGmLbE/bedA
XA2ae8J5qKq04VSI0ia/l/GXliGdDuA686Tq2HQpFeBKxCIZHY1oSMYMZELcSOdyurwWXn9shzA7
Hhi2JAJYqYn4ev8zD/Aw79+uKUosVn2xyOc/iQp2jOhjBIHIbLkIcrUmrd06FV6nIBmr9oku5uN1
1e36OOyqgTEMI3iqn4W0/M0RULHfbKhz9VZ2al9HOHOtOVGXdQ2RFmZI0DGe1s3WRXvRg7O0rJd3
3E/nqJEFUVpcGC8mTzwLbW6tdPWZdQMCmHAOzJuphsLMZFs3UdA4b2oirdNE16UOEX7XbYoDoG6O
7X5407tfChrAsazPSgH7ygEdY1V0O+MWG4rf2ByL0m/JfOypBfYwFJMAd0IuwD6EBLok4PzwARL3
jp2bXkcPZtxJiFvwFjqp+u8DtTtG5vcL9A2M8UYizUfhv+8GU2JjoZ7GTNKdxo+eh58W099MbONI
iqhE0ALMCgDpVyOkkvY1uBch6I9nVt0fkHYGb4L9Q9PXA1A7SaNRHmTfWG6IScMS4CWNl2O3IkDQ
Bo2cbFVhetqTRmH12v+vmkfs5wYEMLdnGPs0Dyd9SygkuHVfKScuhUepKb0VG2Own76c3Zbb+rPd
jWVwtzkM24aPH8s9A62OzfVhrIswdhck722nVUu4pLh5553X5Uj0c0KQqObCEsB/VXqNp0Qyald3
myBG/wbB6Pjfa1Oop63FhnLyN4xpLoo2qxpwHg2H5M77KpWORKoe69tDwiWLQ8u8wHQAiK+4jr10
Izcl5LRBJ1/X754nuyuOQkvY5Msh1hYYgnuIdMoL7wjnsOuDtlgvAGU2VoOZ0+/5QCaF+n1WPLux
jnQcK2wOKLwXB9MPDK4LYNG2Zgbgqos50i6ZBxJpo7IhUf6lgYEyzqqoS+jNrOpI40HGc4a2fTxj
h+dHS92E/XjY9al5JQW7sJoGZA0jrENWYlHVB7w23ScPvxjIPVianyUNsj5TODpv1OZxefbyjOqh
PC7OgAWTAqTts77o0oqmHexXWH42VNrg55bumTz9yxFuvkSUmaoxhcgt+DMi3GpDaU/Z2SULO8yE
vwTBfpzOY4nuAY3SRbdjBHo4T7+J/OR3F0Mp/LddGcANqVVLiFc21Xa1NMx4+whox+tOfmWOMVGJ
bXK0lF1ovUWihR1tC9smclP57pjKHqKbeHSAugIrY9MDEQKVyOR5iZwb7IqFteOOv/TIKpO3tIDu
DpbzjG2L1Do83fUMW3xu6aXJsi5wD1UWEnsQQjzZNcQyd+hc5dEn1qw2N/iZPrxH/Oz/joqxDZ5v
t30H+icpLbP8Estb2Nk7b6lkCMXvHb6DD8SLt4HqQu++21/PO237Ix/VYDa7J7sk8cvVu7hsx+hm
Hpk0XNOtcrUHdbe9SEPdWyhuC757lSaka/pwO0d5yY9HuLhACU9TXRDWQwTbSv/POCth8bnZuti8
jo3BmwclponVh1iuJn3gyMgMgsmYVRT+PEJD/vQBYABosIHX3uR/R5qBIXe10NE0Qbu3b91H8sOI
fXwTC0n+kRCue5I/z2NaNg4KK89cNpSbSjcfBmsxqcO+zKWsysl1SzFNCciZeVJq0xVrGY+60YTn
xACU+RJeUlY2i7+aZYWy0jwlwsuvRk8GuYCAUhu7AZkJnOgwVs8DtJY6luueFXB7s1dkM3+FH4oF
kqx1f+eLuQS6kUOBLQBIZy2NwEYIvfmPscymOM7NSpSg1yWVIVbYMK+O/N6k55mCKdbU5KeQb7ow
8HUBr3vSiMlJyeV6TgwJAq4OpC8skeCztznZKb2CBZbyvX1EKfv81JAKjHR77Uo5EVkrwC6qC8Py
I+PAZ+SlKrO+ViR9Y9OPfVTMi7vk6vrB3e2V/WvmgwMxdoKW3P6K4Of2LMXqe1Td1PnT55JIfudV
7orKmT0R1VKhE0q0vORhmrxC8WbEavgsiar8dUZHK5OoWWShbrnFlJReqbBh81zaHKTVzE4hTHKB
xo2dItrkhZsRHVbN9o1/bsgHYqfPLCUwkbnVXSIKn2aNZ7hCaQe1Wi0HbvQEJEjsWEk0I+QwGWwf
20y//J+4RkxQXLXTWcTAxPk4+Wp3aa64maD5oaTiS5gPMx+soixBuNv3xz0osWovYyaZOZfpSOir
Vcv98RDrm9L+BRUCpk+dqWiOC67wI8JQ0HLq3P27+o7JHHIcOiOOf7TE9Y5IocI0dM4A7FRiKeq0
MUI6bl1mZhhjJgpdOChMG/fYEvNjGErGWGahwUIA5OdcWeqpBmvUY0eFprYosWI55/PGz5xj2zMG
9+fWDJTqE/+U0iZ81Wv8gwiztA7TmytTQr42w4shtLpPTYxPHReY+yLaASYt6iWsxsS/Fn2mGvmK
R9OQT+PkcAhbHyOU3z4SpkUPEzFNfGl72qKoLNQ/s4Jff8abUkcgLL60WZPpMMdLp0Tt6cETvDtd
jwNdCrLSitAJsqckG2U5UiEi51QVmppv5p2X5+ybyMy35JH10OlHo+VaT6JnbLziJxHYsebbDWxp
v4JGl1ixKMUjykD88Kfebsdo6piGcQIWJ9ZZ8w5OaaBJfSQIKikI4q0UsL1MfDWSykRCKYXjgTNt
XwdQ/iF4E/b//oB0Kisrs8tSsdD07a6NbwfSPD55kyeShlIGBYFfpFBvE4xzgRDcEy9RbGbB7hO3
Oh/lNGjUr1d+HZ/jEm9B1QjJMJo2w0xNBi3lb4Yoz5KDp98XiUK1IZep4i5JRhHBNQG7Zsafj9/1
xEiDhCaA+LEIubqxbyKnWgZOso5qJfX25pUWRHWtD3PvDRx8tT4eaTovmY5w6Woo2c6lNVKX9dLz
IjRdw42F/sG8LJV4s9H+5tBFsP8NGc036igdWAtJbA+L+jD4q8GX8/V/L/CAtUJBhxBKHsOBRw2e
a7eao7aVqzuFl/lvFErZTsaNJbuQoJB6Ct4+eOaJVgC3+1UCUIZqAjcaZ6n93eGEWzVjUvWr199/
kh+tNadb6Pd7COqMrp439QUqh/owVkayg2y+3StdIHNuPut6M8fau95TkXoaOWf3JCYm0AAcm55A
5AhuVG1vu/tBwW1T9j5EtikYL48wsUmJTg8rod4WRjaU2u7ME/hZ1y6qPSKmHw9R2xrIsBp6KD0x
HWFLdXAzKWewOoU6QsIdA57M/EBDjKMbDLiXLQb6C8NT187bYYe64DKjlEdnR86/h/EDI5690L0V
9aJysnQZCQBLT0vAjckoTjBfGlZQcxooMqfXgjmwWefmFRFVs6d5zPCawsPk1mnVeN/dKNmHlTtP
ixkqcFFBvGIki7wMgT+9NVuMI6ZNhfhy5GqwB756in5yje5+yvvqhPykjl/Yg2QQSWuh9s2WuVj3
Q9n/d62XP6X6+n9Prcr6uZ7GGkpEGfclnMALN26TQOl6nnyDUchlZ9e3Ir5WMsALUJrtVmhh34k4
1qtuO99ml0z7mK3UV/UxMYxJsLAfKOiMX/cUjp7syy/5EMYklun/OftVZBx+1Bubth/cjitUwX5/
pWS2uxqO5dqGT7MGZRiUg/xzBxBzBBu0BQcgIa9L2QPrzhLWDZwWFugVfxNI83UkSAUyTvBplY7d
w+lDaSoGn/GHt7t5fuqIoZ4nlDDmTET8GE4HDy0FaESvFnHEXZvSEgvrTT/g4fYXfj7oIGUIwC98
jOkQ9IMsR6fF0D+GWBFtuGV6JCipr+TXW3FzGSkO3yY12+9He2DXtIyO2wjKqGHBMrHFWSneMlH9
AEnzLpyybaolokveCQm5OrC5N6BYBtMR0UaCVekwX4flHJ4XflK5UvnOZWLJ7/1NoNgK3/2haHuJ
Ehu6aB0WxCVosh5vKf2sBFEZuYVzwggQzrvziJ796EYjODeiG/+ogZbIXVj3Ngix1GmaZyeQYv2z
9fvCYvyipkpxbMxP1TZQf3h7G9rgorWAYhUvrLSXsJdoRe9kNOPSfk8S+rz3ZSpUZgANqBQxIBcB
tH0KxFCngJWv6Katcq16Fu/47W/qJlHsSTBuOk7sNtX5IQZWtV3yvmJwBx8fMKdifm1LPzB7+sYo
T9QkkNaI+Z6kJA30IPFeRDhNzL0w/KaGC0IEL5/YoTsEDqGDvY1tq3iuFuAZ9c50vwE7TDA31jEx
08d28V1e+a5vi3wR2U3cE+Qr+Xcj8/Flj0xhkq4WjDluWQGmOflC2CiE6SlJlmAsWML/tsx6e7zk
JID37savTBPExhr8XncsKyLmGp+IMARwc9qqVCEWs8VkWqqlNK653GE/aKasW3zEa0NbN3EXEQKs
l+o1PhoC5//1snKxxaadGdh4F5APr2nTLs6qdHUZos0YYOKKbOQujSzWF1vXJEKtfkV5h5CaKJNo
HRFOAVv8jeVBIneAsiQATuuY6ar5aqY9o2Y//ommRyl0eLipJqPEwmNiM7TkHBEsUl3R+pc/3vbE
QhDD0l4Q08EyNyuqpWTCz7NO/VieyuC19BwJSrUCOpsKMM91/adNwY5HaRMiWNjk1pQJ1tLEjA+m
spAeBGQNE/UyuFtPUejqJo3bh9w5Pthh45bW9fpQ5+LC0/tA/Q9MmMBqu9/nCLc66tI4vd6z7GbA
DsvF83bC1n2OveX29YDh9IGs1Vd2ui6lKBOwagofI/4ldvE7U+SJr2OqK1HZBiXy+f/qZcJujOaT
XXiljt/FjIHr+/uUWAbSLHEQsaB8UyN4Uhnp4TJf7G0BrWFjZegUlvgHuVPtmthtK7PwiukCMzkz
FVZ7eTssddf/EYmk5sE3AGy3GeXv6J2LmZWjRbWJuwcqOu0ojl1BY3g6QAxpodHxaZCvcKrWMNHy
Q1Vp2ocOfgyaqzaK7SZUYdSy4sV2a1nGygGcueazLurHUkCmuUFe0pleH/dq+39Of0g/LHq/dTcF
4t5WPpU5KchCWKkb29JrAmgxz/etbc6UZJDtzWBvVLwAjipcoE2FBNIH4XE/H6nONYPktKHvZpHs
4z2veLLV9L/lreDMdX09Lyq1l24lM0Xpze0m+6uVrykLGUhVzWPT+Bo3DN2F9V63OIi1j/dnPXVv
VKwxqLt88UVS15belM6MszfuqY5NpUWHnyAxMGO9eLorRTtgd1sf2uP0yCZxIc/OpW/pyFoxWwod
ND3AXvRCGE1QPfS4UTLLOzkc5rG2dbhvEgx7kwUaB5atql2tU+nblOK0xwnud58ovH3Q8wdWLNjh
5HT77QoMRKdauAEzU+IqSyI8PzyjSQNTDTZLODnBGJi07KEOcOxwfgGg0hQiYpOO2uB6A4euPM48
Ulvpcr+NlBtRxN3OQPGzrHCBZp72KZWwQ1sYxPhArfbsSNGXbGe/GYodMjbw7hCmKZDG66jzjpN4
Qzdle+gOSTBXXc6tgk2EDWZBzbDyvErz3h11CVyT4V9Mo/AaRu2T6wxc1gN5zRTHZ627YNJeRLUJ
+Zz8tYO+pG4S96BjO0iJe5o2NJNRRgVy/87SsJjfPnCyONrDf8MLJtWZ2wEPZypi5rm3Sl7MQZLB
iWkN8KtYIW/gv0O43akew7s44UYhCo3sZCvhpv70vRH2aEgCXT+3LlaPUUaYhs4QkQsLt1Z/z9ea
02MRbGcIt8/ShOSyqaZ+c0n1fKY7O1wZ1fe4oDMahFsn0XLKy9D5mi1xNp/5zvaPOPzf42IhjFVu
OrIVRUnGdbUc6uaIXpBn5VTowjkFfHNlk7CT0u9uwrQOHHM0LhahxTBJS/wWM/vpNKM/XDgrtwAb
EaCLanC/zVq//Qwps7LJUH7lb0MJU4Jj39Ea/gmW0RYlj9tLmoQJEvReTZ025BXayzM1AdVmV94e
ytWOwMRtbstKk/JFN0ViL/3kCu1g6Oj8Yo0e5wlAJE79hDLrGgU3XHhN4bskO8fdAPOGSHpmAwlN
Euy1l/0X8liMmcmNf6xwaKu6noIq+5wvbl9ZE5GOzVRITfoQo/SE/02nTZtcLJ1ESbFlfUS9nrdw
ELPi8XBTF32KD36znJJbixXi2ZjaCRrJTZ9iVXt68yDp1w7Yy424Ml2/ySPRWdxIVBHzvBGepgMj
9/NR40M4dWeWLNPh/sg80HzWUd5WOF4DNwH5eDbDCiSlejDQ0E/8h9G0UlOPEea+T8cdHPu+KWbr
k8tN1FkRYqcY4MJhQ9Eo+XSoevKvHJERk3QmnMYS8nVIK80qEtd02029d8KyRL5sG4hhjMj4T1UZ
Zqjaeym1uA08mEgzB0fdQ1zWxxto/v932RE/2MD8HMUCxZfQWWQitwicFLHWNIZRp84mNwRIf53D
koCiNlcIPShVteR5ANVK1QDY8EcxzQ/k8mEAwS5PC2R5M7rG/aqKE2ffAuV8Hen/A8t5vj4IiYJI
G0TwKICQn6V94ujqfBHu6RTytuHEb5RQnox+PWnHosR5inI67LMIIupRHthU5AZP9/b2J2w2nJGb
Tm0G+rmEU1gjvlPjofoBkYPtDAT+D9MSbK6UZMtQ17m1RGqwbsaoe5VW4pigqUi4n/1uc9mfUQIM
s8lLOtcnkwBLF4JkJ2CuYcGcsPXyYY1opEJI4TDfU3EqoyY0KDyBHAkdrQQlu9xh0G28/bSSF+oS
inUE+ocjkE5wxjfaoGuPG305/XE1Kqj7EQj7sx3avLV0Ooaq5MEYXTw0pHdKvjlyej1MBbn6I/oo
evGERMYjw/jimCk3sD6RiB6+b2pJBv20ysYNKt4rbY2A77veC7M5Pvui4JhE1nzf5XVZsoqmI6df
PTN1L8aV7BoTrPVRom+qtxFOPok0q9sjDoAfVwlXshs4jEwH2n0QiG0xPRKBpWQ0LLSpGqDt5vNp
Y7B9s5JWLau2GWxjtQksL8bK7melgnpr/zKJ/2qqT0AQ0YqKmeiXxdtqwxbzvHskfgoo6VzhhceW
78V+TBP/NvkqnkZygD34njRpq9+HU6dKuWOZfhYTq6cMOOe50lukG1lAPBusdkoTEH7UYLtHK0LI
c5iAod0u10OoINCnLShhqY1X4kgmaXwhTlccTxmOwxsuZT0hdHZ58pz6KsEDDMVh39bYa7hj4FO2
ZT5tDV8j4ffuevHP3ylj7HD6tBXURBxKpck84yf4LJY+z3hpUM0xixzQcazDESYUhjwwVyFFuQRk
AW2M4PyYKH7Wf5mdRmRlx/eUAp0b0RsX6sIGDsAtljd8IGsTcUR+BamswDHCx3tw7H20SDfSwsg4
I2Oq0M16phCK70sbMos5mEzmeulJDXeeIgZRA8iPtIX4TsrAZRS3flHYsuPUUV2F0TMDb4J4tSXq
pXJOTN8SI5UpqlExG+TYqD1XLlR0M30HZDpJI+7vy3M1uUariiNDfAUu4I5+ch3gQSoTyzVJ/Q6k
Q7ocydTwcQgUtkNB/GeKYJypMcfiQoZOGr7fWKpTKENAej2i4oFyudcidEj0aH8Jh3V3N9triEng
mLiy5qTgZXMwC+Y9XKn2briMg1TKld4HVWrfPFgzHRqCdkMW0bUFyVEFjr/dhcVq/JaqltuNXcBj
2hFaZ++QEbZQ0HHt2/Ynpo2BV5ov+hvIh4QdgGCNzHpuY6/A9l74XK+p9M1j8tEIEM3/hXyGhKd/
oJkCMjEvXujk9yQkmrWlyv0FGFmXOU6n1o/Nto0X6uBf1qTQ0WX1EKbBpzvYVWrT3Cs2UXuMehyv
T/HyUdL1JFl0JiMAQIG7CZEkeD354L2CRQtvSc42XRVlTn5Y3BzDbLgzx7qZcw6ln4bZ/deBuRMm
amxyWHtgTZ5kx3CMpuGD0U0+kOzC3d8jPQxi3JuXfeIMbBEf9mQALmnzWcAoEh8zttm4aqXWrTCX
NL4//zsXbGheDPkOg7CypU4d95WI81VJUkV7278K2PO47VcSx3SfBkqZTwsiylWSPYOap/mOd3dB
NwQvNDoxNAE2wPyJFRXUyHIjDYI++f6O+p8GjVthGJ61HmWRVNExz9HNE5CsYz29UTNZOy6N3en1
J0nsKHJuW2sACLkpaO2DCyAAy6jtNn1QSglzTprtP58gSbb7qtcaR7iDocD96XImOwZPtt97LH0l
vqIHAqyONOCR/9dJ7KvBtyKUBAo2xOmJxgcwDfqxhZTRmpKdXehFumgJhAvML0Ispn9nI5BMmnqE
Lxipj8eNZv1XIpGG5bDktUtWgbposMi3jN3s0RQh7gAIYJPgo/vMt6XYOhAcdrQwHv/1JLhyJmKf
0QJ05Nk3NnIt5BhzVILLZ3Ao4z4MXSnztFzrn46Z8831x2K/iRSOG+bk0bYa4wUAAgE9O2sIScwv
++PVhOGeeL5WInHV6N/e/ozch/1OUa5Kfg5wEXpZLSg2ZhtC9o/b6ej0r5Va7tcFKSO2v2Lvzl2R
DF5LFYraTBtxiz1Y2nVYSEbSOQY25NH/S/1YkptD6/6DptlkB+anmqxlD1mV6dWAL45LYO0pdNs+
YGChdgYqPhRx7epbJHaT7qzvc58RKv45rRJengNzxwjPfcTGGKGK3uWh0evPnfsHEOAEqr94QcbG
wYqDLWjjyfRHXbgdv6EN2Z2XDUwxU1iEMsDn73AnpjFj1B66vWIKOsPDFOxPecR5C0gMByT0EE70
IWMeHK5y3ThQEvCafMSYKFtz/OChEOPzEQR/P8HUw0nrvEr4kr3p7Qe0lCSj0nT5gR7l/IUpx4nn
IPaj+hRN/YiLUYyLlZvmHQwtlMETlrPRiZB6eyFBHibCuI57LSPKsGu/D2GPj3fbPX7rUUqTdWtq
Jfv0QL5DZ8KEt8SRuRzvzfem3UiIZfLlkLWp8LA4J6DaqqV0C7SXjD/0cv1agK5gO0l7ljnjK0Hk
kFs2P4/EdWkmNJuz8VW+ZDAy4YK5k5olxr5Tu6dggBXfRmyAdPhJRdozMpNm/dOJT7A6yXk9jDx/
IWJOZMRhTRCYqIoGfP/5P7ATA4rXP9Ws8RxE0uL9B9mxkrcmOa5GjZ3XroNjUvLvhIGo6mZZpUSr
jRGarZPHQoQz+BPGQ6UkW/oZ2OmggMmkJV5y/8ItVqqCpOQ+P2ZmXI9Db3vczclYju4ZhrJ6/4CO
7vgXNv1kYlDkLzppWUtpc+igOgWgD9oeLfV0g3cwfJOELv6QJ0lm/HZ8VROZSteSayvuakA0QrCk
pZbCTbuHYF4CXbrhZO+SuFC9hUkMR23sox6RUNt7kK4geebmHvz60WMIODLuWLLOPdrYra0fwO55
6bpoO77FBxfh0TITQG2aLXD63lhW6kVooOJJXNJ1ZxA0gHQrhW8vFafPnl90A1wKlXKgISigKdli
t2pe2GzHP5Dih+1TobBaDIcR860511NUv5nzo/tb2tMc7WHhz4MD/gjwGv416RyxXzWV2fLitWAS
Jez8UmTZZFb5xp7knGIndhS/MB8Hf/e6yHXcgDrKvpLfKRhobkMyGM7N8uCm4r86UkUoxgDv0zFb
tmKYEwXy8Ue0HtCVofsDOthA/JVwdFGFyLZIHBObk1JjU97SCrYiZnweifhko4lFkCZWuWzkDhO6
DfpbDvhJePNGerDZMJovVYOsGwTjXhfKprJB72S+/v4CUGYVKNfWNpUPFbWM036yN0MP4wtGy76Y
3vMOwCThNFMPHw9wzREEh1vQEMFPspb2cLyViaLYo/POPiK1e94CtnFp6cgULaaUcyxTOPgLis/L
j6ZBsHUFnUBvkLGJ86s/KXuS05fI3l0tz8/Ob8Oy2eOlU88LU4x+Te2UGqnH18JKKIYOJMHFI0p8
oKitGVCJCmdCMneA+9QUzTGU8MveDA/s905kAQcqhwHFHonA3eM35sfN76GvPTaXHbdRfesW4RyV
tUMIc5QJMDEqRSc0jVm/0PfHf1h4i9yrmIcqPDOBOG9CDJVbmfLIqztRmUNb5QfZh5DXiQxCIsil
Co2tia184meRn2C6kDifIqqjVfiUjjkTXFEtkyds8EuAkUpH7mnuZ7Qq+gOMJb9uF3iEBbA4vpPB
xUmk3Bzyrl4wJhSee60yS0ooIdWPCt96MPyw51Yps5obIYa6rIJUXOAoru/dxMaSyALPZLI9RBKf
ELyIpBRuSsJfMNg1WKcSlkAdEyEzA+mh6BcFaqxAVq0qiSdCOPioGEVZYVDGn/LWP/zixhcGKfcv
gE4dKKsM3GJZhZqvq0CBxRbpWKk7usUAdTHHAG8nPOv9Sx64lKt+btGo1wrKc+T1KWXgmJ7zyTF6
ANv94zzwPwIIk5q/WNwZ4YrnmbDU29QoMRpA04oflipjAV/r4QY082VH6LQIlfHopSrAxyxEfVyY
PHB+uf9tQiBeuEOid+D5YVYWPMuQ9/MJxOCZHIGXCSHEZqesU4n3siorkiO5Ss5qUdfeLCPpYpCt
hhzmjsQLewPH2yO9lqPihDPHlTqYYpYZZyFfuK3X3sOPu9044AfMNXDXA7GAJnwq9jrRYSokReBL
FpysaskvQzT3zLbkeaZyEoFvzc/YQszVqBDtUNYnj0fQ8Wnxrdihu/KzXxduR0Rsr13W1mwwXYG3
6jn2Bw9YzoFUT/IQeEPDbWGAKukgc1geZyC8mCe1A3/zIz+nd2myuddzf6tgBB02rW7HttyIZDR+
xXuq3hPvobv1d0I6c24Cb1xVDZDlXq3UR9spKhkz9Kc9Wp2Yt3SAesyQ1TFSesiHwrnI+nU7jcWb
IaJ/ign6Z4+ya1BFdV9skOgy6jZMXhKAefah5Qp3+QEc+Kz37vkQULdT4aQ51xXhnjkSq9apa9tr
2vfsvUxs3GLB0zd9BT2yG2TLwQUnQmOS9H+mkcQT5rWyeKsAaDZKYw2Rr8fXydjN/EqDnaiUseXb
e66m0lPRiUinvtsIgNpMoEEoyQCtCrvtkNBrXzyiFlkwUmO74TZ5V15uEoevQxFTBuTt4N5DHLUM
fpn2vSxMOMT+QF2a5zPFga0Q6rK2HgREyVNqR/Nj7p9plH8SFyb7vem6srUe/Bap7Rwpc8sTQChe
jFW677zckmD71hrCTdZlB6sZTR5mUgT2stPxV6vBSBs1Zik+xXDE/NWvkl9jBDvaoQuxTSh4cqy1
Znkx5G4ciucMRTO6cVvZ3NCy/D8McQXkPPZw/49eFsLLoYtQbrsF7p36QAhXr0bqbHnNpHfkfcLQ
jpth3JkLh6exE1gp/X2AgH3Ja6iKtjaBzo4CvnaV0arvOB52KhU5FMHS1xquvuSMJyogyCsnWbJv
Rs6ErrRi59+DQASC6A18zqdP8w0HycGZ2RzoSq0ITOho9p8Y68hdoM8wjtOJmBZdQUtTp/RrI4Cl
hmq9z7Gp3FF3SLGynSOIH3qBe6V6bmo4w6fyw5lztSL2zr+XNDxEY55DTAMAcuQcGWdxbTDLACrT
GCo4GH5+uBVo+iLfkiwj+7s9RX3d2znfIs5ehTqScmK9KPSd8dtAZ7fS6+ClmuY6sF1YbAa39ySt
8+EI21PSF2bG0fxlW1FbrCaY9gVFgz5rSj1ZReMyd2fCFuRrNuTl0Egj61e+qojUmy3AaewXe8LN
vyk4OcfDgNwYiYZEFYw3AMepr/8PrTN6VnZoivkccblOqNhm7UJOv8VE4vY22AUR4EB8td5zmE/K
FaQBZhCpDk2CNGENck4T+RNnBZViRkhMAvsFaFs/0IRYFPKcJlvyNn33aTY6fv4wbGhNWTiIfIU7
grhLi2ZaZ+WcTPDIAeHOi669XHUyyAbSsyJQK+YoZ4CJa+Lch/RxVrLmMOIxm9Dl9P5IkpKDXl29
024EkQovyg83x9PpGrvBgeDmfRMZVgRGGRjYdoufPV6slrv+mVLwXihDzIx5DaRuYvJJptfvl1lc
KL3SeSOmLfhHVt1Hx26x6zyLWdQmn6zRaSHXISj/TSM9B5RTs/6bAGqyfTbu6Cd8QbscHZDeaLMC
fXIwPsVvXdQUB/xw4M533IbBkbdraC9XsAYXv69f34s83om6/2UBV36BeOycDbRRSvaxZDmEXpcN
kmLc+i7Uxg1JzlY4gF/i1+g3gmcfb2nPQz64stzmfGwW8EdDPHoq6HFSfgMA8qwZFGRauBAQStfv
H991WWBWOjjH2TSxEVE7H3F0W2ZBnarLiivlg81vJdfUMByKq/qRx50tDyc0i8O8BaPYw8GRW2kd
Q9KtqZ4YwJHffv8RHSM6mQe/NECoi+CucOJhw5RvHYQI1n60xPGBvlwg5J3lGwZw9oyvGXWkSlYc
cQiD7nGB9m+uUzs1BXl95w+VS+nA6WfNcaIcpwKnsSZ5kQtfu4E2jE+K/GlAli/+g17+LgAdAIZk
iw6yzSS8p7YZKqDNK1T7uzS1wQOZj6fWM5TTPeimWyUI0XakQTCOIZyzYd/BaTORjHY4nl/z0PAT
8NcRn6Fx1YpixfkCbI6eT14DTlxjG+vnhomNdRRrRHB7LK8tqXR3+4vcqq6QWUPmOD68XcDQNmow
ftXTG96sKd0dRx08I17/v+7W0vrtoaNSUp6WLqmaA9HnWmfx1rORiu8Oz7wNfsafERFmbTWhhh62
F4WTw46m85Z/3wlkwrF0KoHh6in5b5IAqG8QKEFbFo/Xq8/OXcw1VaABocKju6WZvqeq8WaeDdbk
IaXB2V4kXPAzgt2bo7fumiBjzvL9BIfBFsPWi0S5s902lKMd4bRhnBo+WBMqUHxemCzKnGeKuft7
UDJD073bx687AHws8K35+UEmBmtaJaUJzGFcHyob1PTMNS6rMLjgE9cnemi6uQiKmJI2qAdp36iF
fPYiMbbkX15YbgdBPy7dJCYMScJTGg+zvznMSANVUlWwlvEUSgrJNkKj5mmUVnLPDK2N3Yn+LGqo
LhRRy2iKRuG++H3q6xLYjWjZh+PUYE+1Hn+7XWIc4VBlHmN74WnfQLZYUibFPMTZ479c+pc/YCd5
knkvv/aBQOtsuwsNijo7sKgV8WNZ/Xq/MbgJeXfvBbIfZKwp82TgmxGbTPtATEtQKkBS1iaA9rZY
zztAl0L4UBc2LlOCMv6ldoKPnTdrDzUp4SYtiId3lfKqeL88mgdjCIzzh8F9Bw+62BXgwLGSyQwt
axv9SxRK8BY16MOJfZa3Z1e4XdFGyD3HX/2a+rwewVtQKAUcLDDbMTunU4KIiHz9GwVivY3lmfoP
QgiMsyHVXr/RaBCSJnqlwVCKDySH9JUfTYP0DBnZlG+nJ7Ji2FuVv+1i6bE8fux1j7KLNqqoFAeS
9e8z7sDt0HlX6u1LFJlwpvK8Qb8Dr84kAJClAetPAkRC8ZQpYu59zbd9Ks8Ezqv4Z/UodlDf1z6Y
9vXvl+pCZPI+5XLgCM4s/p1ntM5I9Wxvfcfcjk4705h6Omp7Pg/+ewe2vQ5Df1MZUS9HeYoNThgK
c1guC68KN2mg3ZA5f/S7/p31PZo7N7Rfq6v3N4AnGpVV1PUrJH+o6MV4RayWnkN7vjZGkGx0FJ3+
HKXPldIRrkLl/q4yzMMMD5g6UqhFAIEbObN4srm55T/JeMu9QcLLMbPe222zymA8tm1fm/XNnkek
kxXO8Idklhkv1tgJdfYpsXLFup0CkfhIRegJMBsxJgz3Yn7aICBRSIPAC8v7p32uWNKqM6P6HaNa
mcTi8DLGaxGNp4HGNONwAU1m15F3nN7XwAQ71lQqmR82qEbYlWO3fRWnK86yH531qOWcbbadwOie
zkcIvCFdJmCXJTN4fqrlbNE2UyqSpaVpw9QLAYWBrMcVfv1D9SM8in5aMntAOSmU4cKNFzvHt9Ny
48jg2jgL2yi98rkxAluu+1XWMX2ZaZDTy1KMHuhjm+5XADgX2QKJnNU87FXqadVOddn0HUUwwzhm
0v5zkPuYMc6Q16ajiR6oASeEfO7tacKWKIISYqYERGPNmJIMBzcEN8Z+QCsiM/9IfwhtMxjyMCcN
0/xLCpWXQSq82WoEU0jYGjhz/OzoDM+8fWUwh5jdw6+iBZrHA52Vx30iyZjZdv9hO8crbp5Ujwk0
uPp8GOAzC0YL5Gb4wtClbqVnhPuDNqLlnqoKp6hTWjZJjqOhOz2IViTmiqqrrgCiToRfW8YODLIU
PNJbVbf65DtOmsoKXE6xuGsOb0CjTX5wl8DhsDw8YTE7ewhRMU6IsAjASoMk07Hc4gJUMPr8Pksc
Q2E/PEMMgCclhrsXiNtaASnM8YK/R1VyXuN872tkjKo4oLeqvF2c5AoOyqU3l9sbCwWnS+L+Fsc6
oWcmsSx1o/n8Xju7iLrBtPLBOqMgiVF0Qv87x5NDl+3iN8NoBQfUvvg5MnFNNbiFgW9ZQputnXTA
ChV54n5DzJv8P9/kD67alSbWxhKdhZODzdlZAcG6V6ApAE62Dyi/TDAe59sEkuEjV7F5qGa+b95k
63ABQfNGKAkslPmCnATbDokge+1nghUSWDLEbrAoR038T+LL+ellSRi77nvBwI8F1EKGaiYvOcAM
SkiknOU4LinKajA6zzNmTtPmE0e6tN6fiklKUb7hNtAcBkt7ugofEsJrag9+1FtVFhL/C9T6hN/r
RpnGsl9SXAwAxDKZBjcj11+Aaxu4DGyXV6T9yvMAkWweoPO8ix6COo9h0emT724Y4ZrUIW54HhC0
W0L48wV/6Q2WSsHeOEXu0FL60azkfwUYaQkLrKSnXW9voQhKwrpoqPHIb//nXk7OA7iLDr2HX2wc
ZtkZg6nmgENqtQkMsJFv4kJ5ZNobbO9pd/PjwFSUD6cTuPvmhetwp/cVUfLxu9+MCAYcEOTVhjUa
6N1aaNxzVuDaQ/Rgen/pehlHclwyRusCGeiVrJZX2KSFlToGprLnFklU5Qvr/yOLAP3LZTAGUe/z
AOrg1z5/qEYKjYHC783G09Bnoo+4QCdANQbuygoCTvlkvx/WpZgnqBfyUXWHNO2P+yq2kepmwJod
Hm050oCZZp3MAqtvSdMVarvzUKRCBTeHO+JQZxC23G2zaWvVS+OgUA58gNlD8ZAlViNBwaGKsjus
vYOwsM4fmtvMgDX6txaotMxo55y1cftpsT64OsMkr+RlmD23NsnVPcy9d1t3woLguc16TDTn9mV7
oHdDtjRmO/E9dSPUeQsClkS7hpDsvJW7Wx8klAUQlIlGSBPZcPJY17ltzCjPExQctFD2WJ8MAB8i
cv3n0bW74kleEouGdqblvnls4nki8Fl7J5JiY0gHvDzezaRn8TnJme6cuSs0u388nBqR3VPgYpN4
xLT9lGOKKgxFgnZ8y1JFp93bLxVJnNG8Ve58V9K/I0Cks0aqOHEOkgBmud8ovLaJL5mLR/TNpLMZ
pJGLqh2tfOGVZG2H5MbAIOSMZVdECj9izx9D3MT0FVB0v6434KUOozcJRGKzn8zJLwx5LSPscXlq
nNA9Kg7oA4rEJtmWgU8Eos1SUlkyC23gkTBU0khxRITr4dWmK71nwE0UAOytWomq2kpQW/0Rs5HG
cSPmc3QE+QfNTyMFWjvMtwQlCODen84sxG3NTNfm8EehZBa0ZMNbcmFqrzMXImPFnT/wIMdwzV31
AAwc7O4qFw1sTx/RIWyeLO+CobKRijdXjL1ziF2P3bVKvBIVbIJRLTnhsVE97GdT1AMTDkK3HwD4
OwkbFlbkDDzC3jSozo17ZB+L4yZ48G8td+7cSvXp60NfV6XsZHuHc0WgMBHzUx3HmUdld7nbne2V
b3AADell5JyC2GCLVsThc3OTVh9UuXn+islkLEbBCOXgasKOjPAVeF7CA7LHMDvaNQK1J63SQU70
fn823nNQFn88B7JaqY8TdSqxFPMC0NtOQp+3q34VDTHGJAO2q8Ubsxfx0HJs7jNMeN0r8wq7cliG
4X6MvPzov7JwadMN/PYh2ygD+0Cxtwd16hRrhQAyD0KH4GYBZYNhg9pRMe2hA/KE/LRDbXbDNNFH
el6Bv0/u9MkX8LdUZctWBqyEv5u8AABEF41DCv6bFAWuGvDy4SmxGVnOEyM2AzBtWMwubH90CZ8x
WXI+X/MDhwQcdwT99fhOKBiFNPJYvsMMa9FZGwb4ajGs0ADN4xJ69Czvf/YndIkr5GWEp9OuOF4k
jIBUWOyG4piCt/DI/UhZLknl1pdr72+pf/V7wz4zi8YqTpTFZISS1KhScbWeOi9iJqGexXURVT1J
IDL5lHqj+C/tA1734BIC2nKOn9Il0fYdcmTRskvPRcTtJHDn931vd+cWrrormS9dLF8vxfM5E+UO
nyuTUbeUciwkB4/LWrGADVHXT7066VBBg5YVmdfJp8MKAysgPhY6Owtvez4wcdk3pnONh47GW9fj
bm1IFDJu29Yhqlv0fxyJcdK8Ue1w96NNxEQOuJtwq4D7sYOFRpr+Uxp+a3jvZQJ2kPp2tSRw2rC9
VFV3IFTSr55hM3pIL8/dzWUAlDtLJFvwPW+Sj8aREx2kaaVKO326P8q+V5HgiYZnsSP5UYEA+OR0
6PwOQ3F9hZ2zcXH1KMcMt0KyNm8j1B4CT7tJleWgb4hTQPbYil7wHLM+DICMU6Nme8234sEoEO2T
Ce+JUtjUpMtvrSfshOnPUFI7fRpVoZ4aco/hHlDZVRSp/PnVaawCrAERBezOlVuQZv3Y4Bnu3Nqy
LZZGCTRk4diDVYWnOQ6INhgcsesCSeqzbIbydXGP2MTXXSL+SQ3Fyi/8h4iwOEkENThA3onsfF/g
2XY0x7nX/zXRrj22ROSXrF7f3BHA5iMPFa6dKQSz685VtVSO3f6W58ckcFdTYi7N6KIRV6dHZcss
NuYg+0TCc94YbjT3pFTk815OvbkNdnyxFx1G/SbMrDO8sYRRAFkCEx9nxG8S49EsSOaunKVe12XI
OWWLyfteifBmlcljF/vhEsbp0qBmec5iXFdQyzX0ik++nRWqBy2nY04TNNYqvEXd+o5RALE9EEGC
K+wyKLY/+s1vt3unX+z0XABE00y57Ya2LFmBB8Yr/nyhAsH8aQA2DQmo/hb3GrIfMgff/5xixrD1
0mW7cZ5JPJmUwoQHCjZ7H3BBvDA1ehxiWV/UrLZh6smO+trZWVBNebdC4cDd4oj4FacGKYTOcH+Q
WvDGbCQauoXrWERcGyfP6Z5SYCeVDT0Kku2CJkD4/VQ05Qv737KkwFDyb8n4MtrYqCjH15x229I8
EOUMkg3KzJQuHKwUlnoaGbQ87WaTY5cJxqK9NMPtsXaVa8Rk2EWLabbaWm3SwxEPCdjIKQDFZPt3
JkTN/gF9MIdVUspJKUg1SEQfvmJXZlHdekh3j9B5qdLCXiTRLw5OlEuNPVfpaCenSQZK/Gwi6FyL
wbaZZ/HFKIIHCtTpO+I1W410mS7Grmp5NvCCdIB3kl3qJ1pVn5eO0OrfONcIsNzv9ZPFsCejhnVm
LrEv3CNCxge1+2FLknIZTdECSgfNxbC/WjQHX4O1R4JcxQ8nlIdi8ceR/xn9ALuAwRPa65i3t4Zl
aRiImytpQH0XyPKSOu15vHxBqD5S+vYafj+eaOoSf+x9v5HvurfFPLXUdcTUi4E7YW+yWAVyCU6e
+2D3iuRMtMMv80SxPJXAUZWOHRSEl35iMYkPaw/jHgFkcSiSO1eei1cCWJpJjQ+fss01cmQouEEU
S9ZnSiaorlWkW+A6gYYpLG1Cb/Detmnkne9AZJ6ye7daqlUsaHiGyLh3hccgtN8oV6G6vXFoPUTW
1dV4xjJKjIDYK60dQRSOie0D5g+sLxc82K8q6YgczDS33ll5RW+TI2MeCqPUfWOXxsPQwE+xxuBL
iT6EjW9f0ai97zzGFg/W/RTlUY20VupcH8JdkYrzeCcxBwjND4e7AbjsODrNCufqJZkIRDpTdjfV
aGCFeEe4cjEyycVe98FHEIexczV4NFbzpvscQSNd/wm07QvEyvQj5HqnUQdWGxr8fBvmkgQDSJL0
uY3G/IH8bLAuiDdvKRVSeIbHYPpIj9rVjkmHIdsYckuKxnU/6I2HeFP5C47giRrNqLnc4flLgTZi
HKucuAdGLzoNOFuBqOtB/dPIjmy5KhT5uLqe1+qxBXqfaLUeeDw8SO0qgxg3j/FmsdbXn5zBbOl6
DdRnlcFjmHIIEAqYfckKXsp0fGBd/pXRDVqT3H8YPs7q438f3MVvyB0m9lEknnDB+XvXOJqAlnPY
yWqqfPSnk/1YMvFt07TVz9Ye3tzAPaacqEymtsFSZ4gAh0aFNhCsIQCPJqVSj+44Jx959PO2u8J1
7LCPCXBRBblW3cJJcP1EpXTBV11ii+embpjsO7hlHQwvzHp/HekocwfWitI3uvhEIlQd8b3V3zdB
RGZd+uSJ9hblw0X4VSfrcLuxo/ejXIfbBsOmi9zlD6LJzojeI8j8ezAdr85z8c+kUG+/31NvoTld
KHOQqAFEistS/uEYMQLS4ZSRuhmfleH6N/v0Sh5JB2V8ktRf3zP0q1mxonlph7EShclH1EpCUUfe
7QCws0Inxk1sG7PiPRirI5nTs9chRJzicQmboN81T7aDod8ox5ZDKvURUSCcekCDtnlDKzgR07OJ
y1K+0+KgKbAWjccr6NyouOR26b7Q+eYXtPM7jD96eOeBMcQD4LWGEQFOJrcCqynwdNQYKVgUq8Sw
8EBe1HM+E1+UdodOra3mWToTXt8tMs+/1//jGTcKj4xWfMAqBP64MKYn6313VsidKEobGeOhjWH7
NzOORr7AVu19liSatQBT4pxm/C4ruVF/wHLmLSytsslngKaB2aJA0cwHOuXQrwRXXmm686Ni+Z4i
Ev/6Ybefn9HfYFeiWckM4E9EEfejsaGl6IXc/kLajH3BAlTHMI63oKy2RQ0+/Ls7iwWKqol1QtEZ
qpByo4ZQ0FN5sw3g0yFS7tW6UotbVb7CMsMvABCaOMq6bijW6Q+/dW16BYvqeuZIg3jhQYzVZiJc
HkDASvz/2RRLlVTRryk58X322/vpdNT5Hf6l159RQN48oVYtCNuqP+7qiBN3QuSMykjWNLEt8Yx1
cGbGh6NrVjCwuIhouBs6s9YD47I4Zs0BFKmIXidqN7ozo3Kjlw3CRyd2p/uBvxBAU4yCNzMdEm4z
xaLmFAgIHZaItTV7x3cv7T/5y5mXSGdnXCQ+fzfDKs4OobcV2XNyXoFtR/GGMNrQy5/JxyfY7I1L
il8MJ9nmeubYgflLQJhynKQPBQJZNVlBh2CHBF+YMw2A1XGsOckfKn/Bo6FT9Owq5ykM02MzIwbg
9LxNmMQONJ69bzpEXIdVHtBpmIXuJV4CSx0Gd2sMpwGkcRztQtfPG4PTSX6PoLN+Mg+9aM2g5ffJ
qDG1aW9PLQASWjVDjTDipV3WwFbRVFB4CWFB4Dxeb4wSgMGY3YCrvl7R7X6N3KAsJDnzZBa7G1tF
BDoYCHsZWj3u/QKDAdCioaW/HJy9NJmERrP1P8jv8F7rODpJH+OugXvrShXEVYc5CHZSRDSp3pZJ
tNOLv8udO5imdbLi9FvF/SuaCu1wMVTzTO66FT6qUDrt2+LxbdA9ZhrXMomDa3vF9iP2Cj1mztp0
OJnOTy9jH+/8jEGaM5du0FC6qH7/kPFxEaaaaTneq27ggBBOIQLpD5MujQhbAOu7cPh3Yj+MglUq
m+iThNGw0f/L7xfzPLBOOMalrwoDmWPB6EjR/yHdiriSl3cvARzt8BQV7yHEymOk+GPHs1Thb5vK
TjXpNthx6H41mvuvzOHxKvuzni9Plt08PnMZ9+LPeg6EVqHKTTqu+VhhHlzdpeXw4UcAXTBesy4c
o7JGzcPFCXriI3gXFZdDE8hFCT7peoyO0xp0wgzMzQavQk5Y50V9id+zKFe5P8QOf4WuU83Ks2Lm
XxvmGpPLqL/3MazA3GgIAW8IOAwi1i4GlkSrgvgQTjIdLYkMvYbXv6y5O+jtd/FGOqUOu1XHM9w3
TiUfO3vgmyvcxgdx/XY5vNicpDwdanVhi2I1j6ZRmvyUXsKQ8yEAuCqMEoE20peCMBTDf3hsCkDE
TxRLfSlVTb//byTs7kx/NpFT+xqiiJS0R9sI1K2Rs4eGIoEocOcn7HH2U1eKVuXENujsbmSLdnx7
v4Ln0TPGaE/thwdPA6zpuP2BYgcMI1v2b/a54SXD27KKXNa1ebdQ4W3nH05IkTeOyZ8sWIJgZ91E
PaE81R7+Ldch0Grgvjm/XanCEwjxIeT0ZnD/Hrhfo0LjV4B/kDSS5+VVQESx8JB+yBTYPa4pjMbv
lZFtIHnnsPTyDFmeeOhepUjSNh9icWjjzkQF6epZGCA208rAeu0NIDAaygLD+tdld6Wcehgbo9Pb
Utj4PXvUpaoAXovAtHR+zT4oTwnU94a5dbdZCq4+Prwu42AXWtR3DfzG9Fk5S970W6bhOiZUQZra
vslbmOXIY/2GvqWzxSijJ59SO2hIOQyNSshFFA2UlXpLqHaYHNjBcfjq8mjeS/RiByxP+zZUDw5s
90cvATqYHJ3oMAXXfNQNL3cdCAUeuwI+R9rrSeofKKbBNdPgN8tzpuY7BH3VLN29xNxn/jv3THiP
darGKcp+QJjPma/pHlTqPtJQhGbM2YYWxq++audrbfUSr4+te6O55SgUv0uGP3zg3u5LagJzO7uh
zuT2870fgyIpttk+XnFdCyAoMbBTYrwpoc2KdTC+SuBlFO9wkru0YBnKMbz6HBSTBl7jKQZA0+KA
WDmnd/8y38LYlo68fKWiaHYOaK0wbekePwfogf/7YIvBA1VtyTysNFPlNP5hYiEJZps/1RLVTsAt
R6sCUR9QQoohQHZUf+csMvqdg6u9BRk7yGBW4hleNBNSBIOmSHvCV7zPG9TQdeijNU/TaQM2pJ6C
DiZ9Z0rZ61b6JrwcFCaz0cMQ8wyhVwZ0YliHoSNOHewJidw64kEeXgP/sh0L23cQhfLxWBoI/Vdw
C6zpwFpx98/mGMFuMff5VUIZ3VpKn4ClJvXLeT64UBikXx9cCCwmcl5Lp9T+JQchaK59j+ko7bTl
DDBK3HhwEwTcAdGDl3FIVis9YhCIirKHB7Q+pSDvqWpXjJeLERkICKOnb7r/SOJZ4A0TBSZFnBsC
RCV+nWE2KweOGQk0fLITAO0wQVZOh4njmeeGgHSojDKrXU6/idTTNSAMEx6DKYehgFlZtGLeFJQV
JpwaOjBdkh4eVpN97m9in2ewWgSbYq/UDotJFSqsL5nhm84jIQ2Hh0aUMfJOnRGjiKbXDJi95r47
2wCrmlmMNBWkqdtKl0c7MCWHFGrDEi7+T3zCLLiLWXsUecJWmygkFv7FWSQJZhJlu8+/CZcDxH9o
HUVDNKfV6fza0DQHvgIl5rZ+j+xE3E9bqA5tPRjhNVB3o0VRSgCSmv/lMNK8wwvBXjZtiXLVkkz+
8MLiv488M756It9fpx6AmHkL/NCTSOgOOCZCw47jbCFKZAYfrPHIdGr5QJanLqMPv9ss4GpUVi5U
9lmyK58eM0ufTsZ0VAoMByJbnsfzy1vPxI9KXiMhUkvP+fjwdfRRGuTD6XK68L6X/U8Kg6+XmG8e
zqRhWocldAnz8emHcsesofZGqen1n98MjQbmwtJ6e3FI+PB4Xe/xweH5mlQko6PlFo6TJVZWmI6z
MULaJumsCFq3kxDOjEkCW0YeltulfyfGMCusRvrCoZYbOYUreGLCp6PLYTv9czd299tRQc9k8NHe
bTa5QGLm7faxmbNsDhJ7L2hfct244EvODQxKhqrCB3Kv26by3+4uo7yNQtCxY5BxsyctZ5qazL1x
q25jDYv8oNiswflUoGvLCQhknZrwVw3ygFf2FWGfQHte3DWVnZSA7Bn59q2jb6kKDLM9stR1c1Hb
gRiyP89DnTwGUrhIaOL0Hj+QtgkMVCwlh5jDDFoUP9PYgKFY1GDBMMzTDDh8lNzkWZM3aT9q05WE
uJfSdrp12srFyjQ+BdIodQte63XskGCQv8zJ0nz2gvIoIldxxoJmI6tcpomXjwHT+JkJ6mQtgeVF
NrwVTyRmvkOUuiksqEa8pC6rOEOrrFf+b4CB4pcPa/xQRfC/URl4NR8FqLsVVGEaWr4WJUgQQAWt
VB1tjNtQHYjA+JHjl7dXAa/KhC+UivPlFa8OrsTtC3ZV9KMc07COzAdKnGlSSW0DOZb+ibxC1PGr
xm5ziSP+J35jchmrsGpbUgoh0VsdqmjoBbhuETJREwnjS2/aqPU1u+ueobyMh5Lwxclt2ShviDde
6deKvU6vsbUoidCUH8U7++okxM3hV+0mBwXw2fGxQyfF3GCDtS1HKczAHMmxxMfa6gq2mM+ABag6
huZ1G+gFPui6cCXlxXTq8WThySISMO5EJc1yIsrjyN+SyUClSlW09Y6IgEUp4cx6Lls9RfLMbvaT
VLHfU0wvvk1ZNodBo2w222hTp0TGAR4mzhEd01MzyUfjl6WebsvGs1NXtOuiaxGXzRGfsTqZIUG4
4qNnei1g7y8w40I4xuzk4xy07cD8AKWnBtYZrkYWamUgpV/jftgzyIdT10vydv7oRkJA0yEjx0aq
L3PROK5Vj+4WT7JE6OJc5FNOtYJOMBCvADmt9Iuy/+l66KWki03msqeC8WciJFe1QqT+yK/vKqNi
nIHjWRkaL0GnJTEAItDlALVr3FAQYzuEunN5zKacDvOX7KKwfrTDbFKtdnIkR3uu7WIPMLMo76SD
+M0Wb0+GFtvQzOUXoDeX9k5cdeE3ePOEUqyWzBsmrdwbphUyQmc+phAas+S9l0rRlKKG4yEs/Z71
ia/wb9/PkBR62w+quKEE1niAPAWr4eTcBNjA1baR83EVRuMXUK4Fw/vU93xjKaEy5nKfZbxi6tnc
DIsC5IQ4efOQIwm9oH5KlIDHCOyMYXx4ESJaBq0SjfqAaNcTZ1uIgD8V6MeTz9yc027KpQXkS7fy
ad+30xpYOZk1zFGzmTLMWob7D/NDghnMNQYUmvYCS6Oi7TcjRGHS37jitAKIFqd3vnXMM7JuLYne
oHJug58eQAMDKPyB/dNPsVdVl6+j3nS1biIKRYZ7KeoSydOyoaikiUVG98NlvZvpzhRw3cgOJvlk
gRqWfIlWBCaoJi17QBswmejSfKaiq3yHyhgQfyxnIJ0MGpc5lTrbHpOoOW1j5xBG8TIBaL5MQcTH
g3JDQ4zTfwQeLIlgI05E2UqvHPwudYaZJmwZhy+j0waBFe0jiltcsOciAZxGxjaDwNFppS0nAW0J
T1cs3k6cykhRYIEoFcBe+ybNWV4j55mwc3WeoTxb13JwfcDJNz7yynN+GbIUeKEwtULbFzpakSWk
yOAIBTDo0MMP/1111RayxKx1AHZW/6SF7Kn/rZjGXFr+Me6xQrMXB49zV39zDxZA50t55iwpIh0m
yX60uJ9vmeqSrXsA48rZ6PLwWcN7bcf8I/xHA1+cD4NAxGTZHkMC2hutAALmRUVmfVOiJF4ZBCEB
4Cr34lIm+gcGI+BWYIoaLNFVZBQ2bGejv+HZR99BOSmNk9Wy0yvRHQxIwYq6hdsFuqF8qX0UykhD
/DzYyeKFe4KKT516YtS1ErR3DOsVFoGTZrxmhsZvBOe1Y1iAQHA7UcYA1ueySnKiLpZpYpWZ/UJv
OOZk1IkYMqkDesFNtNMtUV+Bd5ncA4h8mlkp9Y+keSpWieeqCwgXhbupod25Wy5HMUfv/6SeeVFd
HpSh/iAXZowFauk87w3UDOuXY10ldDXbu48pNOmcjVQB8Ecz4VZNLG1InCTDykugiYnlW4C+v9AJ
r0uExNZDNr+MyrXh2WPaJSpDwjQOD/Zgd+u78xe5sXk8TSipst0PrOXkLMkpCU9ShWTRbhdRyFpp
BKLUU3MiVGsfTiqhX59SHAaDsaEwWFglrsw2dTxpLX7pBDuNgJNhk9RzlgX9XalHZ7oxNZYWUSzn
dAv4zrgzpD4EYYF6PCEx0MilX0ydTOx9atbbX5xbTi6G27I5JfKRiPn2X94hNNR9Ms2I9swLa5eb
tOzQepJ1Hb71BW8CMR49ZsUlYFnGQ8zCDfcWtmEmxH9hPZgd7DcXZRIx3w2TDCrBlqfRYWNB/hJC
fLALodqlA5uO66sBxPTYUwh3UsLFM91ir0Yb70m2IHV8E1rCYjCIu+TuVS6EtHWaU0fPkwplNMlj
DPPo9j8XKX4vdGC3HHeUcyECwuRFLtFUI/3Lpw1VgzbLjeWbCKTwJ+kZJEQTNZudf19Zds48ESWo
2xs9gwyid9Q/mIIjmnLqiOpxqkTCGW3H2X2C2wev7gm8mkc809bX1mApkOMothqBHN8ywYGkOohp
XsCBNtNpyuNN488MFEp7EeWWrGqxGM8YG8u8mdo3tL01mm7tmKg4E5UW4T24IT1QO2gRWTJbZCPt
G9+g6QREFFl6osRPAiTlADszp+gi+WdJ5g/SlLZl5Ha1ULxl0ZvxrrxrClu7NYnSFYkSG51nqFff
aDpcoXJcgYwNpeWp9WoV5e63VrmSfaQpkXnALHJhgxogVMtlePCSl7yaEPHeQQe8Okx3hnhGPz+I
yxnkl3QMx/uBY89IueUZM1WZ0i/kKa2tOWThHoz0zRlr1UocbQG3Ha9fgkCSA85VsRimdwjBzDr3
2hrZtHVgCk/toU1wYKVsoUuxgKKnnvsLEwF5+Kxk1oaSbJQwWeEyj5x3TWXA0RUucoEqn76zqPuL
t15UTUHupVvNtXMwW4PfvuCWWCsthMsd0T53axgE62ELkJstMyh84tctVi5J69pQTz+ZfOzZOSqY
moGP3obBnJ+8e3FCSij4gUJPpIMwUvEzhIMesIDJ26To6lL9MKUy4E+kmpu/yAKct/WMjokbnUYu
6HwdHCOmIN0YrJJQEQBwPHxC7OvRdzlK4hxk4Sm5Xueav8s2XGx65pQzpm/nDnqaREylwA/KGcq1
aZLmqso6j0ODKIlyvpOGB/nuJ7xGE3zomhj3q+M4Lz4BzUFxYonmannE3WzLSnTy5OceqJLkZyHx
R9DLadXm9TikonSXWPdF7rv49McVqjrSxlxZIGpcP02RTVy0ZvD53jlxLh9DXYgibgTJ3Y0fvBXt
3BUAJbgLNS22h17iGA8EpWkdOV0MF9Oj4vllg5B5hz44cWJDiF6Uklr9RtBNFUfcNzxmWuYZLiIf
9DZ4pLj1hY+/PCZNQ/n7udE2VQZNVfsfoNVOuWIP0dAKKkS1U90XKzBST2BhZNQB9Ql4QE3Qjf/J
lxyESon82rO1sufzbyurT00U6AxbScc0XmhpiyLP+kYohk61Wju4M7dypDqugLw7fLsnCJCHzaM8
da4iTBrvmgouuv9K4nqn7mNKHETfGfMa8AVGffTf7lK4WbTLffqxYfm/tirhh9m5f9+GQmEQlPv2
eHReH7GL0z3u5KyPTEXNvPY2J4vPKA2gRZe0LoE73wk6I91NNXqUTv6IJskMcf5n4qdFVuNZJceI
rQaseWELwTVuJShfYFyuj/6Hc7lOGsF6UH+xRBysj+9dhWWC4RV35auvSexHopWBG2tuwmst35u3
MmYmSsWtCNIlNGRTWuhoAV6F5aYnURyRY1Wm+/0HC29LSt39efNAGektQbx122NxeuXoJcOcMf++
/ptmbX805DtZLqVxYtMNB5774cjl2nZinn/keApC2AiqKWLlI6WFuwOY/RFJJMVupw3r8NrmImO3
+TGHjTcpnd+K2SyhpNg4g22w7/q2Ammn4e2ovKxrw3f4C7V43IrKlF6crs9IEBGxHX+IWLahBBML
goevrTF0Y5QbbXaIuvK4hcFqOPZ+ytrYhLmyS2ZDvYCB03v/z0wZkLpl2Ng8EMfNGP5smW4sRYLo
Eqg3so8bEmbAcsf+HR11d9tmdfTl/aE1A/PVWiZMkU5i9P2E5ubvAKu1qvsVDMhQtxO3a201+jgL
5+hQSdnOtGqqNJ6axyQQeD+iDWswpEExrPJprXAlwhLx4RjDCqT19Ka+UNIzRIXKrJpwoRFhxcQ4
k4dHFs6hNCqkM3dgnHuefM0CZ90IPCwtCfiFXrQP+zzeMBvG6c0HnS1x0v3rqsZ6mnK61npqA82c
oT6WGn74wuDrCU4Ev4zEb9iTGBsvzFrqw2rXsvay8UV1aHTtr5TUZPGMq/6G503a9tL7pMmROqpN
f7eJMEJtrlTqN74OTwIzLFKif37cwhPv3OncFBhLiNgfE4QbOH7Y4010O3zOWR0yZbpeUsJUEVVk
ra+IGR7Xev55y6JRuwgyXbBp2j4TcwzDRiPNMwtLWOAN5oR9C6WblrQoC4uzR0ZzlgRe5jvz6YJA
QapaA3KjN8DgVNxczT/Baw0mUmWQ18tiMT3paIelM+/tLQ+IAcwWSS3vSf2ceLz0OwmYvBcwQAWP
aDgaQWphCJGP6qKNtUwaBmfOPCTHaFX7x6lfFWk7tJdemJbFUrWEN8QGKOWrlu/orrj1+IMDXwne
H8nm8SbGhSCPNdMgYwThGiU9n+1s5nspoyMZpKbBKZFyjoYtpt8bl2UKUB0YOIHF9ZcXFvkIZTad
c/XQl4VtMatBa1TtByNFOK/mXzHwHSkqHv8JMfa4gDCJ52og54f3AX5H3BNguRQS+7+kEgi2SqQB
wqQIVzJ1C1yfi/9JLqhF5nW+qFMVrmvOFDTTLEJH1Ts1Q4+gwDKE5DRys4d57rrkrg3z4DGwG6Vo
O84npiwAL82/J8opXXRkh6mCldJSM8xK/i0M5bIng74Txg0IijAdCfL1r96OwRAmxucwRMUFPtvb
VCzorj4ZOGCJ8HL0KMqIG3EFq9+LXf4X93GG7Rvh52G9CLPLSRPbdBEMtgkOxt/e4co/8Sk6ui0T
3zcF1Qugmjj6YSgHU8++tooE464nu8niaZMzJmktcTV6s4twsM/JmSmuwpoq8JElnlBhlr7pIhsM
CgG3YdRYXyY9Nl/f2cpfzlLiNFnQP3zAmLWAHwfIkIc7eE7B3djr/EtfcYXMXHEicinjyOoe7PMc
58d6bP35fxCp6gWQLwi02v5ztv1tXIiVzYWWn/xpzB1zSEzVtFdBIkL6a3BzQ71xKWLhlomH7qci
vH23jTkLqrKlvML/4H+0qhCMIZ3lZDyCuOjIWJL4Uux9hW5Um6t2njdDmn33MkOsIaAgq8JKTrCs
+nsHr0e+JHnhoMWQnlq1hmHPJZT7MNrDzIO81fRsJwtjxjn8C5zClEE5FEIW0A4EV4OfYq0CL/HY
NJ3h71WZ5Kn/fsOY49PL+m80hc4GbYLAJ6DLPK7mZ5fnzoVXVTPqAg6oikCaP/gJ1glcakmI/wGT
aQsC9rrX7wtnveb5uCBTsO8PGxK+tg+AxoypJAUQvAYSBJD8Omj6dnhoko/KKs+PuaZ6jJiEK4pi
7qfh/pwh5VvyQiH9gC4c5wRbb5WLgZY6UXaAIZ0BcgbSIPB/SeYcganhKGU7VgaTcL64M0QAXY66
/JtW2qp0rK1b2x26uwKP5kA93VGzK1yRghi1Vy6tQXeFnQsMpPZQTf6wqwOx/Vv0kV0RfGTcXIvS
mCD92Xiq92f/wzojStrumXJtmlyF/tL3vj0TZbv6OrOhaPzUPpdfkfA3S81Ktthbb7FujbsEZgUG
+RGbQjJ4Z85tyA2S2FvzLcmR25thOLnLAJ36n30ortVBIzXRyv2LSOPYHzNw7M5ErPep+Ijq7ae0
H0r+rvT2nV7neATGpjIGe9weyS9QxznA53y+dpXfnIQxbLR7E9mvo6zO+oe+tNFEionB1dmVH89O
oGl+nf6zCUaXTrv9+83tPBpw5moJbsOuDifOw4Yhrccr6hsOSj6tUA4I9rOUjvV+bceb5l385Z9X
6nCYF2iXVBYTOvrLcvaNTe//zZKBTdMn8LuU5XYITjRnAMQq+klae0ohRR6E2c3JcIissC2TB8/3
Q6ZeyCAAQ+8FRDEheubIpPdv4jGLwn92QRUHJQ5igQ29ZPgfM0i3mSrTdEPEYRRPor7C6T8q6634
7gVz6wXW2pp3NoDFHQqss3kGr16RxSo3VSauzwRoOXMOa5k63Q1y/UqFGEJqNXiZ2QWnFnf1ugE9
jhvZ1gAA1+rv8iBMAoXXdcHZHxfMFFlQgwZVIbrLEfmBiJAEQrHYByvUoPdh5ORqLpAxGyCcPDvf
YQ2rCcb/bKuKcYGaM+5D8PMlm2ol/NJH9hZ+pKelzhPNv6n3gXsXrSUrKdht48ABFGuyx2G+DA0f
V9CpuI2ybfTmFpzcn7S+NZumk+t9B2uXJTV/Zc6eOjO6lyd+aK4EkOy00QzXpCPYgbkqW0PwEmXi
Ibno+BbMKGJZEHslD+IL87Ze4aH1Q6Fdo15Iap10rzA55T324YHnVGSxTOO1OBrsPwIdOBFaXDXA
qXE3dB8eqvrPB8kFcsH0wfNzMPpcP7TAL8+aALm+d+ME/kAwB3O/qkPpAmUks0ITJk3T5Rn2pi6N
1OLi8GY479NUDvzqoMs9CAsLew7ayU2/SF4n2UcuiWhcil/rn41XSqz7LIJyYBOEFjF9KOHVgTw5
cgZcUb/98crUAFha5jD7PUfFkQ81bOKkEFKJc+7d7HJaUmA9s49e/ob+Rme5RhiESnK8GlZGJpIv
LbqLqxu3iJAoYNVLaFS8odaj1fq1UX+XFUIeqMcp1mE5swjv3DmesBaGylZuApqgj8dsIxTV6Yem
NlAMgvqLZuVKkfynJxYhlTGMSC2uW2AL4pb8uAcgrA7xCRxTkVnICecV77GawKShTnAVEpRm7jCF
2KgBaG7KoTOq3ktHOrb6Y8dmKaieLDestB55cA8KqaOKeAwnRmngeQjcPrt9+nG0MoXUtKLOOmsg
TV279hZAWgYvwkNyx6xGae/35l8NsmMy/yUgXIf0ZAoUk2IapcA12gYt0g1pqXXVVvMYzWj/lsIX
3kH8VSxwwAFor1384F0WfrgttnFhdSOcd8zJnZED53BWJMX+r5o+BxHUkzZSGneBsFf2blfUJLrU
k4rsfs0KebzIyzZ+5sxpHLKI5ASusYLbcx+oaHgqfhV2zVI2FVVHjUu0VdB7xi/myexo8cJf8J7X
GfxtcobZO4rvim+8UtoUqZXNf6rErk0d4FVmuHH5x68bUmDReO0j549euwcI14RHvY1spMCeJ1sk
emTNRu6bAlrJ0CXUXSnX1YOX16LUSTEpikAuf0gcrB7vbhCZ/9aP8+TgCq1+PblzNSEE4f0h90q8
GW+B1+i87DPmxo5CQhgVlkXEhSGl1TB4TifkSa1/mKRmeOgx2Ql+qLWhzIgrO8UBGq5wtJLAnyvW
2UL9NduvCbDjJIfhqOzbIrmQGOTsibdciAEn/mHTJi7ZAvwwPzrBK7rAeBnbTgS9lBfs1bsh7yIO
yYlR0eKuV1nYhv07dSdJNwoHAZnQGbY+YEIjrRLrkto060rilkQLwQ+esPlSJa4Fv+EtXvCZA4rB
QEnouz2Mc7WQNRqAKnoRCb5Mm76ikSDoQk8oE3xj9/MbaDHUPm4XwtUoAZS+dtcwtGmbAf9SX+fF
6U06zJ+t7GYBbkQC5YYBVd2lgOLHRr/idCnM4S+L6dGJubMsMwqdN1wkAPoD/AB+Utfjth4MJkxA
P63sk0IXGqEqMXmmAzix2iWpbglM39a57rB6QR11ZI7yU4LZepnrYPIesVkt0EuPI52Z6C7AibPr
jOBFApt/IUZgoWJHCNYMYJmGLhHZBER1LXFI8SqLo1baREJPolWdqXxbwsb1k+0Pq80CpqCmXww/
AaT3H1LqdLiWmLuxe/RhlWIChMSMVh4WWMu6sDrry16FjzMuo4WVCeaWwPheeFBNwtAyfdWy8Jz7
b6eOWfJXlPXi/i7QIbJqWQGCYyPpwKbSEBFS51gQFyVwuaaeAnyWGjKPKDRJTdRByCd68u8UYI6M
tfoE8g7ZmdCPkftryAx0oVSte7lYGpR3N6vfAgn83Y+NDrSbN+f0Rh3DUNIfdU5TB/mDemzHdpLi
h74Gjz0i6TSYiQRqWLCf3KZQ0Vs4nf160JzpYHRUyDU6OCipyILPP4pUWo8F/6Dg74W2KM1HGFIA
y0vfZ6BHj/KxOlu3MWk9vLxJpvv4zLhqhnYdGacHndIZHJ3aJmviCRr614EiRsX5hjEiTgyNOjm7
A6t1xyz08/mxppw+OvRLUK227eTQAmdYun+Bf5a/YEsA48QaalXVclZLYgO9VFCsDir3j2mnoFPH
mfm1bkYs3Gv5yuT7DIUc+kHuNCaFYcbe+9UHkA8JCRIFHQz9HfYS2Xarh8x5kk5ld/QSNOdkczw3
b58KROYTuH+R02Jy3Uo4yt9lwRdf7+VlFEaWPXz8aRFTdd8W728+TMaqT5/QCNqVJHSpdwrzc4/j
AQweeo8w/sRqcUqUnaeXJX2W4XqsjyGmTyEfZLtdbYCOUV06snoRGrz1CF6oV8lQZLAvsTgFnwU3
2gWFVKOEsyBLEtR5JO8cG2XRqjHYHAF/+ns8bicwYWmPyp5HQ0xpy2kSJ6n5+4OzD4SVgw5e82vO
Gqt18gTKcUaqfTo4VThLlSSDtMnr5s05kCfuxs5R91pxyTyRkRviV/dDRMdSbMoy82USmB57rJAr
SxgLM3g685vJ8BA4xmpQkpJ7yfEX71kCw/u9mGmUsAJEBsZbGMxYUxSm2Cj5fpDEqOSUgf8EvuQX
RGVjEOloysP56wpPxJ0FE7PLe42npIuY7hA7+xZiWI/iKGxoFxaaRWswENowhC/JcHRix72isbL1
riGTzhCnY7keKsdvi4zOE2OLsOpA94MPIs9bDddT0nmyGdElVb8403yeCJLSMQuRgxGlvuvRxkNW
wykyZoRA3FVBomxohpQaVUqCIgynQ+QFRS2NeJ8fj1NMyzwfphtzHTuvzENxWSI48GWJ9Zg8BzDL
HcKiJqnUG/WTpsJil9lOOma/dgxsaC34CAWM4bOLEVCiWsdYdlMYY2aV9wH8SnBclPm/MpqPG9Pj
EkLD1CIlhItsFR6va53p+LHd911RfwWSCLvrI/aMd9iDxRYefg1bHPSZ4gvis7RUQvMtgMwWgqIo
2Z0Z5EW/tIzk4FIOwLY7uJs7bfNtrrJ90lcxwhjOJCFLZcUp1QQGmwq5KVfH5UXAzqx7yUEMVd0o
kbT5MdEhrJ+zAo64zrrEK3u7PYLzeIdd4WuAiLnBT8znAXrE2wOLVtTnRovGZpkI8Lx2PxMCNpqt
E2ywZKItB9w2HhOz8/qcCK07ki16AuJB2I/2YSSdaX5VsTG18MJuCXoBOLHTRRLqodsGBqHWG7dU
X3iTKPJ5kdYbUzSr8oYzJ5zqPxLaaJMi714emryU06wnnI+9ZGswReKuDBsk/t7flcst1MfkPuc3
ljCi4gU90+ItcgbfEqWVUAN3VCftdmksD2HkjX51YctmDns7dEWg8YyHmv1NhJwOXfZS4zEbAqeF
QRkvf7VuGokXsE559eA8BM0GLekYnDRs0SlW/cWTvrvV7cuWRfHSUwoDKZ8hU1GueABsocIUk4fq
Mg9Frt0fR7t0rTfUgTBPX7RnjCbORcpddUmZWht2aV9Z6OJmy76B98iN8j88XFsSdpQ3u3mnDvQW
4anKxr/ut409HlZw1pZm2rYXhNDO2bkfKHYr0G/ZcGXfLrNWECqDNjGFClQeP2HwF9Hv4CLHwP1g
zSUHYp/Kdl1KEprptyPNogm78QFiyA+JoXylunNnSrbMIjqUOif3HrAyqzzBvDQTmcRP0ui6WDGR
XGKjQRYCpezTBW76UX/AeNppznakG7LJCoR9JeKuI/sLywcAPOYcs07nexs/IBpNOsu1xI5XLpIg
kPtj41Cw79gQ/eRJyAeCSoFvFjxvBxXIdSjzRMP4Q3Yg0riDjrCcTNOvyzzJ28f2bKP19p29rsA1
tRzQBzx0Zqn+QQESsGdYqaWxwiw9xdUHBBAcPnJlv/i7kUzjK1Xs6/KmANlwHP/e0kCBS0rttQcN
M3WRlCP7ehrbsw0FJBFNgCVm00WfLMYjYrFcrYF0tz/D2kTcJyAEHO2/GoQdyASdzvFE39paUVqJ
f7m1u19UlZurKdMRswg729eNgUwBAmZ7WSg3at4meeGnbJFheWbbhw6EzzxVhL+FYeK890mXIx3M
gckaMesFISiJKRhob3F/myezOR2NgZjNHsvo+tPQ40fpY/Ao1doyiLRgcgcS/IUWM9N4h54vI58m
rbFB78DLVlXlu21vb/UPUjWWBYcvemdZTu6TydNqROSl2pAjUN1dXy/3mmSPdPoSF91S/oKHwefp
9tmL/RrAH+XKJY08QDVmXnmwgOtkcH+hLe9YzOEEWzGb9XVwUoaQtW7hZlI0FUY0APEwjcVjW4YX
db/zNb51VcK0pNXFfabgGobZS3ZtAHNQN6HmdIxR4OVwJuDNLCLhkLtacfaIZ+jOkgiTfBtvfTHC
yL+LjXBjgk3rk7QM3qpdBid6S7aEM+hloIm21oCuwZSKx21ly77iUkbGXPPj5/KaUXAEw41cmy6+
JozU1Dm+21xL8BNlaCkDqFcas8/KPA5w9ihnRgs4iMYLksPIO/4i5C5eQzmzwr1uOGHalsaKsB5j
juPd4FVcZQerQOFxJCND3L4j8IBlzDwiKL05WMxRXT7Dswp6NeZwULSpBiMJM+wA+AbUrdfc0ixa
peshqiuZ//tg1tdAI+JYIFpsnKjHe3Q+oz+S7byJ6eVM9n1jNbjdTONvkwCtIkxYik4znhQS2AWJ
g/zqbYKX3Xv4x+lV6xYxVJ3xxmILBTqnu0+WIcCZS++6ndQCdq4rUIraP+NKtJtIh9HA12oesXNl
Ms+Yttwg4fR/TdVcLTbER1hk7MEMqSEKXq/DW1gr7l7sTnzt9+kFFJuBIgCZ/DZD361Yym5cBRob
CAADKiY5jYnV7pGBw/HhlcVI9BD92Peof1Gy+IyHuzj29kheEdu8po8k1anfU/rwRDL4SLO7bqD0
1ryxMO/e2NOCNfNbdSadLrknDdpr3IdR27UZya1pBeDx7BpBOhdxAYha1nHbveMkEeqynwHFmfYG
/QjTY0VTdLfWq7+m6sMZf3qwyz15NYbAwrK6oEpweBnBg7ByvBftQKb/yuk4CEQW1jtcNM4Qt01r
GmMSUy7fwPt2XINOGv9sShPeRm58uD6o2NbkDZ3o1v44Y5uxqGKzykWOPKcQrf9jYOnYa2I9pe5R
f0MkDmiOFmpXycnOFe62vF7a6lBJrPyBibC7xgJhQvJPFZ5z8PDAXFQNm3uV0UmmJdwj+hhLYST2
mjtLrlcZ0ArwE04Hd978Isbw8z5zeOFBr6hYnWbu2+v0kh6TI52sWOV7wlXzhUaOhgVdfAcCTf8C
Xb1Ntn1hdntTZKxSlqrIiWnSeP9E7fyj+u04ThJbtlwUkfAVrze5VouoGBqG9ySFDUaURkUm8kNC
85uKsYocmy6nuAwHTiZsm2UjW1Z+9Ykv6xBgmTiwZOlymzjOVkk8JO9kLVRP7waqn55m+Oy2bnUt
iVje8nos6PGSr/Bt2D8wvfs8YLQmVnvV3J/PRowjvwmxGuVIBdCPXTdu8WQctK/MRG7xb6kz6Nv1
9bysZaXfiSO7AMvzw7QkcR07e1WQO2VNGxiqpqn7txA7RptnoV3ZR+oldMMKv358Z1gPtFtqZOVp
09WfEtMSYxBxs9MQz+MZ+/G36hMfosFyVMiz1c2mRs8jPAwSphvPulGegILKEzxr1KjYSvlj49km
/gYbgtYlcCDFHIC1GIrtCycEC3uXSWx+eiGyNDAki4umXXQ0btOFRDTtzMWaktWfigzNFafdJJHa
cdtotKW5ur/ugMmhrWwlgzoOs57teoyYGjicTsiFZoyBUnTgeS24te4a0I7Pa394igEVfds+nW7p
AkpX/tptO7PzeKQyRIwNW2PW2jX2eIPEulyDdJLwlX5aqSF/TeDBXxukyrq2kYsI/lT6t2HmvaNT
QmfU333qp7aZjd5l1jt5dCTVeWwJAqiVQANDvyPxR3rm4txnDfkv7B5lAyrxnoBxuCEuvZD1x/3+
OsORBb0Pn0WpK5bZmW0NWI30R0P10tOquM1dvfi31OjWtQHU1oPEwBlWWnSoV5Mj0iaMlRtC4xgA
eK4b44clYBTJsgRUxdZbQCzVafcwF2xO9G2nX10QuAV1clkEPkDxWWl1yk+W5gN4oQPoUepWZTvP
uPcjiLuxqc//cSuVVAgBh/DCafLvcSEHNW1Ti13iiNxS2nUIV+hyXuPEBiF6N3HJufGtsqtnIy++
KVggp76c4kPI51HX1XK2wJGoxby+I67BjK3a/4+CPxblr69lpx82czuwNIiD6FiZv0hUIOCT+WSR
SLx4Jt1k6XRk8BNj3rvzv4ro1M39LO0NHvdi9kPwGSemI03pajFfTI9aJM9kt4MYwuOI4hVJ3agT
fozjkyfvcFMjafQ/sj5OihHEGBKc/nunCt5vnnZmXchwgB20Fni9T8jk2ECbUKhPCbWfttne7Pqp
cSjY0bNG6QC1sPUZ0yHJsHjHFGR0w21nceVP12w45YD5IhJxnPDdYI1EClz21am7N9j+iFRjCPOJ
ZgEAEvH8HSTa4l+UR1ZCq4AypSzch5dXCtEJcfyGvtF6Z455Zvop2nZ9AIRPQbK9ZbzJgCiJsmSG
plPVeubxqS16AytXOPP4WEeVwnOMkLeUkeg0jn0WPNtviG2OuAGbUfpXVl2IOyT+7qZjXa/SqfSu
EZao16MK1NC6O231rq4/pnnDVwS8ifmsJMO0qJdsqaEkNHrGSuGjntTDhoHkKP9G1xLvr9K4TUWw
namwgfZX6gfFw2ViCYALZaNpFz7aeADi6xclWQyoGEOrliiL7l2gT6JC29VY/tUqdWXb+OlO8m6N
lkgo0i7qfHzjvPdyjH63YzKLwdXSDSm2zAqV6SknpnoB29pwvfhPLXp7rbtU0xZMgVc/UwmFWlsq
Rv0IdGJyNS1jiu7d8BGOVaBK/MYm/XSkKnCdqYZtxdmKSxeAoJqbTdAbfWoHCHSh1R0a2uitfSb9
jkEurSmaskvW9Vb7HRkVZ0LWopD/wWvUWuUvJWDBW3rTFAbYySU33/92Kxm7wAVYrdHC9tcQvpaz
NkQBc02KPEfT+sy9eGrOTxL+0dR7zQCzt6IoOSt//icSj723tv8sJ3LWduzlRcT9KKKOV+J22o1N
b2TseMiLg5sw5n5vf54aEG2UCS0hGLNLudkcqRch0E+8ex2cH4eqvY24HubMlA8lNngT3z/2/08U
64gx6dnDZt90kSMozPQG9SAAb7AVKzEnYjnosksM7Hwjx1LbK/0vuzcwTEctFczRsSdEI6utrrBG
F/g2BUttyy42VmjX9oaDqB3zELIUT+5yUfxZ23M6wiIOaXF/fXo3XSE1f1S63iHuLHYF+utVmNt+
jtRt9ayMpFcEFu/m23LXuuePn5wlktiU3tG3gv5ptS8ocJn4ivGQBjugnE/yI4V3cfr+IlQOvnvl
2QHyrRpB/pRwXEc31du2laj/qbHfhPqcZJ82CNHg6lVumMsLTzXjCGfu4AvSp9PcmZXVXy3RtRS+
2MMVZlhSOadbHbFnf2aG1qk8/QIfTXIIF1M6NI//j3pVnXHbCYd++pgGI1aCNUpmZKhzii5rETWU
dTudzk/ziX7RZVjxXTuP9SuOO5n1nDZiVdKALjKz22tfd6GvXmZeketGbft9SkVt6ZjiJwwl9xvY
cTc54u2DnevBwtlAc21Z10eVAb9IfLbRZN2LQP+cR2p5sHKqxlhnlkgjAdEMfWp7AvOxjLfARUDd
fsJaYRDZGIC6X+kHmci2nmToiEuqQQ1CSYiNfYO9IJy1yhxelMAr3m9zgjARwRoz7xjupluQ/U1o
HtwCrE7lfENS6JFhqcwHTZiE7BedfyXxhBullZH8Con1haJlnIm7627v1WbmMk8yc26T/qJSZtfy
vzz/RokdGIvu/AVtFhFONbQ6rYDFy0iZOYvyHtSS0oGbkRmMHj2wbpWqQK9vtxl8QevNko9iI84c
t5Yl5P5nyyCC9t60BczD3HguNHjIcx9/36bFDqhYLlKju02yZEh6YY8TggzK5K9ad3swtbRJ/OuY
G2wZNxtJkV8n/zIPYSuTsuxD6wgRA57kyAZVWJZ5hDCR9JAGEJbmfpQ3v/KJNJclSdsm92l26MUf
0YGCcutN1JNN/a79K7hDNm5peQTNJUDM9ABou6+VUb22AZdxncD0Dn9kVhlVMkA9JcKElbrU28Yv
gVp274oFbjVqKt7fia2vwurKIYC1pb3iAbvFiQ5InWJJ8c/1yT3VffP+VjY6wGbLKpPEPD5dpPY+
svWU1zBm9IYSvEk6Mdd05Tv5bR5LDQpaPrQFfl216VHOc668+lyRImEVEc+oY7XqNbvM9dFKcwNe
ueHw3ND7ZApqx2iYag91lfKIdo70E0EJxonjb426YMUEB4pI1ZV6xDoVN9svt2XNIDBwP/J2aLBF
LXD3GlDoxHYomdyA/BSMHzAycSqXzk92eMgi0gz+es18L06wpr9YNeToP8AwqiDrpVHfAKH5P+d5
F4GqX+ssm5M93LBgWC27/QRoO6XsrxYB4SE8ONxJF+MWlTBW1TYxAetZPrVJrD1/p3kDpRb/bFGO
sbXobetkr/fjQ9gQJ9Y3/LoA/UYTdfB8s0guzce1B6cV2GxHExDwla+NmpigvrWK1I63KmfaI/A3
hz8GiD4HPrFGom2SGNkLoDfLx+XYVPCr4JJ+QiE2CFbYKaCQGINHrT3DSajNbTcAnAocxcr9jd6t
9CNB+jxVl7SBv8TaS0Ro/+67kG9piOLEpLSaBdfPMm55z6datBzNVOnUeqTSI7ud/NRyZhIeHZRD
ngHVARQJGDWLA9a6/SauvJzlkH8LdA2L3QhNb9PFkocaCmgFDH1K3ar2Ci/kDI+P7W1DmgfYpg8d
TljAk7VV7wP2FD8ZZBDUWl7R7Otvs/RFFy06/wq674ox4RW8tUHLS5/6CwHV8VAi/Ieq81rhDiUz
Y4HSNwWQpMXsN7atGNAmgUMDhZ86IRr8ojf0LYy4N0o1V0eNpmaxYzFtRZCHto5IgMTzj8ntw89C
Qopm1arMhRhpxZ4nhMlsRBGwdjcuTLF/6tHrcoWoQwFCie+Vb2/RwfPLO09dcAQMux0iitO32pI1
X+v2hTbe/JwiO43psrJgmmH/hypmeoSNz46uPTF/QzHyNQenXGjr3V5XtDGc6r3SoJ7yi2mp6kg/
6noTLnYi9myb9z7JFOZV6cO3nLUKDwC1mup+GqW3ebg+IZ6pnbrJuVgjVaPGUpyzJTlrrVRCaKNI
RSa+/75tMUXPQAwjMWqxza/0OnBhkL1lKHik7xhsn8UlKcz/LpspyAP1t1bPRsjLbY8tJqGRBi7o
E/CbfvoJT5FAHR9vC1q1n27eUYX5wWZiRT8SJt8OHJOLBdReqOI67MwDa3ky+ihe22wiU8/UJBw0
dixt+GP/uAg41Zez7o3eBqQL85iTGYH2z+5wMkD5JUGaA2AyIVD29597hKKROu8IjRJ2xUOa+MHH
csyEyqhgIqYWaXUZ3lLrBWpNoZO84VN6gXCtN4eJ+I0JnNbh2OX+ktGvwyKaIM5Ctc5wrIaeDDXc
Lx3M5GUCjgARSVl6iN6KnFmjgNAxhdSzI08ZEcASmLp9ylV12lQKG8TpYhbKAYkmfff2/BKkbRHj
7WZuGk6vP06SBsFcgezJp3fWFxOFTWZhCfG+lKgDTC6WBQlr5rTKSG8kEvvXyv0J/DcR3Jgk37p/
DG+y8RW1TDr/DXc28xsqsMuUa0HDqRYgIYGW03dQ2VEWjlx8el+ZZEzDp3XRWByHED+brWx6cm3R
zJiQfWz97iU5klHMFeD4OHp9NKqyeqIG+qxmOLTuYDSqF8RugIXvnWByOJPE9yCCBaul5eIFXhZa
BJ3IzAaqMwP50N51rvE2tg+SazaxezlIZvacYtmTKl4z1L54/X97rJ/ty5Sx2fXs92T9N56Sm/qp
ShZ5bqj/4UmDd+gMVZU6pAOfqCTadNuDJKGuOv4DrwVDsaFmRItrvAUC6i+j/UilaYGj9BFMeG/1
lWeLG5PXOsYZOqyhLxSQDiEReEMHlojUbbAvW0CebeFQRuYoa3f9STDl44cSjofyQcFQ0DlsaK5/
g35r3PlvCfHqIDGHdfSjLoZ+tbOsAU1GFGyPFdY6YvE1476I/cd7UU3CCUVS+9GEUWsz9SaxmQpV
5B7tshvIee2op8v8FP5IgsNTdu+6OS6ga46e1HAzBhIkWfh2b6FyQOlHqISKzIzkrSSJ6jiiA2me
OOE97FEQzq2m8aL+KLqGIGu9TtjImvhLA+aTugZAYg1FGso6skkEomYG65Rebnbm95aRfIZUl74c
FvR4GDNTciiWKgIQp21Rhlv9FLjTQ92/pvPJQR9Kr4BjvpeDc70q4eX8azndkUU4ogMqkx/iFOXE
flrKCGwHzrzksbpus7/NXFt8gbXHICx9JHDVrnHuXjRUj9SkIW/1mXT5fuenThxum+gHIpIXeOSS
1BUVy9+cD6PHm+U9F2+F9HOd8OZ3rAjf9QAdPK+UPELojAJ/I5SswJqZVzef6TPpeCXrCop6pUYH
ZV33RCeShXQHKS0NQ0he83UuD0DZfy0Xih6G0QOTEXRdPR7wKJTLQi8gzuxnu3LlYkIWIv203l7r
JMlZixCskMYUtRyDRkoaq142u0QjViFRGT09xWhdyCH3LWqd94ftLEaXdzs+3hY7Rjm9RaBmiDSD
3h8RpiIfi91Vuf1rg6YMLZK7D2kFjlXnGVGGYCnpgNihIwbYJpSc6J/L/BZCjF+j5ktIjTjcKLQr
3Q0nILUGJJ4tEM8zbkCF/zzpxI3DdWjZwhqe+vgWlfOX2aA0+3gH1tYc41U45dAnj2h2qj+HSQLD
gZJ5FUmvMw2Qin45KFVEd9Pri+W2O+3QKCxnej2HiRg4hWeSBZfU5LKlwJDUHR0vhdwEfZTrktOI
BGiMZP2DFnGolh0caxawVVCwF7sYa/MhB48YT1Q7p5ktVcn0s+AIJYRsX4JrARN/AoiJEGj0mUgc
tkY3VGpqk4fbLC1/5Nkg+Dmuo4ET5OyCK9v7mSNDP+LSKOENnBMujTvM47SemOMCkR0HVK40DHVg
2TKVfu55peyekVryKTRVfL/x0z1xbH9HHw6M6xn3/1tYUgSob5V/4GJj+pRTyLuWdzB/y1cmkMjX
+CldgrzMsb5B35IfZgosziI1Gn0i/xSn7Ip+e79m1wxSh9yvp9GjM4LuAGj9gQj50pWNJnGnEioV
GmtS2Xs0ApDS8T1ZQdKkZn6uhMxquhADt8A28vqwTehGzLWhpiJ7ml6upfnhs6sXTyXbvjIBiH7a
HGJmcnxGN+NUCvctBDbDjeqO8mihqIqPpQYrMiYRcBGZZi1OozRY5FU3YT44oHdSd1XEglOrU2yR
NS+zyMD/k/Cj3BgZUoA87tZujr+VFykh2J9A5ixKx7bJ0CruMIc7mmnO93y0R+T7KTrzoHzNE7WQ
opbPXMp9BlakSxmqslbbZYr6304k69JLYrn/aExE9/05QLTNkgtYfH919zzvtJDTBodEu3EDuR6J
6DQh9Z4/YYz3SEv4l2KGEkOWz5cxPw4f1F+AgLL1A6KU7Rh1Y/XXYr9AqfJkCfFewc1g6KxxPJa2
orJ8dFcGQ1Ke4E91VmJmwmLLxYEggMxQ7AWm7WeRKS64/6W93WzqsvhFLepvntao+HYFO1kVXhsC
9qAFDcVJIqVvw2VlUwWHwhbR0yUUFMFod2B16ymduzQsepwR48joz8dqZE+g5pSeVRtbdo/7hj9z
bFsQ2obHmc5FxOGyPqBhtV3HGs5vgGI1fVf15A/UcH7xzXw5xt2Mfh54gUQEE1JUZC270VApyACY
1i65dz0huGGexBoKG7HI2WekidtEPkwDrz9/tc7mUKXdfjXzl5311fru73v8nDkNEpdIprHU59ht
LzUzQa30B3TeqBlY7Ier2WRKNXLdvXUMv4NGvTH7HRaH/hC7pGlHxrkXDK4uOrPAv9gfW5IGboQ2
MMScC7ApiJ23S97sQBlp7Qu978+d+LJ7KBn+HxAMSbu/u7Jg9/8JL5e0JNK9206xWGDOf+CbaTwp
pgUNZ5pCbp2suxTptc5Ua/VEQDMTergHO4zIz/+841OqKLBBZ1ruIMS28qVMBNLkldfKJbqy5Oo0
ZxisXu2VGiKlHZ8nv8SDYHxy10eHX3j/J6kem9hrQoAWFWSvb0dYKtMuqk5EpCHT1nN3t0TAxpUl
I/O/dUxvEkdbPjOOqvc6daO/khLhc0zRHGpIz2xXqfKe5mB5n4h1VrALgRz9cRljmPn5drEU9eaX
s+OQU/OU1EQ7gFZAtzMZAd0RHJTUVZc8xSMFbE+u6Six7m4SwAyjtDhY/cPKC3fZu+QaltDRImAw
d0qkJLH/RWUeX3x5kZd5+HHcm5SAE/Ljuv0lDuas05aaUM33FbmmlIDiXNgThgx1aCFsfbK6ervs
0141qpb4W4RrZ5h72wDjTgMxhM6Ld7gafSg+vDWfFgwE/9IiXUderljtaCOLiKgz29I6933urQt7
F/Uv78oIo71AnRLGjOKpkfWYEwoMoRwEXlwGh+McyMguo9Hf23Ab3f8D5pmmCHgQFo0SaaYKxt0J
NgsLfJomLTKZBqj0jagflWHS7c927qCra4Y0W6pcFG7zb2rKi05S6pX8ThY25IiEX7mEjauJ3FZY
3M7X61ZDI0HtV1CQqDoGFYgv6WigPONUJA6wZ0zh6SLepyVQsa+L5WySDlNc8wsrk5L6KqDdmDhs
VRKHIPLvuZCtOXstT86tEDmLBmCqKZ1YWp5jZBGMSbpx3oZX3AbLsWuMfIJX/DZzVkHXtkHEhTGw
dp3mbzvHAUwsY9BCuClBPZrG1Jzmec163PDmR8vyMLvFwP8fWkIn8sQArHggBCazkEy6TiWYx4iT
1yaSDNv+8TfU73zzAUtnCRGvmlYDnn9iRqKNVoOOAIc8zua6Qx13LWpUlTGV5l8Yvdv7lRnFsFHj
PxfgOrZfEE8Ljr1Szmo/RCzoofwbHh/bo0RSi+R9UrQDCFeDN6WiYYTk1BrddoQbmo5LjjrFEXnP
zu3rUIrdtkz4zgDrE+cIOoUxfejWzIglEieeLZzxj+/TAMnHicai11Jm1cz20kV5IRXEz0coebe7
fDTUvZItHHfUUOln5wgFyC796cMJEIyevNPJsYAp1m745wwqOFrMCI0ZZOJSlzSFNfpTETqUBPBo
Xm6KBlNT367YjBjfO8O4CbcVJ7mOw3C82CUIb4FtOEjgvUUh0Gxj7c+jyx/KEogk72Zx8pNN42q2
QCKwdxbPYj6pTECkQNjSD3+oiQrl089vQVdNkvmBO+yeRDm+HXZtx5Ja9JiQSx52ZnamsLcckyHw
jrk2MDDNc2kBf/hJzuj59UAn/ud2q1rmwosYWo8kkp5Ir8eiUWM9F4fAmMthISVUj5KweZVnPrYG
W8j+hm9PPxLV8aCsAP4HMkthQncF/JBocX37VFTr9GbqcHXiRU+H7TUnWsQJ1HYZlAADBr16mZ3f
ZMR8bD6JD+tynlPxvbZ8+dPZkMg2CKlH97nPk42L1UzNU+701DXNyVaA1QaEYEaBC/qvjdn0FQdH
xu0SPRwB3zlvvI9itu04KVH2dpGcBFsNCJ9+tDpz0TGw/S19t2luqDvOROAhYlUe2LbVG9WwAju7
1T088qwhQ/og0zwkuWIiLqI8bwq5F0R/+lZrYxgpaG0jEWni7Y85fNF1ZKl44AKiVzeM/nMsZLkP
iL52Hjz9puRQcrXcy4RP4D/hViIOsADOLy9aM3K/JXAFjWyGqsnQZH9vbyvI3EuHY/ac8VsL9+GT
In58OwK4F6cSAJIQiXj5H72ibeN8w/oqLJAgxMTsTtDpSBuXbyslxU790mmbsWymfMpE+F2hPBM1
CuPYQzsLuOV9wpwaXx87okvNLBVI+CzJP+aiXKIFnjZVGdLUEh6BzvZc0N1v2Vp/pYa8yg1EfXtI
ufxIsc2bA8bTtDhyJYDxzmxnAeCiNph/9YAM/uyQfgksQSyoopoerJADptqBT/SxKma8idPrxUmA
iObZSxeaN8XjnyXj1y/cYpmx+uEYP9UQ6CGDcn8NQaGCNdyB3KM3TLhu0MkR1OvFn00WBQ47WOUx
Qtg5orpwBu7IK6Y9Xf6xgUheGM3U1GE571JY2r/Vq9Ca9hrQSFqZ+stBPrdOSTM3Q2sGaU4TJcoz
knnph15eC3NaOYdmk9gZyWsvYMrHggd9wA9WVXI75QB2cS++zbzLjJSKiniEc0DOwREV1a0ukJDG
MzWddNkPSQk62bzpFn/VAzejrqAd2bTKdTkUQv4YMY1zyqpg/KxE6hFOQzq2BU9SlwCcY54ZcCGe
he5BX3Gb2jSlX4ciSS22eKAjHp1nN1DzeLTQPgiMg3qrniKBDXaYDApStYEE7lZ0hl3LkWfWseDL
ya2wi8/XOR9txk9QkYIZfvWUgF3CkvzaBpNe1NriOVPMroZpAi7AkD4sQ47X1FciQOjJ8cvM9Y9f
zTbuRFbmf2OXMRfExmHz7jXQ45g3m+8l1Rk7XzWMjz7Mzy2g89VUL1uNJLrA5eE7s67SElhtOf6r
6c4YfdDza+xsyDrjSXqqXMIhQhsObsoCChevTa5dC7Z1agpnwbQoue7vSnUC7uB1wTlLbdxDMbux
aZVTK9Yg4VfrmYi64U4ZxbftcEVFJlUaFFl2NrusB2bakbtm89xy8wzalsCxbyPtt9GJaez9VvBL
/H4RVdyFmbXnUyUDHIkO7L38kpQs7/DpfJPhEeKHWT/HXF6HzrEIRerAWfMSGtL12PdoGx/qCtwm
Ok06XyJJUC2mDMkJ36/81grTjaLnt+IoJw7BZPlu40xIZumNRRGdHP8Y89pNbrKEq8NHKE70df6q
kTCUoduXT9HSpBljBgqVUjk5Ao+4ZYVDPsn7DkHpzyOqOSj22E+e/TwV8S3TYOGC7bi82AwQKAyy
n1k9UQUO2eNxRkc3G/JQSQ5UQ1MjGUDCLUbCtjWGd2n3RYYoe3zptFI45M3Dp6R2rFFg8GUUPLmD
04Q4TYxueDnmKBOMyr/RJtOnklIz1IWPY1yGtERoKFuwAHiQrUlHVq+Yb9mQe/Y+ELUVNQ4seXj9
xNCbUyh1rzuKMDPDjvzNK8bfjC8PiQ/MY5aKDNklki5o+MpkU+/ol+H6Yv2JJWg5nPOSOgR0+v3C
9GhL/vK89uEYQ5U+9FZy6B3lFE9X4F6q34LrBQBIeF+TCXfRP+fZyv00WCoRdYrZnC6gQsbT/IgQ
IFhXtQ/Fg0Plc7hUFvm1zMiNEz6Cj6MoDgOFAZkc5/Rvg0LtuC2PqxCN00pXRTmJLbmA5o6xTa2O
8zvIb1vVlBJ/REn17lChNGirp8Djp6aKb/2GrsnhTS1mc4pV2Ulw9ezDY5cpYkXgKPw/9l3Nx1eI
eoNg8xeTt+EOus0SiQqXDV6jwaZh2tyBIxNDbjkl3COSwMcjXdlTU6x8Hoy2EO1DhWeRLIuKZ1Zv
v67TWLgksOe/OLxuhkAmoouehF5ADlQtyDlW4xrkAk+ZnyOCJPoHMOR/BBbJVTvHKxpMbohvECPb
XAMNLYE91zZxC7jZAGY4c28RN393IC92KWvkQXqFtDHe+MoaJf6vJEGc6Cgh3/oZhWSyI7zjgN9v
haCSChz5CQ7cocoNPvg5ygnmfnMcYviKpETtr8Onma+seuLirXnyEbngv89tpts70OAULcAd5kDY
WSugGIOh4GkN4kIVyejNOjhhSH/6CH1ci3M8BZKNPSAMXq49Z/EjtaRtUp1b11nQA7F7EJqhnyLB
yvIan45sbRgg9Tu5Q91+RQrHayGncjlulhT/4UniOwmyo03A5+7wRn0mLiuuqnGvb4jwPXZWcT0M
XyclPgAS+mSFSMHAGocK9IzlryZd+N0nyDnXkMCv7ycEVQd4AcvtE/vOnBGAiw3Pm22EgTgBrdlb
IRKaj7ENXHx+GaMbt6I57CIfbet+/Tv6hMy11kDCcTSMnyGQEN27oozhX3MPtenw9JnzzeroD4pp
wO7tKvdYvM0t30EdJhPOY6tdXNR1TC6HN7gZWXZ9Nds6Bc2PIRkTsudiCPPJncxTbpVSFluIgAPq
3Fx80TYdC1HZEu1ClrXu2Ut5NTK9DM4EwSRWj38jAW9JxEyS2YszI5CPbaq1+UCKxADNnCOnhIOQ
tMBd/7TAiGYGBOKudgoEv9AT8wDtUPFsW3CfKjZ48FJ5QjIxz8ZKO95yLklveIQZColKrAgn+Zq/
FaEy7Mh8XWpSrZxgtbHJYYyMxMIAI4ac/u45tvr2miQio5FCEtQMcWbf3LTUIcDWmnJXgDb5R5P1
I2y8EI6NGgAuwshtEWGQpA6jExyCgqdC9h3SkI80bvSRhma/fDZDxfsphooGcaXR+d2Z6MxavVoB
nLug1lmrvU6vrKK3j74h0rhw/xwgIeVKtN15RV2BupiJljoCfT52IRj8YZAzR4zWOks+fkQhPcez
365JeJ1Da84FOmVI0Bj3xo1fwcP7SKJU5G2pnHyG0dMGAVqMEhbeC4e8RW5W0N4htWhosKjtMags
0aaVLR+oh4v3XvSRsEK57zUSBRfHMHXg1e3qxZy8QfFm4hDl54a0BTMdE2Yum/nCCdqgiDW2bwD/
14gDj1muRZEVnCui+OkxdvlD1DShELAV4og5Dy/GP2Mdh/jq5pTzpY9sjoK/M9wocHdOPCzw8OoW
z1qG3LBIohQgmA5HmcsEpD27cwYXKx/aNR0ctJKnl1k5SuGD9CxyMjNDDGZtKbtEOSBDDakLl39l
V+FyR5hNVEPYmuDOBYBZtwH4JZRCbgMg85Y8t7XKyByR9AsAo3DxEk42kI6Q2qtu1KzB7dCAzNru
tsEJPgq3Grm717Ccg2lW/yhjdzMhZt42JZrykv/vPK/Qn2ZIAVXdKBYn0wsOnZHxCwowBTRFjVNe
4xPLOhBNuvowBHabCJQgkxRws1nVyLgugHcrx2CYeSspfUcxePW6EybJpAuCGQgEMrf7NVyDyVBd
DEuOr8yeJ8jrGjVsQwj+BfyfEPuGoV89HruKv1ARt0AKLB8v9rQsaZztilzJ2DfZMSbVmVyCE0eL
44Qedkh+Fy55Oc0RosIIQSAo2htGINgOM+4p2zQQezUBEgOgHjt/H1DoDcswRq4GPu2ZqjS7cuMZ
GOwdi3sfie1wfdftADCefphDLG+Tt0DSfNRSw//Ahxa++ulckRkWQoEYiGmWHZFgSFdLAMYbvs0T
bybsc8+wS9NQMbveRwn/NsdPZapD89wRQqdy4lMHS7SVcD/ucOvvGuA7yLzEeH3iszDGClCcLFu9
nnT7+18CyB3lmJMe9neg8NuyULvwr3O5w4ez4ty/bLFlfjvxNoj5FTiGMVTqmMuqzjwQH579ujrb
enzpDOB/255XzCAKhI8/tBjgFiD3aCj6R+Le1ANkCTP3L7AlZuuS8uo6SYCKE9Q/3BRKg++hDGyI
TO3YYT9u4sVLmm7wYxMHq+T+296IraV43qI0KIBJsxdW3TZfbMEomwzuEFy4Gsn3ZRxHOzygj0gj
iMGJVWxdXdrlOuhywJZxMI2kp9daY+6crUop52uo2/rBA2HpmTbYspIuHDCm/zAAg9JGeRzozSZo
MHs4josJx0gv3WQu54fbkMRq4y4JFuccPT+UiDX61prqObWez+5mRWfuwMDKOXuH8Uz0IQL3R707
n9v5chx+tDekX1+VQNil51wqDlw7fmxl92SNiFaHkjdC6CIDbVeU9LpScidjRZfniibQr0DIwdzZ
K49+4Nw/lhbTwlwGeOzfoEz3yTNq+LB+Aui7E2XPKKiaQekRvlc7Z+VbpTIK1G0yowJSxifO3fq6
V/1aZi+o4AG1O4GyOYOTnjnE3T3DXXJtTKYOULFtzeH/NhCwnSI5AjeTd/JgL7V/HQ97yXrA4Eth
DcS93xlbhgtfucEDvA/aaKdP5auhQGr+8nDOVefuoqWocIrt2jMqK3pAPGzrwlI1TdF8BYPDNNk7
R7e7viqSGqo/NbayzNvlzjAgn8P0bdz1jiEQ7V3cjekJ/LKQ6c9jJYsFeacwyBs6oHo/V2wVFsu+
zaw9T/6A6ec7VxwZANmeHNHe3awkgJaAmNm4v4/GvMK6Q6QAxW0Gz+lSFm/kcSQuEmUTYgg6NWfs
t9arjqvlRby5grQaFFwnQB8SWAlx1g8C6PZ8vIGv9M3Ftuw4el0rBZ2BFenPTwCMxO9UnsxRnNA9
83C5erNyFzM18bxWoKZHebtnqGKUCOO0tkr6773K+HkePo1GqrHkxoa2/vGA9qtHcaCA4dZkt37r
s4Fvb7JS7TtBLd7w68nks2h/gVF29owbkoggugJcnpA9Ste6xvg+7zpuD79Bf5d+6bSlAuQo42yC
K/Y2Wg3jzYXlnGGVHae7OAK3AXPk+NY+pC76pZgwgKO84jKp3Z/6eNgBUyVDhCwrRkqsGdORzHjz
kogFerRS1EnJq+qqhOH3FybcTYUV+TnUHP9DcSWDZNiEVht0x7uQvdyq0EVK5lk4im6kKMC1XwDO
ZU4cVilStGq1YehIKkfqYQFSSCLUgtfOCMlRPANiiIEggZtcVuASho8JqyxqUfraGM5U5fjkeaT8
xneOib+lZhh/Y8Px36PVSjXBd5mR2Zj4vaRBfewY2gF9wI3sfxqlSlvLfMm3Tzr7cr2FB37V1Hui
G9DCSjak7yAINCy0GL7+MuhTXU5iCirpYUSSSyfXNxovBKZSW3DwJ0GFphhwyd8nm3ZPH8uXJgum
OJ9Lp2J0qBjVQGSJ4SizMu3aT5wIIfI3UVqKfzH4IrNa446v1fYn6OdqQWOCkCOo7MJdVonJ+CYl
w92PvT+X/JDr0Ku4J8ei14+f7TS5gzDtnONxcxQ2RS2h8ZZ+2iWAW6ICYPTOxSUQkrUYY6V1HEqf
MG4VeIGyd5CXP7u2+sKetRHj0BMY+DfNnNcj8sD8b/Lv4s5e/YuBLcQ/wh3z3fb3sv7I3O9u5bVK
r2qipo296AtD8ac1XY6jy6e5Egc1oY0rm2B06r+OCMCZblz7ssIqCu0S8ylJ/lSEDkqBwE/F+F3y
Ln4uBrZsgLgt3HdtOefPr6sFx38j50Zm6G5cxmnKWgmH3hVhYuLtvhX+iM7aUgVfZQe/AQfhshXK
OjIkVx7/T1Cu+4g0hghP0um0oFgTRcgvnO/P/Ta7vy9O+TCIZFSbdUchchYv5xOdk0G8DF2/XW1T
I39Oda4mHSfwGetPtK5TfHRi0/i7/6KyoNsoKkcShHrKZjT03jIhBpuVcxLK3F3l1yVNd8+trQiV
ftn9/uWs/MlhftR/zNIcB7W4AO9HDB6kpRlutt6HIOBfcJrnA8ayAHlitlYMHQRso2qWIluQ5FTD
2GixpYIRLxZ+F1jMePWVzgUa0eMydX/ifNI2QoeszZEV/h4a+N9c1PvtmPijh58DITcu02cvC7em
fj6zooe4MeMW1/8+yleQDcCFj8bVS+nEb8IDBDPegnulupKR2xr3huU7+vrn4GiOaRprf7+4aYue
vHmWFMARjfC03WaNuqPYtbGlWFt9Bhz4WsM1kPixeVgNIwu7GBwiWHN194PSXK8WMl8qqEYyzyL4
5GbN1DX/iRP6mwB+OKO3RTw2qDGWCq4/gkLRoFE8Uo4S+rpCUZQbTuK9sOcFxD3xoA04//reoLps
SdXkDG0629IyXnAwLdERz0p2tCSPBCvJliLrfI7zoLOWYgsZ28NNx6/9AVkEZVEXYmRIOUhZxzyv
Y+RFrMS1DfmrkV7eu6dvj7dAWtFM5q2wsCNBqvZILDE+cJq/ge9VRHcLcIlH9rjpL7p3z4Op7Uq+
dPgB+QN4birFTU9FlU2bf5URpLaG5ykL1DYKQfT/qMq0SaJRiIlTLcQUyY6WSJEu+SvOZt/i29C/
75pwyG0h4HTnhdgc/L+xuBCG0rI/0ZwUb8PSV67owbRNO1Hcu3Eff0DBWMxEV2QaiNpSBl4Txv5a
QVbr9J1seYqeoibbFFvYs+knrUEPh/ml0zY8bAiWOOfw8ED5dAFW5dUSw0+sy1uXO1ih3JWRCAaz
l2GOw8oR4ROjhju8XQ4Cgs+tHolNyWVYI0mZO60JzLYu1nMut7wIML28CPsj0TOlrByxz4+onxpu
t/Faz9l99BN2x2Didykb0+UDlpJ5FZiPYZ+fZQqJhtWDqJgWV1x1ULiIfCO4qTxoHfKC9uA00AdO
Kt7yvDCCkOIL34caCpV1hDF00ZPrMFsde1M90OCQnq2qBnhWZBAfDHvYPZR1Gw4sQxj9M4MYBIRh
SdSuQZkWDSYYyEwNLBbwbFnEkgd9ALJMpr/0hMfgyuzldXhSQF5kohy2kGkEh/TdgOR0K4ckzOPT
K9V+lxN9sfqEyK5O3kEB/TaQg5gj29AW/GORVlDWXdaHvHPc7iKP0wJqUqLos0iLPpp+mc4zNJS4
FBZJBrdZGFw+SUyp1M9uKOEuSqMiulhYhK7nvI2Jmj9XOVBiBT7L4V5ZQrF4j6rqg8c6w6fijRsu
ucsQGPDRk78L6zuC2O2/fiNf608PH9CsHIObkRGIzYCmOTvYKfR0nhTiB0mAOC/HqtEnZ25QQ+4O
ZAp9pUtcZwru3zKBriapp33B8URyDeGzdPKGnyqG3wBNqt0KPRbHSyWBlwDjFVFuyN8Bcuvywgdc
X6D0fb8SRwFidE8zHzH2Y1/6uIqvGBssOe5RSXg2zGb4rhjAsRsmYLXE29yT2nzZkjfPYCliWF6f
tlDfm/CjBIzkDGEeOwfsAYhySoJa0WWrdYy6ADjVmGtqgOntJdOdiZI5MKYOhRPdXGzvR8hRreJC
YpbesEC5Xngy34Yeum4spoLrTvbfW5wYCKeZenwRjz9oZBqvmWgdPCsf6POtHIRvjASI6qC+SBh9
I/Sw0hq+EdF4r8y+YwgySTQ/D2evUhZEh/cyJ4RXU00FgzB+81Ao/o2zo8TTr1Cq7HBo/COE1cCD
l/NeGPtpx5ZELPpKeIJEXiqI78mTznFtlvYvIco4rbUoMIAfKmpI2Ypu5lBtc0LAWJsF33lYjJXR
jzFCKS/MfCpo4YOhKrwLEX++sQn8YH2hISVDkuq75Y75ESqqu19eALhTCslJ4ocujFXZIW+iFZJK
+rhyxFlayxmt8kOPQ/CZzrsdSe9Woyf5bZeC0yE9DgMgx7k7yZPz4NORvJHkY3ZMnouiKTzprxHz
uQFXQ13pPH2t/IWtNiMEjxaphSBQsduhjKHQhZG8qMwDyEKBkiwPRtfRWZJK8Xt0/yfKyUBTzWs1
cFRclkEQs/eww95bmdshHLdtwJIzwsKFY9/Ttp4ae2EjHYSU4b3JATuU1VehkI9rP86D+ZyC3EFs
XWfGbO/6jVX1rxmbAFVE8VAaZWKe8ETCiOLbPf4bykBunk3xGtiopsHZr4qeKvlZBQ/502nffSxi
8iL+Lk/O0Ru5xOkmsvwE62ndBuxCa8Lxs9RaRjkuKtwyAkGy+PhdGsaK9zY76Sx1xpamxczJcyEs
7eDHQ4HX6zT7YjFjdX3oD/m7FJ27p40d0322rgYhLZj41CegqhCbw8xsKAgMH3WQOYabQ2Ud6UJa
06OWIfZSAY5uWrk9Hxx265p4HghR7LyiTIYF2vkpMcW/Oh9DCJEKcKE2JdkaWBWUc+4bb4XeqXNp
Qo7+CK1+3X7O1ggTNVIaB5ajl7oDXzjLvod2ZSO1m2XY1fkIw4w6aIdXtnNLeSTlYSL8W/u6oLwH
25ixpik9fX6Fqdnms2YmCj6QbitJQgOj53Y6kYTrxWveuIGHbld0sOFwNphPJBx0/2uVqQD7gJ0o
bkqngEmyXx7HJWgH0RLB5VKIkuRQv5ARod19XXCzMkZP1SZopm+HTLi5NAIENt/0BgFTvemo4ZWh
DyUsLO+B5Hw13H/FQpBJ8d6UOj6RN2AYQAmFzIYbqsFMGqADV4V5LUkcBZfUnGVG7xWH7Ja/o4Gn
FOkgSjDyiMXXr/Px9j0Gai77LSEJv20Apcwv70zj0cMizWrUMEhxBoyAeOkCnVPLoqc2bAmAoVYs
YsJbWfR5l5JlU9QGNRxUaHqz3XOrQ0kag9dmtI0pyT02jeAYvYEpCX0OC9a7bXcbl1QvyIBEsBuT
S/QQ/JFRM1sp613uFJqqFKx8TLMaQkeHT0oUCfXplRyk4aFFbg1/i2LUnLZtWHsBzUzEkW15UCVS
FYoFW7cxRDq46/J0BjEC75Fq6jd47zwgyJpGol8O7SY0SSGTLHu1S/ya+cI7/AtmKwHnU62g0KIC
VEfWcm+V8LSPtFKzPJL7qWY5RwXyLiinPufhj9RXnsn8CGQARC15p7oeQUVX4d+LKyWs5MsfLKUw
FD0BULTc7gcSItzSgbd1xzOTYQuPEssSZB7gfs+Ah5Modfg//c6Ja++TO0DLK7jZbqfAo7c36e6+
GSH424bhCh0uPif7/Wm3VQp9P/sXS/6FjgXa2rZz5Sm/czoSOQZ8Q9Cqd0w7dSuFEsoafQQLATFL
hlZMMccDOmH0yQ2UHka9GLFlNr0+AABJj3uKXhsrq9PfQxLtSm3RYnbaN6TXsN2zC27T0FtpOukh
d+DzkSaHgmlDdHrjpFSR0mc1Z2wW1Mh8QwYxsZSRAOZYOm3mZirarYXuDb48opigl6peQgsBs2Jm
bQWi/rpupo9nBtoPWOIESkCG14Y3We+XZ4TcEWKt+OUtZEU/0XcabuW9uEDNqMhMEuydn9iB7Jma
lygyWudyUTQyesCkj1BkGQdnOhzg2vECMevak+TtFJxDE9Y/YWSr3kR25W0MkOPoPhTch0OFfgOX
5uEGqdE+NDvRFRQ/LHTrrPBXFoveZ7zZjZVfapQFTKtdirQr1GKM7yc++qc07M3TUtDwQrsSijAo
26mQz0nL+TRk994KY9ZTibW5Fb5NnlUyJf8IOx3zZafD0pYIVEDf/JFXfJ7lE6c/rMAgwv5l6TsC
FMM6tKvx9lQCBPZ0q8DTd+M3siyrZCZZdqELWLSOLf1A+C60dbtT9vtH1APoy+QfSmLiN+FeienQ
Pe35YpWeLpcOWB/zoioe+b4V4ehqUNcAz45e96el3eaMNMbai9xK4SnmdAihFduGcwF96VmI585j
OK0HSNy2HAvHR5D9I5P0Dts5lNAnXIAUCVuYrz279JAJcKpadbGfqyfK34SRHczLiCehN9TvwaUv
s/Q1PyBZGcUHO5MZgsv9pwETaOc73V7PdZhhRjV2eDkv4e6p+NfH58500r32u20FRbP3P6KIA+NW
bk2pmVuBQbvMIK30uTnW5UwhAI/9wcj+WlqMu0RkKqeLeHQLrur7mfhpFnlTrxv3/Vtnc+6XV8zi
5G+mM+15UijJQRZOxBNn15KIQSagyEvccjSSVq2tOXBvLqjgvqQqp++DclTQY0HHH5wDA02upd+J
meWfIjwj9KPwrN745HeFhJpjCY4sJyN3hpnhhqNppzKkngtscuCo55kX6Aj9fG6yBhUjVUnPseoh
XOcwiGwkHX1Wu+FgSEVTSkMvT0M5dg9kbQf4nwXPMIGl//1corXPQ1mqVc2kOWDTWsrHJWaN03bm
T0KcK5y7oM0IvTO4xSC88iKf63QCcOEC2FYzKU0tIvrF1fLawViXbvIJnvnBQWbcgNQuH1ozqg3q
huW1WG79SYB5JmhCF1bar0gJzauzja2se4yVrzreEpr+iKST3R9PPNmpSeVZyrNH3DQXU/ZaNIrN
y7p4vOdXp8sE4uF5Kcla0xfvRe8aP21MHxfo8riyyE9bZEWlNajpw2hJGPkiZ+DOI33nIfRIqotm
xnC5JfEKTBHdYjsQDrWUiTht/9bZ4h2wUbGLjcLZ1FeirUBTmZeFiXemSd2GXiczuQl4Ky0/4q6T
zO+KVFdXI0civwdkurLYybJFzrizSWfBwPttr/qxUQQhVVsPKrkd/LKlkq1BTfpsuo46/aX5hYk3
SOBIZPO/3uGVkYempHX7J95Vs27LbuRo1+M7Bnd0dOwvFVw7s4i8uti06hZSbX2ZJs7i0HIRyMMJ
dzIioNymcH2FTlPieKwwefq1z4E8qTnGVIfXRxTFiVulbvnpE+r8FmwB7x5NlCcPCSPPGrKuLnyl
iLt7PTjanVno95aHKsMCCiIAx82/BrVud07FKaDmBdsTLqgCu9v2NZAJLaIrRO+n4Df4Zvy0GqB2
Br0lAVsshHelSgtXoahnYZ13fvybn608nM5XMAvVVx7dZG0dGiEGqun1icCiikAfoYkGYwaWwuNq
TEW0Y+UeaIhtIvvmsNPsHA54PdeJggO0RPTh33zz4cLaIe1bqnnlyfz8qRB/Fz7BEBaCAu2pTkTF
47CxjYl6JZFS5fKu/IVrrWOw1POPaDchNJbc63ameYjr7nDXXhyp84zYtXnP6zKUTRhKnrwEgF6c
xKU92AaUAyuDPdz7GEOm15T6r54OJQ+qsuTj8OxIviindfFFCJfiAWKFRIR3k4umfl1xLU1AMLDn
wiOjWBmDJ7+chTRoHXzsJ60T/MlYhoZV3ETPuftD5+xDDYkQfiPHIXO0Bc4aHfGCajAW07or1AmG
pJiufIOXJ3BH1KV1cBoYjQF5xr+GzzfGnJslhykZwDqo0kuqwyaI0a8CibT3egLsT2fPOaooJcaR
zUPA5Ms0GG8BUbe3zAlMETsHm1wtkz0eBrlo73SJseeh8gFfqVvU67ZZ2GaStChkHd6BSwujBEig
UMto52RcPNtS1gJQxu4cygthLyG1nPo2/VN3OPp8K6ZYGgVPLAlvy5lFc/HWVDJL09qLk+llw0eC
t+3jxqZ75lZhVPQWZODwF8e9mqej8rRMcrAi9Rf270EIQzkSfPOhFpf182716g8hYvGRxzlQjdTj
K/eF/reMUacOy4C9PK7e0bTW5782SkN72U7Q88yEBJA4JLMiOXnnQ9elz/4WlkAMO6zydRACGKGM
KUmjLDrKvNWRnVibGeGmadhsmYf/C1lVW0rD/auFOBoC2PH9PeswDoGgscpRQI3PvRssyPE8RinP
r+LSK4y+UQgPXdZ8TiX1yVXcUZssB+Vmpmwu4adtkvv5p+pmgHZGLOakpcTrg9peEYz3q5BeiONg
e5Ph/MVjjSgWOQd1Skp/WachJU2AJRapJbzPCTOsdGfwmrwH+FdUM8XCSo2cKmeR/+3RW/ETy4l3
b9lwvz90t0JvV9ZJjoOuKe2NJUx3c+u4eTkxhgS73NUBcc3/iYsQqC8ZUH2nIQ1JphoUTmRY2IPY
8oVLV73FDokeEqGT8TAhgGuXQCFOOz2CMznIl4i4T3B88GTBhfCPmGU6VXFyLd19pUhfxLsRTog7
RtOZTEUJF/enfLIxumG5iy8WJmYGAVkGBBnqaaJcitpaoN5CDKtz+Zo0GlqXsJSsP9KH2CSb0RFY
8HvsGeRpfrAkl6Ph9/ZPf15jumAzK6LDbhwyHwl83ShZ01UhO82FNcJmupV1zsS4YQ5XWCXaMWvp
lIVeZvfBza0sDJPYm3iOUl92B9M3aRK2OHB24N7vo6dXJWQpFjRuEtr5TIcL4UQJLyz907FVQq9D
oDMBe8tB8DOlWZTNj1b5tnq2VjZj6EqSRwYm+jGe5SU42lqlItp+7LtV4pFuhtQNycPv1K8xiBKj
C6fZl6c7Wpf9vwbXuatQRmU0lRGAYb8nITxRyTrM2YJFOUmvs/bftXUnVW1RopnFbp8gsANBIKEz
hPNlNgH81lKtb5phd5PgLmQOyuvLuROwJgbcs0WrGoJKcI2t5UnyO31Ew6uT1tzMt0S3RYJ9L8NL
uNpC6pUqDbDcamak77ZWcSnUMID7yKF/+lJDcded434kbJCCQrGIWStQvV5tPKEVurHm8lFnkqdE
hrgjldz/1xYTVuw/Rjlrr0+nkOnLgPtnhLbR9OD4Mc8y0SRMNwUDNsurEJJnPaNlnZUEkVlpcWwS
8tcALXvIYuGcQa3xNwhf2ppWcJ+Kos4hkNtBaNRddCjl9Hj+pljtzi7P49HAwvxAq9I56vQXEV6G
4OABVplEsWaVTiUA/lrTAo3zo8gC4oVmAtbbj+CMx3rxpFeYKjN3vwYWgAHwKi/+9cR0igLgSpKS
RNpB2adNwU3hSUwQ15dDpQblN5N0z8Zu0o+jo4JTkzG9tGnyjXVTkIT++wUgtiSYI3Qe9gSehm/H
WKrC8J9kE7e/cXTBA94ngonYUlnvV33TY87i28spMxPKi11dQQu50XZiA2CsqjrxXFOSdjhAgaGV
I4CBcO/txY6LhSwz7Ne8a1qhcSrdMkK6WS2miZezaW5edOEM3TfMxHtNwA3RUfv9YGtOKrHPEamU
LtsLXX412rvzvqKZ/sUMp5//4w0CQk0Wtcb3zYhNPtIGR7hFMgLVGia0J47cfW9BV5t188CU7SOe
d/w5MX2iPXxc2V/uKTqbG8i1Mj8Je2RaFjNVAeb8PvrGEEUTCX8+RIETiaMvM8V/7ETrzX4ru5r1
pWrY/+01WsWc+tdQXEsRBCN0tQrm1djRaxY8jq3EwdzoqsbVRrTIdvx3KBdVq0lva1NI2OGtxUNd
q2EmZSonhG96vYMEbGSW+HqEb2vpK8OD8sLr+oyg/hiobmwGGXDDfyw94QpCGFLmabPM0i4RIcZ0
tdiiIJ8KmaIBnYCVGKXs7wJ1NndTL0iZHFV4ENd11r6nmp+2G4IFRAZGlUE3Vu69lnQSZhlvdT+9
DqQlOCPYBYbd+CFJthWSqwv8T+vxu9X7xMFKA6cny2U1zd10Y+6fb6hYZCGU4Zxo7hH6FKNXuWdo
tfz2hT9UF2sjnuL8eleqZAZaQuDaOsuK/FgSg9/VphcLYrFd8wu5TKW9Ej5I6O3VGzUajejiodaK
n5TMcgXkYVxb0v+GIUKNJVgfamwOturbtSZhqmUKssRmtsDgwzOFa6sHUP8ONkeG7hJoeP9aKdIF
WNdKxC7AoSWBwf9LONNpPRqfqbonIjPtJutVmp3uQHs8fT9l/+gvFl+8HxeBYHuObwA+bBzbsN/3
2w5U9eZ54zKTqYi3jVhC0z1NdfSj1VJCZH6t8KIvT1iIv4mwJf5aDprp2YNUZ5OuylJufCUEhwDQ
NXEZCOSZMUx60tGs5Udb0K707cYBens0RfpnhJF8dN0LuuCpQ9Not594sYOUDhPyX/5wdeb7NIyO
VN2Hv+wKY89h8uM10HVmAmvjazhL/Q7NHc11pDCZ46k0cocybqtK4vXrlZrTxC7Cqy8I+3qLCPXJ
lLQz9HAtiEnm/3ojvuO/sUbtXoEH56SzNsV6V80d2LjnX0DySbu20MAuWfhBI2y7wyyzceBp6stJ
KxqXdQMOuCRdWaref/+3AW20qdJ+n7Xqs6JUFOxkj9Tfvz05BurTlS9JCfUsEyn71DUfA1HhrYa6
3vzgi7Xto4cXQfK8rmVytuK/4neHHDXauIx/1urccF4YPkCgHibpP64bxkHNbtkt2XtREWP68wOi
gR3zZjiXoBQP7ZoaGBjzljPWC1Ii8UDYV774ZIEqTFSCB44osr2ifVlGVkPNQRfJ2dFeQwa2Ppxw
iXrUjDSX1MEPljontgAO2ryGYWQK8FFZX887KposUIj4F8Tx65mNGtMaW4AlbGLDLsTkg141xsVe
Z1mNHvj6u7Ik6jCt3RHCA0eivzF+V+Hch8wsMzYUPGGX4eDeX+XRJv1XDStgO9DTjrUrSLFhLkIC
rojw3uBxx+tT/BPe/6Kxi+xzIgMYcrHUl8mDI03/7eFQ4Z5BAOI6gp6jh05XaiiLGi9Zs3zWAj0n
zKOnNVqDq8TblckUoVUGoPYb/ZvxBJT3oilx6z7r/6uBXQg0KzQpTUBTgXESUbm4BfGaMRE0Xmgm
uFXkO5EiY4+Y1TUsrwVgowXuI7MSZM+MNLsggCHvD0WaGrh3zgINDPhZ/TkWO/z5CDaDXblaET3M
v0bJZm2OfXS51/rE9Q4UB8dzkPKONtBhIuM16jGR3D2axuKPolYQPNKGwpuIIYWakMQ2X0pgdgBj
BKVuwky41p7jLsg2SsGqeYbazayfJnd/k2yV9VAqqK99Tt9H7xw34D7SKBb2DjNgyRCUMziElVEr
QwMh7Dk0Q8ebI1hRg2p9On1yrwvIwdGdXuCKAJinOCPtmPruAp68lBZTkO/yATN6MAYrDeOCwYw8
aqNh2PZWVTrdd1OVrHc2dF0O9uktgMgyF7hgUvc7iJtDsyNA3qqkzTfKEbXm3DyQ3SlWEiffzvBe
fhUkHD+cydWqc08MaekWfF0cwSM8pJjbK3R7XQjyFEfYVumerMm+kgeSPhlvMk2ejCaFUOdV4cvV
KYHpyykRNZ582mmYng0OPpukr9bcMtWMkbpF3Vrk8oN1DYR07UkjmdC5lHzEbatrNmM2ISLpR5No
DjHanBdIXpl0z4JriVfMJv2K8UujbmvJaN0sB3FGKt/21/ioOLsYcuA9kw19OPfPqMEoP6b/cFVE
/TpTPeUsDDNbZsqm5ES5TZMPGuR+lXd6RFdetcn3DyGp/aXk/ydPyTow9dKOuCkdhcTFkvJfq0c0
xAuflE3QXF716G8oS+HOK5p/WZ+Tegu7cFl8ahCXkT+t1SbMqMSSvLpvthF53MFB/sOxi6NdjI7T
ckxN8ulP3P2bncSRrSzmbcQH/6FMeYQoOixQzwEky5yxhxXU9O3FF4MNj0yNpeqrsy85adbIAd5Q
rnwa9xoZWqw54Np99s8Wr3QeIfhmhGtGT7fA9333XtJYeOKXcziL7ZrNJEleQgiVWWhsYGoWpZ1o
O6FQUvf3QY2UhjKHdOd1Pg5g5LO4pO1ApBx7itqpp20tqaRBTcg7j97Me0Wnco5H9YWsX9KXHFdn
d/0Rg9YYMIxspbxlP99CrxW1LS4IpYsyiLFofi6DyFPFloxzaZCyEUZhLddFFM88Md5DBFMVDBaa
7ef2iLPYI/7SAVqI6Ylhivmz7jdWDKAdeWgWGGqDTQvxcL2/Sw/h6vGZNL5Zo0bkkeYTK/Xbh7Pl
6QI/HDI2sr8FVempuz1cmOE8eNRuyT+/CDIhJKMOh/D+o93ghlAnNPWr9XozkDh3SN7oSkoGDRrN
E5QBSmwu/dcpmzJ0BChx1Mfy2IG3CwC3aM2XSNG/14BKFkKvmRgsilgYjjsqZt1zOF7fhtBXQCIK
E6bI47vnQ8aviuCUGbkMu1Xjyqs5MUxSXnX5Jeezp3MsTfF8nYI504Ja0X665BZakFV9Hnpkq2uj
qZadP2XlcNL+hYTsYBLtXnIDF5eHP2AjlCMDHrjK8uKlu8iKZUMfQ849TforxZFq6mVyIs8rdQgM
n4pWsdzmSJaTvUmab5zHTTZSFPrlW7bHk/yxtiiLIE5EOu6EFgI+8fTFCug49w+GGDsLMZv6Bb6v
8J4S3OuTnsDAT3H6RPPNgnZ6l/CrQfmmoOaR0tUXqyEPOkZWIu4jWOR6+5AlQSI/NhQ6Jl5oZ0Xw
u1RZnmw+chq8ZNctxvjiQybS+dnyCJw4HKLUgrBTuIjMVyGyurPZuL5TyBaZW4eY9gSsEmaMj3+v
QDyUYSo2ZfohoYUzeBvIV2chpr8GNhFq5actj4z7poxEf+bnviRQNeofUvKQRfkn6eSDkh5teYWL
aaZUyFYm3QDTocxC2F91InwLvMZ6iwxWnlNZpEw+Pd3QCjQEeeUEmJXCIb10oCVwu9szvrf2leH6
D9lWBlxH3PUdw9RL7Gp1XEIKlekXndlzPSWiYaE2nE/Jx9+ZW/Atq253t2WBD43QW56YKzqtGwvt
5k6g+2LN6b+DDehoH+D14I5ksDALywwHFsA2d+aJe70uB+VRB4SJQbFTemc9WPO8RFrqfQLRmRQa
6aM9A0Uy1/p9qa4nsn2n5A/YFzJAqGs84HTYFsK5ofhZ2ByijiPJ7KKwJkcVTbtWPGfW/TexYFEk
3D0I4NNW0abZB3Mc2UsH3TMeIcBN/3Jx2C04Hxl2Bbwd4ACss4qABHpGbne3USb3+4l0/t+SQ+Iz
f9gFRBYCUI447TMI5oZLsk31F59aqP+RCQ7M4KFYssrPu2RioSOr+dokrR6C/aikeDjqTS5meheO
mSsEhq3TAjhTsiewBzFPcl5dHk8BNid66J+bMELRrYLUeq8pfs0LmOULSPNXhscCuo9uePnyhSu8
VE0D4Al84wNEUeB2/k0PclD6ZtZRnwI7wzf5D9MC3FWR0OUtqHFZ6KeS/O2BAiTL3QbXJ9RwniLa
PnJDDPNdSjMKKwX0pjnZejg/O3peDQ50Eg1OjwPWqwCxALV1PkRsiMP2qlCSaOVKbmk/Ule+NqIb
q9U1n1wuX/Im2gLO85oTq1lkdBfB3z/QGdpaCFVaS/0K1pQnMHkz7LSgOEmYCpPcp/0Y+LQvuxAL
vsmfkqKq0KA8owU161RFfKUBlOIhGeIpwaNPfY4vMHfKqOvCjZI+AEQugiJeTlc6evgydNVR8I7p
4/6umC/AcAJy9KLfY4M08HwIE4vHnCdc4yCXlTxRnpK0M84R8afAXzK8jc+VkaF/70xOo/zNhfoW
XBgB5ge5ucJpD9f3Ea17Usd6f4s0ebX1FVqVbakpyrxdmyVMgbnpyCEE02e+T+d/ScinC3Sv2IPZ
MAhW4UCVlBHMoZpwiXkbBcU5wjYPI+OGeSYRWSksY0kYLvDqZyAEdcCwvoZPYuieLS2CcOmZpxZm
WGEKu5Zhrn79F9IMDEDVXcyjnsmdL748fGsZm9/t9AsvgZfrJmnPtS23KbamHOacx1mPoe0ZDi61
xC7dFp5Vt+nBreGVsOgoLpSThy5tVvsKKKFzjf6yZ2nXqVQNuyJ/DlWauftrl5+GMyQBQe+6h/7z
zOpiQj9mKDfmy6mag498czew/up1uKo/zA18bfOA/E4jITRdotJX8JXyfpX/1nOs9OIs3D+X4vOF
7FXMo7zu0GEcK4vgZyftA4tDu3WkIMyQwGEicIAXgnghJS9zNNqoaAHMAbSnkCFzWHoMbiQ9rAFM
bzV/o/NB5aocejiYX/lgNFAq8JdG6GKzHnWvIcFsMb4wyY08B5m7tqpFIu++E6TsYUiKXWgbm2QD
bUvnG+dD8zuysSntF7IkgVEQpYXK0r+KvHNhHrTFwGy602D98ngvjCNWocglq5Su9WPhd6/+5wIe
QydOZ4kWyojJhowzQkKvYQ9jQxqXFz4kZNpRWBUtF+b/umbOe4oAgKXNB6FzJpr+W0Z5vuy2wcG0
JqCCPwvMhhUMOZt77XXXeKjO6XXdXsGeNY6o8cujytr9JU1a2yJRFVc5i3VTVK1mtxDehnamTtSU
2HVFf6WbEjB9YCLLXbvY2J8HZ+i3S17iVXTg8cl4VP8p1VOVVsqi5/rnzTkEGyCQiFFrMDPlm56D
WtOMyVQs4+nDvS8XwZSHuzoP58Rmc9Itjc+R8LgDXDr/e1CDxox+MtmjTOt2PritoU0K+lKwnCIq
Vtu0EoHQH1XUPI54f4jUJsPwS0a9/xpnoAm2YYxrO6OKlTEA+/KhyGNimPlkKBjGt+Z3w8Kz2rFV
ukQaz9QgwYCVKUjnw6LCmFsGhG4t3V7vOEKA0IIvZw2Ok5h3YzNJ5e37HZZU1sZGhaxDU6ezBdZ/
emnR/XYB4oF9WUDAb+k2Z86Sf12h8Te/bcRQHZH8zxM/AwbByZRNo63I/TjheSA59ofU/ReGTAEQ
Q+mYNalJ8fEC4+nGKdrjjIcDlzIeGJ/5/nFn8GGrgWUmPmM7BaHR7h0M4dQmdI4TMKlqF63e6aBX
fJfNHXjGlDSm3HEHG0r4VjH6JEmIEARACO/1kfIU1YddtQYgScREXcSKMQkvmH+AWLvWf5YQ702T
CY1aIjRvl0zMkBIuwS8FXbKDvR74itIJqQL2MyUC1mj6+U5l1O2nb9vFMti7fm9nB8bing9cw7aE
HvOQkGD1kWFzxCD2G2RGkLofL2u65Q/zB2/iGC4vQH3otRb/FibFeCg0xU6zbyZ8eLxRKNTRhR+e
cFLZmtChwnsg6Xqk1+vnRn47MXYEV4cabzX1VLULn1qwgRo78NAmIo0f586QW5t1Wfozu9G2MAUh
/ssIQXR79kGaIqyUHnneLfX2EM9QdbwfvZ/KRWxsZGR3dsvgxtIO/yMmCSx+NNPEYf9FhB6oP4Xx
tdCJbnm+M8A6A2ZDIjYcJVkhQE+/Ha7klopvSlki8WX26L7B2tVqWbXByDKAKIEIbW9msllmVchF
O+P38bQSWTg04MxW/6D6MxfJ/kRCo6YDRC1WKoa469Z0JNvPvw7bNNaTojhLIeAdfWJnZHyppvZo
swGIKtHMrtTXc9XajbrMA6IwfNvG+cRpBaee6SG8848ApEOIGr9gPjIGsfa3n2xAy/u2fmDRGYvS
xT3s9pA2AGlTv8IU9RNBxPEXMUMQoqO1xhN838dYQ4zJ5PtSCzq3StIh/GOxws+kt6neRJXWHDA/
mTkgHZ/rwzpNOGYEv8EgYmPWmh7Mu/cMdG5pZcVh8/I5xltrHtVST2/Y5bCuwS+Cs8R+qOMzJNRs
oeRmLvvnPaI+QtRF8rygOwCyc3sv2XsLnTnTHYM4+EQe3SZjCJdsgame48wiKiCi81B52sc3I14u
DRGCHqpUFpF6/qFaxeg+nNNFabJKqgAWEHaRSPw/6tczh1+6R6zkykJbcQBqS4aEP1WjNBNLREfs
ilYM7QvTE1Ud1MzZy8BFKa84Urs73nvz9W5oU5crlnQmTTFdzb+/Vxrgr0EXItyyolt+32oYKpnp
qUPXtLTGaiYgopn+TSeLoWsS05t+tyUgBjFxVYDS8e420B0WcxJYqrabqwEUCA05BQDiWPUs8+q3
GZ86/D5aISOsdRIzDJmE6w2kdB1ucYAccwUWXKwjU6Pu7fC/3fMt94VHmv1IClE3H00D8dhBc3gB
TzTpSF03siRWzMrluv2KOWfCe/kkfs4Q9poIu7Tcg/qde3dS0hknt6oDeid8EenKQ0BE6+iLz941
oaJYhBEzkW/B1qjvZCIRYJ+lcHPN87oGT+0tVx9ZKMivoxsytF/6IEUL4oujvvs+t5OOO8dv8AgR
kSBa+OkCGOoGnKKdZrIQ+qeFAVenoC7cOLiUqnezguzeHzsOy8UNTdl8GQ1HhCn+4kvWNQ1K5Wqs
aArYRJ/KneZ8o7YVqft1gHt9wKyvwNWRGce57FD5P7+xDkhH3sQWEN4HLKh7yo9L0nt28Oq4B4bX
XtoeoSyUdStDBAnogaU7zneXJictHp+R9q0zHOtSSKwAnEmXnPf/o2tLpQkriZoXAYVC2gg4PEOE
Y9MqKO0cs9XlfjVS/i4ocmEEb6fj+IY8j9Tjo4YZiho3A4PaOrPFMM7zniDMIKTpFiPXa2/KgHBf
UtOqUxIfprZ1XLE6j5cI5XCwXYTRyflifeVGFJifHlfe9DZDmLwE8GaEEJLV9QtiVVINgiZ6wl1Z
yrdPWhXekMBynu8lyLlzWGIUOBCb0cBGB38krAxxdRbKzHcX+/AGlRf8eOnFhYhniQUdYcPrqpGR
aPjc7dykgnEv7Mu5+E85RuwFNAc2sm3vR/7esaWrSf3Ui5TMsiYk5fgvdhO2x/edP5cW5yuKV203
LQE2fvZ1Y1Xz8jJCm5v+HabG1OoVqW+0ZKfdeIX0R3R+1eqtwfh4hJm+73LT5l6OYzzoe19QVDPO
amuVsTUvvO9SeStDNQhSlr8JWDszIcDt0O4p3SDi6vUHM9klwuvRXbUrW2OTFF0h2YlK00zJl0lW
NqkBfSB3afC6BqeHEbnJ6FrzBeOskJRxeX/WJaMwUQ1j/z4TgKDqqUHtdXgvO8LjecJTvAmbT0jB
m7UYCmPEq+LK4szT+8nGrwJB0N7FH6Tq2n2bs7UYub7AhPpxozV6uQJXCZknE1ovqJyTd7YVIGuw
xiDukoLIya9f5pqmA86bPdFkP2UXHju16DI6ilCFNurNQ40LKmdXjuiNnjXfYsc8tK5Nvzaxa5a1
3MXHlCFHu2udbVwCkvcytX7RrVbVSxXtqtRbXUqKtNPAsuflzHGyzv7EDGPLaUSjJllePmDuqIZp
b4rBN2emu1jYZWxyH7aAlJxeVtB0TNzz7hIGZDwQQY8RtZ6DFWkdalg2TU38VMMPVqH+OT31YfQs
ert3TVEknh0bFmTopXSU+hz8SSXMuAwmvGij2R5MUdCEwpFvarlC03TU0C8O+9wkQinqNsf+vdSQ
jEVH77ubi9sP0Yml0cLsa0ygt8+3GZnGPf3+xenqPoSw88A65/Zy+m/k5Zp1lHuqXT9tVLu8Ggy7
bN1kHl7hlAcPDsd9bMOvX8crI14tXizGgxs5Nnu7Z2LGFph5ll8yl9aNwIYHZgirS01Jv98iVd/C
eYLR9fA7yGr31bGlgMCMFZQCS4YEY3NLIuFI46tFbgOamZcJdUPmq7DR998IaOP9D5FeIDpiS8WL
4NXsl8RisFFIIbWnFJUqseUc9mr4pUbK0fmvFjQdaHH9YeMmyOtWB+Wib9dXEcI6sKOlqCSy468K
2bquwqxJuqowJh3R98KV8pHBfePC9Q0lcsVU1tt0k82RbgqClloz8D5m8n7lRHTY1NnAxQlyuL+H
k59LIy2MsihxC+aiw54H9V5ufnVtTiclDM5zLLUDMFoTRyLQ5lo7RUvBIzJwksOQIWPlJ2C+RvtU
QJOeZ9a670FoknLTuTRCYJ/uV156JZMOBrzJxkwvZmj4sID7W8zb5Z+fkKNG6dOrO5tJuWY8tSSp
ER9dnP4gOrBjKfXOk/h1DvyUuk1hMYD9lsfoEwffGQk+CfaAbtVLUA1uacbvKWm0hHiqBY0l7WD9
uGzxMnpw0s2ufXQYwEDa59KyoxQAd9Ww+imyYPpGTYypPdKGEp1MmU3uNzK+aQ8xs6nijHywhfSo
l0273j03IIwf2wqvPERxc1Cpzn2C1LrIjCIOsRq1RkhOYMc/2biL0Wuq5xz6Qz64iJypNPB48q2j
992I7LJ/1+EtXfqe86JzTPIZFADecNxbInFVwzzRQlXPUpeIjknFyrRZK3ZYavwZh1jyzfOaw3SL
STa64SUb/JknmtOsn1YM1+RqAKlxqVbuf7kk8krgfJdkRnkwyHo38UzuBFmnF/rX7K+7l0Ckq9VE
dG2zmmer/9Sh5PeHVUhpPAzEZ4ZChhyXd0Xc7+HZx2861BaOFY3dfPUHaqGlgnO+gAmjp2GKqQyr
hNbi/7nKIzFdrltZhvJicugBkGe+hp+Ycmh2pxz3O8X4Y4KyB0dc09AjUMNZ0W5tzZ/a+lzaon/w
HZ8yf/9nbaVHKY2HbTkWaBo692vRd1DyhFK7HxzSNx1K2qg2flAsIYSv6haheP8QYfxf1Nn2Ov8f
wS+OKYkbtlVbYq6s0jTyKD5QwcrFJ6ojKF2n3oPcpd0/F/C5oChzrbcGASXwyybVCAcmp5szQS9H
gd5ZCsWNMJG+1LgKaoe01Ij2t4YOqINVThwjRnxgFTFVtX4/danZR+MZxW4s1NQ5ZyLRF9m/lM7T
U6SuqPpqyMEiOVewzvqL6idYv8f93YEo/CQ+Vgy88rz3peVubRHF6pbIRCsJOzm+wCKQk9jAR2qu
lqDguVqMFrWXFmpxkBbRN1bGzFfuRPLMRxekFDZIGtEDYWYx5DgUGiEzGNaas//KWpakubtV6PCu
Ez89+V6OuQpsNLIKqBRkoVIKuGaYnW5tk2sCIws/wQLyKc1fn9wOtcg6YjDc2PwI62cWU3E2uuzH
afyi5bLov+AxAbzw4fNJrLyHJB05SPSuDFkG4MwmMtLIK85wzJaMt5Lf8inqLAzwo4DS5DSixiAz
jpGqT+wGOunRWhjHXv/q9FVijp+Fg6PpmhKgb4uHq0YPiDHQqA6Slz74TynNL+Pnx2tbsG0k0Z/M
XuHfsQl1Yd86u8qE4XSDa2bbG8JO4lbv/fr4yuiNUBAk+lqPuFgCth8v55fZqOpgaSJonfuXH4Ff
StqfMfvll6s/cSCUZ4ItTbos+0VFU6dLkNMeRzu6EKvywcML7vgyvWQB6BvZDp6iNzdg0yBi8MyD
mgauTase0UGWWzEJG0Cz/fLV8Nxa+cBpA6mSd6qyDMsVYAodKU00xX5/5E+ym5N035R/6UecX3wd
EaPi3ueNZOi7Irs26MDtJ83aEBEjQIeL4z3X6y3NSsiBbUlaAhi25nsMC1RaNfH/PRNWnv7CA0Hv
9kjFj0TE1+S/WgaDcfBC68nrXFKc/4/qcLkJKl0M1JhUdRIhRMjTs/cGuAvIgr2p1JGsIcP0M2fN
twtesDBD6Qpfr6Tm6PXkmAbHRrri2JpNEmRSJNe4gaIqsQxSg4MEUvE7sjm6Spi+/GtsECw45/jm
cT5JSQ7PpM8pMVeZt1V+FuQH2NXgx1eJqIPr7G8mNNrnuuqsPbmFvFEIgsYNFluBTN4+ZBCQcxvN
sCq19129B9iP9KiqGw+hh7+6v6BQSa4YLgqBiHJ5VQLFcQ6UQumpouSb1l5Ex0oXZmcbg7FAGGTC
cudM3Ej9VyBA2dxPZeVTAAZ60BAS9p9ne6ECScGm+wp/KDF1OU/g5noWcojeh/arwgin3LiH/+dZ
nP98XG3xM1F/QlMbBpZ8DH9Rl4ZUQSIR9ZLiCUbicRYR0SADjzv1QBH74OY55q31WKL9YlirCBSE
tS7kbzT+Ij0VXZFOL4uf7rZEC/gUrgtBHt4+bVSPzajoKfViwaOFxeQE4xhYoyEyX+bBHUmquJ3l
Xn7mUqtaBvgbxE8CwJqPnoXFLmJwXZTNHlU6kp0RIfZmYbJhMePM+Q4ZtwcGxVpVI2dygaf5EYvJ
IWKMhYqNvIfiMfBf+nEttjBXkrC8sdj2uBKV1CMXKCPe8HLHrGkpn9igZbSiVJMRjuM7j4/ZAR2d
jmp+1JFg/+N5mEOsS9OrlxC+yLSOaRN1Uir70AiCmPxhM69mXorSrOx4QNBaoKf1+IiNCEi/U5r8
ryQeM3eEt/NnnCqChnVe6hqu0OBOebvZ2OBQuSGBSLK8RwgHXUZQUp17gEVkIKupa1rMNk+G+8RZ
M+IECSRof9ioPnNiPsr5YsdrGmCR5EKiTGxbWFdT4b0koMzOxHFn6IHmV92TpujzQBUufokMgSn4
ZJ0QuG5Y1Ke3SL974o3kM5NNo1ycWTbn2sUGWOr2/A0Dq6HYD3+U1dkbUxwiVTcBv9hflHTDeGZv
STu1uJbOiTXB0JKeUgMFxbkwYcqAwnZXK3+9NtdWc2XZGu0kQ3nQk6j7LtrwVltnLaB5XyYVcomY
gXBYo18hg8mA0RJhT5QD9/qcpfrMccP7By9rC5XlqEQFah8eoatPoOlvcfi9dyFbActyFlkKLv4O
jb1nf+4vc1huiLO3lFdyETUR4jnMLozFiz2hUONlV04u0pM2j7l4tc7CHCswAArdZExVNpO6YDPP
kame7Y6LzQwB2qWoDp42pJlF3vVwq36E/F32Y4Th/LSTn0TCWKJm8vGBfnxoSFrbQdQ3soNd0eAb
JyGSfQZAGEFjI9P2eazZP52bNfmhLmcf1va6zVsdoqfOnsDPbzPXrfhAQ60vT5Wn002A2DOVZopD
zzcrBdKm7Lq3Ys2iU4ugZLu1ugNfykEnV/pT4g2bUDp5zvIE94mmjSp3ceeGx+x4ofG2iPHkgyWo
bc8HhZLSjislIoMtPma9CqH+/y2xYk+h+KYAQWX8V1uxI8QUB4UHa8Ldz8BGL15lxBtArO5trIDu
Eb8B3aZY+dNA4MrI2Hi/m0cJUoJ2KrHeev7BD08Nx74ItGGySokB4Nccq/wfTpKZdSIRfAc/ata3
UL7MtyDRtGnDvPnDqSgQjXAMpEDv+zwudVUpiLjP4sfV8X8Xk7+oBHmCxwytF7WOuYXWwdVf2VsJ
TMStKUx8Fkvc8l6pATBbavj9pXWEiy0TTpFD0juhzuhFB8muz02s/+2syrHtpB5iTep/UMlI8gaG
vMVpoltTtsz2MK8DG0MNjUbo41HgEXjZfXw/X4Y89ZDAy2RkwkkPXIc9aspe2hzQNI0Dadx2IMhm
lpo5QZ329wAOCFLne4TVp1qnef+WYUME/jBy8yrgVL4UcxGFLBo+yyHZ65dha92LsyRLekXPXV/R
gTJedZD5h5keldlsSmsnv02oqGWXjFbu6k8rej0ZJUJDu3H012Myf0ibEeWVK/9N5m8r2xVejiGC
NmxxsOZ+N8VEgBr4IOKI4TKmSd8rBSZWAG9dP/S4GbqJSXskBrEE0R9fVBos2/nJr04SkxNpIA5z
5FotGGX2WIHQjfucEYO2N/Uyo1N9pv0prC/dAypzexkjMDr+BLHgd/CW18enrBHaHS2B1oAmwGKJ
zGnMk6TL5+9Kx1Y8cTWGOS2k1YR4lUfeehsBxyt0KgqzsDAXivni/be0qoQ6HTRKRwL9WUTYJD0m
Q4WX1CZrHUITLEUBtzpMXp5n5LjaXMVa6jV8PX890f7q3aZYF9peH8elilFKjlXLnp4ffuGmSAjJ
iIYYoEvYT3WBwgxgiuRuGUG2hrHJI/+P+wvnQxmkaffkhMhJMaFrANoLwCU0nyV/0zvyqJfR6fMO
7KCxfXpS4D+k9+4xn6jREjkRl73YlNS/2T/a068fdJ9txBMeQTl5TPHXK9k1O6nd1cwVE59Bd8cU
LdoAKeZYhGIhKrM2e1GQpEK6MkyZsThxtn0YQvhDZrssnd7nHAuB6WD9gJ7zcU8+BZKVWgU2lW2H
NuqzxLVELVCPuFvZEi9kJDysqaBE36vnr/ePMSOuflJVHBS3ApOifeMHUHy6pXrqyDQnMkCP1GJR
EJulWtv0ZL3DfIB5xp9zWOLVLqENRwRLiZukSu4H6U8Be8bZpkMH0wFohxkJ8o+l1P1BbU/WvUWv
UMMebtzlARBuaYKkqP6lcze6uFGfFCXUnFdMxtFPJ9BEBlMbrwTBk2SufdD524wJanwMDtT7mpXS
nEuVAdhKTBadp30kPZbiD3eeBG/Nbtfm+TdNXbuN1RIqGmwZHsdJTJwHIkWqxI0KRMXxIW0LH7jV
pSWN9DJea7DH6umspCQdB5MdTaaxDXZ8gxrMKZzeUfLqLnyWJcJz110bEAm+GCj5CCTYyfhaVb0S
bBqCbM4zqTVocXxp2/n2mhr5N3NkePQ9d3h0I3ewhsL0XMwf3dDE+sQ8Px18myagh8lVwBR0075y
+qXj+uvc6iy7WGbKtGEuuZScDTojjwJOyZeCpM3wtltec6k3g7xEVeOBLVgqmNTGOh5Kjl9HuwD/
IvBYxeYY4jEszEJB1nP34YLZDtWMsfc5iQjDUCXogqbJ3M4fwhIAIlwkRlcaunRUNQmsrFtx7720
CtLPnt17xQvbPEaijtcV5RxyvDT7aRF5XvIa1t36lfYhhJf7sNV5WIVealLN9KUfwyBeTEA85v7V
PzI9hj4sMQB5yxNl5y1Z08w5W3lNNCov5s33DAzZCwBq0ilEqixfW+vIR1FsH2DsOZojmCMajnwo
cmGxNmxYSSwTANSGdOUNUmoryinb40EekWVCUxI9aKAaoS4C3WaoD5U62OT7qtT1Q54loT8r8CNY
vpKLpzcNTR7ZV/EBO3qBCzpUDlUCiO2S7B1sqg4vLohtK459Vb4Fq5xKxHELBEbY7t6xjEunipmL
k0S3z2t24fH2LU/gqcXm+RK8Xyo38xxq97ffzrdC05n3EovL5hg7xRKs7rp8y19RXUSteRb6gNAu
cINfP+ivpYrFcTm6BI5EHvB31I2gax569c8FClZYrGNhXP8NVq+rXX+RSUWshwY1VMhsZbLfXxJ0
NLQpmb3uZHNyBaAZRbvH950vn3vDZ/FhfUnVRkq1cg7niScDYTDmiUwr73I6gVLC2W6ma1wIfk5P
9HZGmvjQvsEUlfOUXixsHR2vG5tslfQHq6Lt7YqhKHR8VYN0zgNB0LCggeNvcXGkKEWlJu2eCwkG
1c3g2Y64z1ZZFaUCnjShHTAq0Bz8sp2beXdmS2cAk6T9Wgwo7mrY1RgDpD3OZ+RwwQE+rFgT7NiF
92YDn6mQfBLeD5g9CWN1vTNYZjKmoXClxFaUolX7LRXtexTK/39ARv/DFiC+JlZ3h9uyihFNGU4R
rZAKyQeWkuOvRyiOsxVnqsESoUE2D4NAMPg+Cp+thviUhoxJD0wAr7rTddSkRZwLdVKsYlOUvAz0
F/4R+W0nYXiwCDXBc112tDyDahvwmO+lQeDl06Zm+r7Ir5rdMdeETQSOoyw9CFUEZnkYJQWfJhcC
lSbMwz76F2iGFbdHqqNggFJQTBN5BiYAFAB92TZVe8e13JUubxHgQ2P2fYczn4+YsDcAJW+CFduC
gYbo75mlv+IXCvxy5n9b7FgTlLSv6erN1zkVAtG865KqzZU43mIL3Q90Woh+Ak8n+qCKFVXoW0u2
JBSUyGFVJnNj/Jb4wSgTvnSQjlk2qY+5GRM7zO3icuH0tWFUq4Z0Lg9yoWIaNs5LD/cMNy74tQHP
o2XOv5QrKcjnP+wxyAItbXdhO8xEWiV7GFoot7Ud4vcAXNFk4u+U4Lnz+w7PhF/Ft7zZx3PCiAP2
9KpgaC310Hp7WVvSdOfpTJ/5mmGaDLh6BTDa0qdNcy52Cbpscg8brv+PmH8sG7NrI0gdhgfvP9bV
McOe7GL9TkSskT8BC48+Eb8kbR5WGAp7Jx13qCHCvPpmal3T/rNV811ZGAZjNKvju90w8fHw+T2X
3vDml4PVuCi9PhhB6VjSdPOOB4SaenJo3lbtHHz3C7eF4nBgDeedhE+S2jPfs32XrR6YimSVC3gi
KKo31/ZfInFVFG63ZlZnaovhg9bMixaYHWLGDEdkE0yHxHlRaOZFLaQhfeaJP0hrDh1XFQhNI096
9/gxbe16VqfMGcUvNWVD4bhDcwrldT34KdyWTvBTJnUsL6GUON6shRFrdsva/bw4Of7Slh/3oPs9
7ys6wR/Ehhnib2sucGAkjo3rYNpJkSdB1TamcxLJIsD3Xz+dvptgVtudDDHqV/BZF2Nx9bZnySA/
9Hn1tGdoi3BnsX+kqIZP5rbXhMKzS+7/KMawiP9S21BCd7W/yMrCgr1VRgGcAi2dc7zqLsGXOamS
OYejdd2h0eJADTt0WpMseUgegqoeRqamjTYYPclb56KOizXJjAVZrxbY43F3i8zTb9twxadPI01f
CN1Ah8dZkaowFXLSYRTXqeEZY90dPu3iTV9/SNpeUMqI79aG9rALt9RSPwTM7xiZSIKvZZNbTHa0
ehJiEWsbQL7zF2LVC+YAmO8VeZcadiE8DIdg9rT9ZRxgfLbPHGztuFzJvUBZhC/bYuurmgjmldgb
J94rIm7e2qD2uwD1nVeIKhsevpsU6M5SAU7dZH+dHLd9q3dTgNTFp7hCtkabDdnIwyrXK7/ga7qW
Hks68FSKU/+nx8+fz2v1mFZ/lvWr2AHuypJH3Yi/gJikbjFUcdFeNsMrCogwIwQRcyEUQTA5I8k0
ZqfYnTtX7yz+omipNsARJyGQ3jLZVk9I5SKUH+rtGMsMiOmRFBBdj3ntRLuwjeuD6s+Y9EVTjQN0
K5j8fiU5FzSWn8/E47KmfBkKeJ5DkUKE/S2JfSG2iaHAM0IXDMTurraZRM2NRhUJdUsmReRo7h0k
YKeavYqWkYEVuiShsI7QVfVoDbJMcdxxQurOWLHAW5kNXD3PaTtQmYSLZHXkCYMk0I7LRn42LP6T
w/OG77HQSFzL//NJo+BxsuiO5AjcdWDZ8Jd19NtMn6XDe1X8NZ9QAgIq8nhkF5E9yA9v2WhjRtxb
XUMAoxZBekLhKY8dPutNYdH7IKgJuWWvkCnshmEp7dG0M1Vv4SxSo1pmr+4I4rbn5dGZ+3xux93E
1eP8dT0OG8fy8zNn52KywSTiUTB0Bnt3j6wmghxN4weGnRpi+rZQJ0O0FitN5/yuZuJFc4b9jhp0
19+Cv/jp4NVY2c32Sy0Xkq+gGc1FWDAZvC3hkNDTpgGKrBUDNOrL/6eoAV+pvvZjjJlgvOM/FJ6z
HzmelKmiWtWz56yVSqH/VqJLr0v3KrtgAH96umgaWhdJ1B4aowp2LE8jXf0ojQfBmI/HcJYfLCNQ
lRQarCp3NSJPHAGMBoXDchnxUMNzP97I++23GlFiuWD/q88hEIgxr1Dm7YWY3kIgggsFJDs4cxRI
LbTFFXF+d6hhNMDZ86KMErTWd2VhOuKCtBfMa3P1to5i6qgBSkcWJs5Ze/QbtSiGFsr1bUwXr6X8
lEUay8AdkBYg+p1wAUwl27pP9pVevXUogQ4GK9FP3bVmw+RmC6YvwfFv+zZUOwImpMChwBgn8TLY
XkgEafPnfdlsxg1q5QqunRm7xwQ5MhJF5PLYw1yvZLubIwuUZPrUC3RB01NDcwW27SDxGhmVbViL
9ZL2P5ViGeNdJ8i3Y0nLtLzqy9FiSaEgF5lqX/K3GJ0qOC8dfpy1vfaKmGa1iC7LuV63b+xdH1+A
k86ghYFX9OVI/kMOYnzoR/SE/fJi5n1R3dzBjvFbJ8nd30yJ4sO+PNYXXUMbVNWI0AEHsYQaEoNV
3iShyZZESuoOQR/lpPLL8pNSGmYeQ0aNtw7WIuAOkBtt6QbB4KHuarF+Ab86HkpxCzwV56siLQJm
2C5Q7/4fum2aGut85mx06b7EPcN9xaoQp0Z5BFindy3ltzR2FRB42pbJ/xfF2cXo2w2jHix6Qeq0
9znlASkwAsSjUqMwpsysM5kQIvrGhicEKeQ/+Chr70iCQe/j8JbAh9FaOXRkBsRQ4dW4o/gfSAmf
SilN0AtJoZyOu+YxYCLl044P5aWggjYA4/c3QqoGCOQPcRq9vt0v9Ezx7lArezrNUBVDVdKvl016
HdNeBkGgN9N2tylOcVIctG0lo3Txul+or193/fXYXHOAAHMxYBJgWtTF9B7hANlMLIhAOXLFGy2c
nRNwXq82FUcndslZ8aCn26s67mrepemoWABwEF4AEq5HSM/Q+qaodwpGEwx6SbkhrMpeW7VmZy4g
d82P+vHsFzoUm5H6+G9JtTS7Yjg6V4OIze61SHov7tST8lzoYztfYDyVJNCtN5NQJFdi5UriqAQe
e8GiqYne/sKS6NwIP7dy5MuJK/zfBKUbw8pOtaOLpqg6hkPgUDFPWXZBDCsSH77rJXaKd6IDWZnN
5hZMaxW4y5ehZNJqWcqZE9tweXfy83e7DYZjT+QSn83G+/zTsVyZIzPybWYc4Tis35TrjBL/BTi4
BT3geEacuyccS8fENV9S3MJya6Q4EBk2Cxyp5fucgfclR4IW/j9tC2eobaZ00E/wbcW4X8dys96B
F1bWYnb1ZsSxr7IxOo+EIwZzjJ7WTU7EkgFRAgnhqpYMtcxQU6pI8oQbXmtWqRYhaY3i63uAwzsQ
gwNcp6Sa5Lxf+pcDkJF+0wT4Xr35z6TdnISJqMeshawHmDqMUoX1QMUcK+UQvKlVgDcNo2T4x0xx
HqAmeU4UzEOFJetwvNhqFAv18gmrfI2W6FygfgvEQsTNUTGYVP3b/UkP2qYGDyrOT5s8Vts55nI+
How3Acg4H7vYuNGi8x3OimUIq8O16OdcBtqDDxcKTJRKnF/AHbRsDc4/YoNKQx2mzHbeDlEoWeJR
ughbxz275t4Q/K9ubFZksf7TfaCDRadvSoYyUsfTDfYUDS4oMkcUnAqjCZEgUZe3rXI7bcEpQp9w
BYBDZSGHsITaj7R7BYDT9iqfeLRwJoySuVRrKcR/767iyD5SInjJhSPJcsb67c7TmZziaTY7C0Xj
V14M9bf179NhpcfYTGG9VQuX3EUSXrLF1Oe9eSe9f8ah1M/1a7qWDnLu0kb6yZvG5Gg+TDlkaiWJ
Y5lw9uGsThIcE/k1Wts0NLshUc8VPtGFMnZy79YUdX3eqRNzjKTvD7ekejTb4km7R8oXVV/WeEOo
ZYEhVBx72kvW0edxFB6KlxsVFtxZORpRswiUv2URqo9PjqI2CoHI/N7eQMd8tBi/lKQ/uUVccrsa
8Sc3yFk4IypwPyipUQkbPoKF+WNDwt+zGiv2IIn5vHC1ilzQL+5Ko5oCozqd3k8l36GZxl5QNWXQ
t8sPRkofl4Sf20rCevOGX/Q61btJDAC2zoEHZJQgEIVMxN1gnuv+6vKpl87MO3O8nPGzAYG+04HY
FrMKh8HS1MZUVGE+YdmySIkYL3V/BbEcYb14bQnRl/auJy3nr6dgnzI6l+S9nddYLU4BS247wsM9
53i8AwqQ5qneHdAls1wYvi0ae1t7tWKLjeXLYN9ZOgbn7/rSTgZUrq0bg7aj53oOrfaQ83ND9IsR
q0aBvWp5eblpgNQwXqFsPI8XuK0HFl5n4aULu43fgm7xu+xVhT540I51C1qnlM5Zx4VZnkLrGCJl
wi8j6Y/FFLxPjhSSMXRrJAojCi212ePExmRGYOBI7FmNYOusUQkCZWuVXLrQANhhSUF6leqapO/Z
MFGDp+kjQBgod++WyTOExrAmCnM63FddsOZuh/XRSePGb7YC66Fu+UDyBJMCiqGIn6FgohP89g+d
7k+N/QgBOd0TD7RWPyMeCTJ9ugR5rFzd3ehn6D24eZrTT7+ZBpi2c/iWAEqn3eAcjuiAIJWk7dH9
0tvVQZPDGABJ4L9jHmjODyuVz8qn5eHsU+qL8CgZvoxyf9a+RC3BLwGvJCQAX7GFM5iTKPRacalO
v1HgDZ9rbJR9YVLirxn832PC58NiVnV+4GJD+zyyvCTIid6aZXZae2VEySubigxq7/w3HmypAyuR
dMJJzc6oNy1BE5WMSDdHde+ZgOUou68fgAwa7tElkYgXJ97N23rpHes+qf2NPnzCRj28JwcnfFjg
yqO21lRY4igCHYsMOiZsOa8RCp+72/eXsGRN2HeRnWUXvsbkIhBeoA8s4F2XpJhYYG/P2nCqVNF4
E1Myk6y7KFDrvVJHRH7o9E7rdtN2IMaM8ROt01ZC6JcYqKfgImCdv2gEWwbZGZUfDbewtmeVNP99
zD36MCUb1M1dzIrjt12IzJeQHhufnP1ItME6mW/MxB0nVTDFLnBntUdemiJeecGMRirT/GE+Uifc
pydKXF+e6WoV1cif6J+l/kjh/hWgaOGdEyBz+p6HM7VhXtNNFUzrOADjKRkS9Xvu8puaPHLMca9z
jA7Es1qiWo9DJQe4NpYVXiVK1Pi5NaEvmPCOsfEg8KwWDF0NMXZS4vfxGNDrTQgPv5Pc5AiWuGRR
uO4ys7k7pyhYokhsT32vqW/BBGttz3EboucA8lhoRolBhWKpmZghuuJi7VYtiSYZ4VK86PgOn1s+
tUz6lhdWb4MirRgkce802XBkw2xbzBPgAqJkw18FbPGMxCcpmAYDKBLObzBngxfPNfztKwmCkgel
ewL8WGMbSwaL4D2Mx8k1ZsQP2yaNrvMW8axVMHdDeM9OLcfW12cx9xv+xioF0bdb2bYuZsdwV7V2
04QKCVXdKJa8EBYDY6r1htoXM4LkrIYav1kDmi8Y7nfmcB2SMFoIHHPqrRJhVHkfBJtNj77dkR9m
BZc8Q+rzfAL7OnAnQdZJ+QkK9BuH3thQ2bhxvXft61WHFpsvgTqX2iH3eVHRJcfM7R4YLhV6TAdi
xH9NIzUy35jEx6IHSgW9NwV5ni98AC/JurDxIJsbrdlBmG8eKmleST0FQgzYDokevRFzATA/eOQo
5klNr6og3pVRANYqYjhAnnjfSfJxsIfY8O2CLdEeuQqX1OMw14w1w493iFKB2s0aNDzIJl/duaJ5
zt5xygMtWyPI93IUY3r185MXkOh05rH3BvgeV9HcevXh0Cyy1yQbmuTi9Af4MG+5So2XFgqXLNT4
b8QPVJC3gxv2SsVI5ICynv4XIWy05RwGYXSqMWjpRGKy7pjTe9i99gMjHrwpG709EhyzSJ+J3Y95
ns/i/PfVJfOaIVXJNzD1s+IFBoXVF/IRdJrG6spiH9bdRZvmDS/381IgA5PYvGh5wAr3AIMWsapR
pmH1TY5bMGCLdtqefrQcDuso7dYJRFwGtltlI/bSDmmS877z97/o720OYMF7gOwoMOg/hoSRtqA0
Q22T+gHHyD/3FX5Ug7QdnBi4M527LiwWxew30Fvz1FBUfTvbbH1+YrvYVIeWzhDJeBjEp3MBrlXv
BGdu2Iowg0Q9s+Mpsr6E6rJrmRNdhjyeRH5tG1Den9KmUP6Yx1g0BgDpTamn2R7B0Z+K0TggTew5
PQ0S9Qt/tzgNtnJKWDf68M/tnhlQATrXEW6uf7AQZR+a1No86i/rv0jHag+PuTTa1SxKiDz3DJFo
Wvmi99oQYy54UjKCxRuUhePrt5Y+4mJ9XpFwk5y33ID1bKNUvAEIpJ86aXM+NI0IIvGO/ShDH3aN
7/87ybR4LHJdRIQ8XScun9B/WvD6TTsLm5Z4J8k+3tIw3CTQJUtPUAokwH0pw6pKMEafH3HMo66j
hr+LptTp8RcxvWBPjhszYHJ86Ic1jyhwCjqZ5L1KeQqTcFRPd6xdaEsLnKzH7bHu8cJrCZa89shk
2/84/BFNyDZwcj7Cr7jWtXUCGJT+sfGuRNf7jnAQGkCoiP9Lcc0rYgQrwl11MUFucTJKEdY42R22
09csTCtqIAJgdmVGJvrYwcjCYk1n2bxZq2Cdgd/UcYJZ4KbFLXElBmaetcNbEBGT50yD+xRmBKm/
q5DWQxZKXATFFwSxugoZxB6fbz7DSqFezlCgnqxWV3hVqC6DcJue51TDK17GLX2lXmw2nZz3SjYi
mJNJSBmNtVdHgAfc5j5q7z5av5TNxQ31Ouy0uc2O8/QEw/hlFg7SPYyj94XR4QAFrGkqGkZbw8Xz
5uimvPtP2NMk2RnhdBTJPwixEWs+ZgpeEj7yNG2pchPlxSiKWPd8XFhFEeR9SSiawFPHtfkYtgIm
8SvOrZtXKZBLSHpTpSd7S2PRjSgfnRp1xEeT5gyxcvGSZU90eQq5tpwQkjMIL9uyQpQFl0sMPd+3
o346N8rKs2nIh3xsitcJs9PJR8uYKt6MHVCsSvrhaDrXQY24p3/lR4xxPws5yEoibw1cF36fIDPU
nA06l1YqZWnWrz/YU7/fTN6YFrbKreR9YBl1GSVWLx+hjGB9FlXVXvWGF6uATpbNG1FW1m4hPIuA
F//aqnkxSzfFxpkRZIaWsoxUghkWdvV/V3LcFHLaqTJgvKli6hllsGswpk180fl4Gtv5u1hrh8+c
sPuA/mZnB6lRRX428zq0L8Tvp62nLgnlq0nIH9x236fcE4fTenoFjNt/Eb+hMEvZNbfGhy3n8GoW
GaSPyWmlffeHQniYuoJtWZItvu7KdQauN/xBN/TrJfKU45OLw6D4n9p1EixhD/+wVgsDPoIlHRmW
i1Uf7YA0fB0YFBLoVFfzuXBruRMjqTDqMGa5vbREzdhXho+ZUK8Fw1aftpE+k5mroCvyGkLsy90f
pbeK9Eu2zKypfDsyflKeO6u7TpvrgO0HGWYQhQudyIfs2pBBitKg326vqOD1B+KareAIQb7H0/xE
SI2QEAxJAVhtwwTqSjmwtx+Jp4V3SVAHos6DhzNm1FDoJMOm5w/cFRO63sAA9N54pzFkvB25nJyJ
cx7rgdxKCPkZvgnf/TRo1wmEDyvzlUflepAou4wK0BT+pI/hHNImATle0BQHihxOZD8bZIeTZjUN
PjmZHh3J+DqvMDQQFWCL1jiWTtfAWpQCOy9IX9nhWX2FOX5GarPQdPcxM7Q8NtPXpSlKvtKKd2Iq
rKI7LC3m52/OLGxODxua2uJ3EmhdImF2IusQb+BFZPyfoc1V7x7AvyhfEBMe5TQ7NRWiP8sS+Fn3
7ziDAeOGshPjyr4oFgytaEDwqKcwoLl98ohThdBlhfGVC/pSVG1ghYprXI09w5eQGVKxzhO+AKzI
6y4w4axKE1xwNH+StGjZxEByZW5VAvByCDLDoT23LSF7sAOjmToaP1IsGL6hOapLPxiwuw0CvelV
QxH+j9QRxvR5H7GwC2mskllVsczhX6HyLw154PCL/qqtzmTW9+XwcdF55qU4/Mm/kRbemSHpCMLM
ITIAh/01RAstUp43SEdXtS5mjUCFvG/zvK5qlPB1ZxiTkCGyjI0Leu2XlrWV+zK/GzMx+nD322Bo
XKNHmcd53/QGITKkFAKIV0H0yyHG9pVZkmhyi9V4RQ+GvyB2/NANU8oE6zwET2jjYOzD4wt44Mn/
62jWcJb3fzcCEzPw8Qvg87v6FFWEiPMBPu/wmtANOw6EBopgssXVEa6QF+zpyZxby//mYBCxLa7H
4damWB3SgYJ/9bRATw3S2E3R9zCG77hctJR1PysSSXMQE35SEx0FWRczVDwjy8QLZ9djbN7E7EjY
CWUgpuemf5xoEJ20NnEFkxHkoKCOwU91Xo31RmtCCpDQYuGU/N27U42YBBbIfOG5ejesl/VZSI0M
IK8s3HGp0Azgg1AOp06PiiNHvWJsPgZ8V7GfAuPJsAhBoEbxmj8+90NWbpjH667jAQG2/op/tAJG
oRYelkH8WJ8e1cD+1Jwi3Wd3BleLgPaEwDUc7g0Q7RqC/RNKdxmeBlSKBI4HRP2XzRJU8UtBJsAA
yAn8KNfUI/T11K3l7RfaSSlOcZoIZF56E8F/fYelCvrGe1410UgsGS7CBwaErHF6TBexWSEuEoWi
q4bciNqt2t72Cr+Qje9jYZ5GoxLCapLZa/7fp/XvQyRWQGhmCACvy749Blh70I4Vtuu788OmJnbj
2T34M6lRcQvYvtRoYhC8cS8Gk6ryaYC8ioe6Gqmtj8CIs/JMvvJHU6qobbU72PdCwKzYscdYWM9V
W+mdGklaZJvapC2wTiC4yhjPWLmv8b+qPuYonlsqFU3BGmB2MImqWMY2GIEJY2DarG+t3UPA0rrK
IzW0++O840l7kKGNnqOn3TRxyfp34CRsf8ibBjMeQo7DoJ2ZnJsZ7h7vTrfs8e1Nm4B2JjLMvM7G
zyYiThobfKQmEhpkSt1LVwndLFmLbg83G0+53dounzYQZJ7/04nOBeDXIv5tYEWroGT3rGLpNbc5
NvfxWboXfxPS9WiBt9oRKXtyYMkizYU31rX83w981mJ2zBUdLBiykQT/hv8QeeU85MZT9HRUJep6
wVvuWkxzcihtWGPqlzSCxnCwu9Qgt91s86HHtIQ321LZQggJnSE6IbZ+oTb1xr2WNoPl1LF7lyKI
5/AWtCD6yeAmUSrzn1K/fFN6iCRt3/nI1VxYbBpTLpkL7S+z2okC1KfSy81OQbn5W/QRapJhyLJW
MQvopUEQl+bvQKpE8whH6CBnhh9W8bdWDj+DN0x99SafadcSZXfji3jbw4p/Xg9ba0T/ftj1cHV0
imeqrQmkARMgkjYTIMMck2kZ8PT1XGjK8HWwmIHI+H14GRXv641uAkL9yJuRNYozlpedTk1iL+ph
v1nd8uHjdEUhVeWSFYtLwJ86LOt+FZSEv6BDOOCsu2Gku0w3choyVqbSXbGS78XfdxGvPx34lN77
esx+O2VVfAI/jZxG46gm08JhbV3qhf7lxp5WMj8ZJEXjC586XEPqCDgTKIJW1dBUhJDJAO9t16xi
zGlSAO2Q1+H7QbkNmpmLqOUUWm+fsQdwIjeK3jSAFlJiCoPKgh1+93eifl7JdskPrqLerEKrSBQ+
P6Y6NBCD4cPrWJqWopfYNVherKkUyxwSdiTV7PkLpb1ErPVfB8OE1dhQOsFwQXHLhuv9CirwcsbC
fQzQGKYj5CYp1SpRB+8eZnH9mf9U6RCVdZ2HVt/6ByhEdEA5ZUI6auyQEBsNTW2csdfUthMrKdf6
qZrelqINanmB0OMOW3ofeAyV+3IPmKd/4C/9V7WiJxMRn+aSHd0wwinHkpcdlQpRyFUE1lq1ZOnS
sdwhvOlnoZ3LX8gfXqP0a9wsTSp1AEsH1UC+NkHUh8tbMgH2c0YIAEu3iZsMpZGTWq18LSotiLbw
wp88lqD5B1fD1XAmz7tMeW27r/XBsWqO7AqRi0SL7ljbFZZx/c/6uB+er/lMLyX4vBA+IYvnCzBl
ni7GUs+dni6SScx09WDZ2mdwo2pG4a6XATDuVq6fm9ub3Ev5C62QmbrbkhYevyUwfLVMt10oJvWd
MfLk56QppZ9VaJ/f1jiKFfBdIf6YwSBiR7RMDZZKlmza7ciuit9jRDsEVLC7GTpzMvOzPPJ3IRFK
GHTJJ4dUuMAbJ4iC3ojcOppbrhVFdD/s+6lNH8lyy1kNJEvd83C6lJRJDRk8qINCTdNICdX9MugB
dG3GEtKE/j9/SrqJt26FduYYmQqog/P9p3Y8JEuPBKaH88eow04XyCGAPBW34RfygUa9g2cIuUON
BER5REEK1l5KGFKmL8j1Cej97xmZ8aKaKud46OKh5tECRtdqtgq+TC945mS7kS7wWVxWS0Pto3kX
hfPleGCR9td6MA//ZTwJK6Xdht5KLuWwZwjp44pPl/BGsSCrgcrT7Dw9VkNDy2HTpizggoIvskXI
TV+YCfKbMwqyevhvoyFlntrmqzaXESOXoGDaOfRxuNKFJ4/FMASwRNKa0WPmdrNFcGnHmVoXio2j
VMZwofxNk955dRcRS6E2T614G4c+hz1fnreJgbWUHoZ8xP9qQZNdAMOOk8IGd+UiSVemIiieDbn4
wA8PlGzUi3jP74aoi/6OmdBxVQJwg+62V1OFJ3jCGs7EdnSLOpmZf9uT23PVL3jL5GlmrDdTN3e/
5r98l6iiZIiFoqRuc81AtI5vJbf7iwhxG4+pcYLHFjMeFX7hYsdl4VBKNTkl2KsESrQErkS9qwDP
RQO2ACls4pXOXKPehgHsLuXLC4SvPVngBM2yOeN6xb2uGtMrcQjiEQ1jYFlmLF0//CzLvtDLEjjV
xWeRvts8qAatesN9fe88SIzrkFhPLaNaK0RWNOb5YbKo29gd5DBGLVrWAUnM1JLhC073YZGhh4mA
Fz1pJ6y5a7t5kjmMg1/Ulqw46UHWKVL0Ca7obcAwuIDAKOVBji8xBZn+yAhmSVdxRjjm3BjstZhf
CilWbn6JF1jcG7au5rmEd6Ga/R+SaLzioRQoner9+xiNvFlhjRs9C8Ya7FCUOIvN5jNm3uyTFmuO
fRpEY+nXVSFPD/JqHrt50SzfmdWGE1xlaX1Q6Fm0N1ivc33Vak386oASAzERBaXDf1oD4R0EOSBL
uZw/VpSQ4f0KWLZWl8QcTETTsVXrREjkICw2VxZTqujfE84OvBt3jgT+GD+ICEs4yHx++8DnTgBu
FPhxBX6enfQUzDsHPlIUzSwZ9hX4RKucD+2CtH8WwH4Nymmvpy3aiNZ/Kpsm3KI8CjJuzeZEVWKN
1V3zn8U/IEy1gFb/Pu2vGXXKOoE7IpJ/4jor2c8n1ejss0zyJeNG+0+jvo85Vezr8HcR8suSUw+c
NQc8jpXDrbz3uU1bJmE7Va/8iGGNT2xIroa1e7I9TpqGKPe3iaXEgLZ4dvQ14bNpMDwtjhoVce09
t2mL8SSBgeV3buZt6+9El2w/IQC9MHgQqhk5yLRz6BUa9Hf4OmvkS42oUkaAbd+9u50kL0MN9W5M
nNYu0+6r+PPXygJNxD+CymcF7TZGviRKSrSkjLdR13QX/HkxiwoEBvCMJDVylpopT2W+FIz+vOQG
f6rSoOijW5mKetskfkuCUS6XVksnWs/+7DZK6Pa32ZjRCf8W2SSIYa9wXTv28MipyJfVjYGpflYq
IcXZbK3th2YezEQV4zcie5/Tt7vA+AbJIa5FYvk7nQrwrC+Sh5CqmCC+eQW7/w4NBdDKAq3xXf2q
I3OCuP48wI1ZL1YZpMVh/f7GBeeLxZR3NoEa+2LE7B2K9ZUD05TiXqDpCdf0PX/cDth6+sDQp+xT
J2TvgBi8r7Go/qhGyCE4D3P8CoQFcXf7GMh7MimLdRLlzgIMzrLFcv/LxGERaEOx+eV9adcEF+vr
UrdQ85J886JWgUKJIEyZpz+K0QoF2XxUWUnk00SyIU0qqkPuQT/X3ud2sZmX7asRbYcfJN/7t5X+
XGVdZieEGTOUR+skNp/hGlvJQOXTrBsZvjRgbLAc58QGq7McnEfm2PByYLFYyng7eXonBWr5Rusm
lAJK4fCeKAHXbEMQWqjM4ILJTgxFiDytoay+UYs7E+JEXMYMWvGOgshSd5HA0zjH/NyX5TJzEl/H
x/xvnWDT0va+Cxt2omsci/FvJxBLW2fhdKxMpgHrGj5BPCRrrqhO8HFDL3BePw8Rys1VKVXaXoF6
EHJvG5uZaIp7LOE0VUdwYQQ3d8lkVtn70afI/jn3racI/1rHdixdX3clZWcqHt9ugddSETC+HCrz
zrWr5Vq+nvbVjdPDM//GA8UjK1prH7oFejAWSnSlZZZs2VJ0NwVOvqYO0FFXUUa1s1tg+tee2wVk
XYZA2p+g0snN8zJcOoTLhD9aQE1uTvwsWN1AxBQ2wdMil6hoaFkXWf4eYTai1aGJ2RSMJiKMoQoY
8uSndL7Z+hqGgVk1dZYRkyjdQ//Luy2b82jGxchaeBdm42X8/CKnX3LOhFbpqbayDdVjw6b7sWLU
wZP0G0wtNxnP7lkb7bCznIQP4A8ReXZEP8HvnUL4qj1OA57w4RGlYfm8Hh2GnPR/0eXu+rQ/yQah
KpaxWSxmSkGcqLDlh7rYc/B8M8ulHtIyOJqFwHUK6ELkPP+YBZeIKZiruCQML6+JZ3rZa/aoJ2VW
dul1N6FrdCxVq0rzrZATc5boDu9yo10OAGEsXpudgZMVWp/B+S3Q0qlzSzCTiw0S3wV19BIxX5X5
sG0EdJhx+lUaIMiiRSWwLQEytzvqma0OKsT5vujs/arnLt7uUH4q76BTZFib+eiHYQ9W4WNrTrma
NV+zBddjCk8pSpKJXsGMu0/E3Pbfq5wgqygdWml7aMWlT3WcLn+MlE5GnLAvr735K4PMKsNdDByD
rdzSPJmVnxpivD48abyrZ5S0F1nEyFNdLYSgnTtgqAB5PrBrGNRddY5JtLxk7CJTeCoaBdJwk9AD
ddJXEMH65pzDmrxwSGALatzEnmAbKuAZUz417ApLg2p6B7Idfooj+uISX+O7EHDC1c21cA/w5wCx
D6JTBJZw1RYTbv34yzcjuJaXjf9pA5H22cykeIsG9hfOlzEFFUUwioU9azrN/C+y7Z1zD0Bf0ux6
YnzVN8YNyqPv7j0lX+hDxXOzUyuO0a5AgrNnIoZsAprBGS0g2izEn+aHagTc0qw0xTbvKLygjrRi
xBOVrihyz8JflbzfKdlZP0xsdKsZikXBcFhvfFVDBjVclbYQmutIbwRxUGqDVD2xDbx1d2shhINb
DnQkEnlZZadPRHHjj1bk2XXdIGfoV6QdA+9yiwn6pJLr1weuYcYUgUcaWv6xfmmmMxiW9z+XsqXH
jNH9as6d9HwWqy6SMzWpWgvknfDtSEvESZYQUZY1l96avCssyzJkvbGAD9o9KkiXXQhFc1WIro8v
UY8UGZxv+ACNxIT2DsinqX6ZqiDUVIswgpSn9oBof8d4Kc8XVcKHmAcYgcRnvHocxPBBGoN7MG99
Ik8kanR4cvqHc7LNTgze6Omnmk3bvKpTFhfho/Ijp8daF5y9i67jIo9zDpriB0wYjtYO/Jaq+lpi
zXYIgqn90Ha6KyK33AMqt1sO/rSofakHzEjDdz5hqQLct4Gm1D0gTuRphthJwvbVTWsVRw6/0FeI
OrwRrJABaEG1+6SDQxyu+7+sEE+qHwOr7XWQQjt9O/pBqWRpR01iukJzDwAVohMUNlIk13ZKcQaR
aI0qD0BgRJxlQl5Um2Nl/9tvT5qi/Kbv87KDNyflDuWtl/LwhU4JyWmrwX3EbtKwo8H7kgU7eOEl
P2Z/06nQEwZ9zZdEYn2knFhnQRjQQwCAnlC1SntPlikhe88RB7N/VObVIMIMGlC9cFLmfw9rvdgE
tTi0Y0hiQQhQG096wFQFo4c+2vyDYDCbMe20dqOw7yu46mzceFew99eXQhdVSRBhMhyHO2v0MVrA
PXIw8JT2FZ4xltZQtSlhIVpMFEC+gjM0wzfFOUO1eu23Cmz+j6eqrNXyr/Bu/9dJWLiUMWrtoa2W
HqxsQXSCzt/orfDfgz3AWHwW6zfeW1GFiwldnkKQRSjbgWWAmdatcN04SB8/5J5I3I3WVpYY/FLO
pqZQjFDZdOIFcEaYy36jv9X9KDV+jjk7FMSQoKdzO53RfGycD7d9wZj+iLt4HkFrlVeV0i2dpIIJ
/+ULzEopt1ckeeaiLDS3izsfRJwMBLkyl8Bwa94+RWwhZpbtATty34YzJDd/cvrdxc254oui+PRt
I/1OcBDda8yWLvZ0C4O2s0KVYsXoM4O0DN/6+bNG23LWBa7o5HWw4Sx2fOGROAt5kiW+t1tLK8uP
yAsp0G3cTQS7lU1F8z05ssNwXXmnKu67Yct9Avq6v05a0NuAONPFF5S0o9//XQuF123u4f1WNODu
zLdMCP1nSd1MgPpj51+h/eaTriAODYNyidBCZ0t+gdaSnvM8JqGboz2Tp+uVe03W3pzHkDctW2Cg
GqLCOvRLZ9mNygTHMaqRIFbYK+DvK5S3Tc0mVgm3T3vBqUUYvRlH/Kh5k/PR6a/cy71xTx9lr83V
EmGbb576/8FfPrR4sNOf8vikXzKftQYug826RSdclEmrZi8UDJth+QBhCI3ffQzhV+iuRlDRFB8Y
wbJtMNcE5trucyPlihFkiaimlXKI4nz0Ad8p5bXfi/md1UpX3YOjLDDFTOqpysVNPLsZXg695/E7
BjL+snvmuHeLEQlneAOdHRnGXesBZmLMGbD/zbfaJdtub0NkKDK7D2dCVU0GTeLy8qvN4cWewaN3
qHE+qv2K9ASyRfOjDe/zfHBQqeq0vJYx+qlLNOsJcHnCCYHiyKaEfwPaJnPmAuBC78GmUlIoteeY
Ug7iHzkSyvUCU/lXSwGDqJ/BjLvAtjjDOoSNEqUDjGLiXRKZ3+cRzocbEKuIPJjfug+OIj43AbaM
ls051lhEIcmMGnuS36N8Ief7LpG8zx5aJK2UGTgIXsQV3B0d97Vr1NcYewFuUfyRweHC7gsbpp/x
QhHPTi05ZWOPgIdKj3QCLBTbyD76KVOec3wkaKVRFJBsrMH4GB4jqSlP40MyB5G/Lbzq9vSt104e
RqteICb7tfO6iZ1uFe7hpuJG2OHDJ+48BkMfAe0IdIzTHSsFGImXekvaSikjsGgOGbyDkKQc7Rnj
8+TEyM+Iooj8CudeEK8Y+8nUrzRnxamvk2SKxikN/jMzSWkTNWmyYK8Jq7IjZSEfHuRR3peiQhwA
V2fSi6aCq61qcNzGWgaePI0uub/V8abY2BWiGPbmdxeHFlSdMQ/CB7Mb83ljCDl43tKLrkupmzIr
m+2Dy6jeo58gAvUwLEuXsTev6d/7EBxu2W6mM+gVonYOOAdpTsgzTaOeYfuA0Eoo5VudWz0cnoxK
09nk010j0Ltf6Jc4lD3dGOHK17zDMl494nBM/96EQ43Iwof9D33R8RKyoMk0AOq+erl0CIqYiKJD
nJMyvZYi+z1e8hiNNMfZMM7sF0y5SMahqmym+x09N/Wc0+m9xVEj41NcW/dKKj9el62c39a+rtAj
+3UzsUrPr01t8xsY9miz6aZoXQx8pvXoJZA1EOYTRG0Pxb77rqeU4Oc9US/1D3oF0Rt3c4LlpeKt
4UzdLIZhUvXjpcbAq1jL3zhzn9DW8X6gJ44A349+rOa5QbYFJt4WMQOn3yy83RqDghQ1rmFoYNRX
qcaPajgnGHdrC9unAwLjpuVYmjN9KNGQV5ri7BfhjR8d/TVYz0AO2DEj4biske9HRWHTzFSJVuYy
mlF5TSCs6XX4G3kOaN2PCKky8tyVKI/YBc/5iljbW4S7TEoksRQqPdSLfjPUOEphkgfmHjtAU+jc
IbT9Spg9PKRHvwQgTNn5tUw354E24TND2W8zOXLemd6lbptTafJI93bAVnp7XysShE03sNE+TY8j
1PtOsltqkd0TySv9DalNljTTzNS3gU3EBmZFEqotfEn/rdThlkZ76Jp76DzjPP0fh/rvKdsWuh8o
hIeiO9x7bl7V1wDZAdyCWC/kIJ8HxC58bZsFEUrULnkWGM+rgRIixlllK1RGJ01YtIroDpom7i+C
SxJKaNzItYTQ7gCxJfo6XfORmDWSF7OOP8nYzCD+fGZ4a14848ukSHzUvZGG+ZsVvSpBrHJXTa8d
I1pzf7orv/yTGxbE/V2TsNl2o9mKSPqv3FZhBNYdCGgkplRPpzhRTK6/q+GCl9nXF9F/w4VYpdfT
cQ4gAF28yv9Nt1TjIheWZZGouxtLb7MKyBPq8dAnvw+FMuDctI5PJtFc2KrSIgE7Vu/2Kle3+Yyo
pcFMK0IEcqzmx9AKwSoqqm1fkjo36frR/4pnyl9RLwdmUwhcC08MDLKh93g8WJlpukcZ9WPBW5Qp
ZEjiND/w+W1hSKjnED0Q3u6NQtTztIBIpEyRerfKLq0qCQ73blWkfx9zqU00OsRHynotpMJ7Kdoy
U7SDhHnzkmefB/m9Pc1+QF988xad3FgRGEiurqN2Nw4MqvLDNe5YJAhc7yglmNSUKGrMSNBhVxD9
IE9Bh7ORyUA1heJoh5q9ry1WLC1I6/cm4GAoRB5pKeE4l9TZnRKDUiDR8z5dJLTxIm8HWRt5aZxF
DODuu7VZqLG61y87w+78r7lXV8Wh9eou13yADGEpPcqShzw2b+zJCknwsqaGGl/eTMJ5Kcoqp2vd
VuTON3OzVsWcAx2Wj4teZDF9qt8RRl+S3XJovXbHygu7W+2H0FvpRirT7GqBn638PdFl6kXuh1jl
Gk/+4FEbmRf1EoZ/j7AsO/qqI703RVSmp/VXB9z3CM+WDWfwZyLGMkkF0ti/wt7xdd515vXBtdLF
ucW7fBE5Q1beRVxq7q6L4m4QCCu4jJdDHm05ZG0k7JETsC8QyOUCun9mWBWCgIHBagnxmOyT9Ja6
CBOqu4kQHlBKCiJenzCa1gmj/3Q/qY9XST9UgdLFD0fFsAX/1l1Hhqtj1y0FPh3oF4I+T+hEkYN9
XeZxyLaEkc18a4FpSn3PYthws9fVlqX0jHxJfC5RjSz9F9ptKKJXo7RGCTjibFT6gMPrWEAMrBiW
/YqFh8E4fSEqQkt2VPS3uC3OAGFJSUB+14h5yslnQX2vKLTHL87QQoiqcA25THyM0O9d05nLgIeY
0OeTVRlc5wKyxlWhz9vzxWnBmu5PyUomLMRbrWXnxMmPWON4yT1nNUv9h+ry3DydFAhlBidiOYIT
9CIasr6KkDEOASGjPw8jSn8ZmpTIuMH9ixAh5jFXmXMD4EDAKvmR1IJl5GkxB2XlR7exlOY2dDvF
u8a6g7NjfBJP/XhpvJn7oawKJ6g6iszA4RCNUhEWGb1XTZO1BSq1cCdou7j229hKQA85hw1S5BNq
ExJTBxqyUN5bbgSJ2wFLmiiUn0FsF5tDNNhE9lR45bx3UlAWWMRevQdW8iCQu1AVmcKrslT4gkZ6
q8GkVDNNoxaYI+wTQzBljs5bFDI1P5iNhvSpSLm1o7CHEj2TNmWjkZsWMKDqyuzjCZ5Abe3MyMzZ
3K2ZhYGjHg2Xq6sTjnnZtYymlLjL8RtB5c9zDJWqn6OfhoGRNnY/+PzcHO/Adli5/m11ZadcaFAr
yD0B51KRdit4hgos62Tar8nbFWRHAJPTVudxCMo0ieQ3pI/u4WuLCeE1TwQSgM+tRqmTvsKRUGso
YpgFjR6sdX22uNH9WRb69+JZ/oKBGwIWDhZVDld4wc6tKHwuENFuClWiKNB+nIQrATnQEY8THCER
ZMizJ92LkOlphT+Xxe3E44PSC2gkXADXXtMvyaaz6i0goCdzQjM4us1f+ImRBdbUFqyLU/ztfD5w
hkzxotymUgbSwJcbTTF7hmElpk0yQVfxrCc2r/2FI9EtCdlNqQQXZMkthEnx4kl5jkDV6ouircVY
vnQNsprSltRnuJ5uAJHVaKPEdMeYQoWG5OWfcV9IVItmc5Twc2QjvfmNYIoZqaWrQOna5h0eSHjA
V4cDZqwMlUE7wNvpB1IsNTxKnlY08sPeG1B9NaMXduWE9aQoQyI0VZi4YrhV9QSDDUc+kO6Q8Mdb
aXKtb6CZ3W24uYJwARoAWMg1i3EtdclH81HDcrhJUQ0V3QrvTVOTME5ohGtH2427div9T/kDr6oV
XTmc/0gTYlqh4bGlFO893O9lzzt80qOlECnaQnelYHyIIFuLPknBNUJ8RF0CTCEGj7FgeHdt6pMx
b5LwT9xYu+nDQO03Jgs7mcNAt5aUicIzSp89BYnWI9bE4zIgWu3iiVmQFSjBP1TUBFOqvY/WwzAR
fdzbk2BtJ7byAmuRUjiyXR5tZ/aYpqtbv9GdxJja4Ro9t79i+QxKijpFR5+4Ye4ukfGyqt0a/qMQ
qFUrOYi2aWWkwYs3xXeKyVj72oIQIJXuNwNDM7zDPIgCowdHIv3mwEBepI3A8veEBGGShkT8PH7k
BKsrXmtEb9zkb7UWuLbI253xD1vVo2rjWnMl7zkEOF7IL/pMbIyYbK1vephvP22mvVLfS8E0TtvK
Qqs/TO5F2vk1kNz54MWQeLRFXlPiF+fY/ZYAAKkEhDeVHbTbKhGQH3yoG65mtjl9KLpR5vVBITcI
5MNSKcV35TYFw3Ln2Rd/1htDrTn+fWMRWJtQ0sXY++7Psu/I3T7kpyrLKPP2WSd7Ys042Hcfh97d
2cHsaIDaOelQssptRUXB9X5HE08JRTTzJ/R0CKg0L7T5zL1GtL8Dc59H74mtcmlA8l9uF+wH6qAh
h9GvGx/43WutCty4b9t4PYAC6RXxPRfOxSu5Cg0ljfB0xoT1XLaT/3Cx3nDQ1SFVIQhBFuxvDB2H
p28dgxcjP/QtqTVMN2KxbQTK5S84MKbQ63I0igM2PkEzUhk98MoIJU/CoIsDdz/pph5765y70F1t
ma8vrLepfzqXdUVMRbnAHkDJSJHG8lZpE89MlxMH71TJ/mNdpplqDY7k2cRSd5LSsEN2HFbilWiI
T2JxvxGT89Rbz+pXJVx0hLBdDtEwqyNUVIqzDmlCGsQwGHAA6pK8Fzh/AGoV0wxEGnRH/6h41tZX
7NYkrI42YbZqhFCZtmX7FVRoP/D19Zv66xK6B+UkA0d6Z3Y546eTsrkWhs/9dgCWBX5PaJlFktAZ
oGBefQqMFHC8S7CfoEGk94pTDvg1S8y0H2/HgbZW60GVKeZrcDIflv0cBIT1beBOMWfp+D0g2cSp
hc+1InpmMc68JCyKD0oEpKT49u8lZ0rocyRoejKjGNkAEtuMcXzlmdLHTd9bU+toggWRJOhmbW4H
ZFbzI3oxpJPzxglLGrMQRTqOeKR4jvZhqU8mCjQGKCX/iOleJYYo+De/EEvgrS4xErUaNRaWtosg
3L5fsT39zy54gZj6NpVCYDgmYn/GkcFTBcOblBcmZ7FlYaXtYt72XnxsVa8xRszCbPF8tFg/m7cw
dMn4gULKR4i2dC7IJ0HtzspmyEyG+b8EECouaAqefMnWo5JfUjTaPidle/uRjNFCeM0633vVHoX3
VVQaEFakkWL7CMTQYDTOdxeWvbG2/p21y5EqLvB8lTXyY8E7/sF0IKkLZlpi31MHCLMOqD4euxBH
IvoJrkmBuYBbn8JjwDVYURYr405z57vko2WYi0UsJ9RG7rnvVYGM/fhsvlx1K1nQjL5roeZmPAps
UIdvI33v901aRQZJcT6+plM9R+DL3GeZ2G3YagvrJ5mKI9t80mydoVsXQoRxFex86BA34gcIWOJ8
TcMT4SRL0yuEb6rOp5yYzyof8PwP69khr/fiQRdaE6DhnmQj2JWGPzCS4WXEfu8CfNczBa2Q7OC4
2cvMQogOprhx2wYeqNR6eTvHhEkbWbYuUm8V2O7PgI116Zd1rGxoJfsMgI73H7wsbhs0CRP9w38E
URBN2emxZl1XiN1NTkLplxO4/0zJLuk7X+JEUC9XjBQazhZr0mslomzYPEqqV8kixx4QRmXLTtEG
n9z6Wd9i6G16o4EH3K0v2WmoS30gYW+DPM8PERcnOdlbqlLJDKkZJbFZycVMK5xBcj+dpyoVOCWI
7QrflFzKEBfrvvz4fn9Xgyqn60iMNcy6TV/YT1QyPCMsUTsU67e48ZhRAWZIWI146Vm7Q5/u53+H
4M6Jh74g7HNSNZAg2V1aVF5ytD9HAPL3d75ZqJSTGy585YYqrubEto+9YViX6bCTAk+vntbm0zyr
G9rRPmhes0k6jqQs53a/j7V1UKBeCbWOtGyR1tveqW/Jwol73ZfZVVXXX43zBFLkJgJfBatu7lcI
bLsbkdbkTSF8hKP/j0m3MiI//s+LubiDr/KSnIRdVBaAwjVZOFCl56FJ2e/gwaEjgzU9DTF1GZsa
YeCLlGe0/5D7DilKBoGFkF5uN5CyUOgdXLOY/YZGkx9O7TtJOo8GWdL11PWQSzhrEyTKSH4zS416
0A6rp8pZ9NAUWFNGHA35MuBHdjqBgZbjFS+nGC6y3aoMFsBILKB3BD2U2w2HF9/Ly6a2xlwdLYwM
7JgtApaqPxi5riZJeDV8AAC/ALtkaur5ySmBS9jp3Nq3GtOCWi3VMFCXz7hWrjrWz8+wmU1UTCb4
0KCcFPr60ztuAtS5EeyEwYuFIUfyE8M1Wfd6675jjusnOJCaXlasXPZM3DFuBSjtG6Fa39nX2Z+R
tg75Sn95hPEfc/Adu3yTnXbELW3hzKRkR2/MrS+Lm/Jqhu/a0m5q7C+FhwGme7O669NIUcP8VWP6
i8+bmrO9K38vcYesuQEPM1Bj09fRmKq2drPTHnou9OiHHIKWyiHO2sn6okn+kA97Z5ge9SMSzJ4W
SutryV2oDavLCQEtChWHO/clOLVM/cEHbaYLiJrXZg+uJrVcmhB5moX7LykUJAWNCgMs0l5W5l4J
EMWa00X7V2hhmim8GJXXJ6aF2pf2phJ0zQ4Hibg1NPJYM0lXnfnhFhjKGFI4BDs8ibuq+V+43DoC
zYsr5kd+4cToCwzs0E9bY/Dmk1MMIX5XIDEijKK2rn9iJwiYshzboNZ2Jij1EYIDGKiGWzV1svkQ
h015HYZPTio2M0J9c3+1fEnAA5CO/rAqYRcymqR7SGyd+pkA+TfIcg4W/DV2QoMdt8rWhkg9wn7N
nXc9S9TkEKW4VyXKDinOv6PuuUF7PVhiYvWbDj8k4rBs/vfIMADIBBQ8TsbWeSIoXQi4lYnQ0ZFk
uEi/pfYhyYQSsez/jVX2UJcPsxvNFkHnirXOKi5sIvVU5cQPTK7rSSE4gknP0QFE/exvlNTEWzfo
ty4cJV/jsAZCbaAqpzbOgTNRD2eoCb9fUYwv9vaBbzWPWshoJH4hALU5FvjTl5QAec6OKOyzW+cZ
2h5xzCcMTz9yAyNKqVX5pgQjnHBz9q8GDFOxW+jtuyT+zRflZj43PiDQIbRTG+1r2Krz/20Kk0F4
v1/BGPua1kfPpLxDrUsLLIPzyJtW8IDW3O4oRuSugBLwbV47Rh0mkJmEQQ1IAo+DwuCjYrw4puFL
lWHLAex3hrZZ5GVsSPdBnmXvlm37BrCOnkS2x3nKuOArrXSaPtaxpRy63sTHtpacuNSGaBKPUDx+
0zFgdJLNRoY+Fatg8UsEU6SfpluYTLcgG/6kF5czwGktz00+ANvOfO+/O4bnvvrq/p72ycLbkgHI
9vFcGQ07q6XxQd2sYp4MfTDVm8hdSWdgPnqUJegTTXnEc4c6GnVE5lKU4ekDE2zpEEHUIubhooDz
wKCL5eVk8owqRABv9brK9A1WGFA1qSLXLMltC1Hi9DkjF77nDg02UDBqwHZe3vLh4NjkPtCWNDSc
D6fA/gQ89HK5MTjFCoIvNlSMdCBvXfTFDR8/YBZcR8PZ85x3PF4vSzVdViXwHRDkDJ7BpKPb5Jbg
u/rfUxOhYv+uKBom2iTrV08lrZLN0idaFrpbRLo8PB0G3bbiZ5+zumgGmpUPvely7avgYX3aKg1A
fXoAQRnNBsUh8rEGpTb29vAQ2hqhY9PrEpM/8BMh4adVEn4o1snfLSdGhQKdU1bsTB3tTVoRwDew
NvRPaUwQzTrzhiGzF3k5pTrNNWzqrUFNqPQGi3r6/pIS1RlGajAq+fDLPcsBlv/ln+MPr7rUyAG2
lKifb0ZfPM2D2xyqr/IPlhqT/IJYQ9IsM+SpL1lBugEfdz/+pRquf3JAq1tnmK+pf489hmErAKDA
SnTQSsbNmedIfJwXUWN9Z4H1R0nKKLts4AtGC0QPH9N+CcxB5+WmsRlARCjE8lUR1tBEWgYMH9bP
UAQmFFgoMnqGjOPQvJCqH3CLQBw+rnxhhyatV/7vRVYhggmdZYUUF7LqxvDNIYM1zQRIDrCXGP+x
lMbCWUztL6YV+ApTjN8RhAZuw4Fu5m52mkTsEiIZCGPYsmdrxZm5H5vjZNU9NOg3mTQVc9eYXWmA
ub+m0yJL7J/4zLz/40dyZRpcMwxpLRdEEG6mzOvIeKkOLTzJF5MLGWu9PmGmEX/beYK+hG8Jw0MQ
v67ZyWG9mSAO1y004D4fnkv6zKM33S4/K2JQ+a9T2p5nfXCqHdNJdN6tdiUHCrRfRbbaGkB/ywno
FIsPliKOcIZ4dBxdy0D0xOC+kPQOBZ0Gbf9OrE0FADg0HxTo3TW03hIo21/4+PYFvFcm7JmEoKXL
K1x+MmBC58fh5LhO7OCiPuyERVzRjNpw+sLEqkVtmjx4K+JjCmNSgUex1r21yNX9kLN6kKYXsFtf
aQ3e03etnRaE8KVFXYDh2cvHqaq6SelMX7fkepTAqlpUakcW4XCK/9By9A88xIGjTYeTupWYRaQ+
7gphMyV9TMg5cpJ8Fk5x8fj/QCNBBuJSU0P7LJhC8UZTMvHLMX0ZS4Pl/oUJTo3AJFf3PN7vzGbe
M26bOMBO+Tc+CG4V39J+e2KZGGiUS6opNKPIqax4RIdngXfedooDX+BEncwiKLAwZHvm+GP02cpE
e6qsBZmyhck7cZWYSY6TCHbprDunItM3p/MudSgf/5B4ZouJf8LqPxvb+/eDhOBzfXQ0sLjlNRCJ
2S5g1hgDLvS5N4lsUHsllZQlydmhj/Y56KaApBiZA9Tn3qU3VWfFbhWRivjOPbdoMae4EOLDcmeJ
0UlyYtb/aaERX0UE+pOA7/TKtbD3ZFVAV/bJv848AvRTk/s3/cVFm8rMmvqOxIN6Mmy14FGf4+YL
j3y8ngLCaJUsxIaLTnZcW+uW/IHackmI//F0hqECg8wfP0Itc26l02Lhlf54YCdmunbdPfnCgVrI
teMedZTvSndXJRiOdzk8S9YVfq9PNSPh3ACIV0PQ+Z6WeGapFItq83j4+dU8hkb3b7NQt4kIUlXT
j+6Z47EnhxCscJ5+8m8ENhLEFsyG5PDDcLwuUkPFKUhotgyS955OFqeB+tV4VtP7kJUfynjLGr8P
iD9ycWof8aR3LitGdguu3Fm2vsEb0b8dkZz2xCpKn0R6oRacBXmsRPaVluyQd8DwNmlbdRgDeDMp
c+eOnWzNV2iHLZAycEIDaZdO1PvYZTAwvfOW7LKOEWMV/8N+db9+mRp3D/73BgfxeF+zthyKm3oC
Ia7KcylMojMw9OiPl0+Gk2caeYwv3gBL9PbCVS9X3isOy/Cml5I0By+wmuSgaqebDWuLY9zCsCTC
Au82dsLGV9WSOS7HOdq2aKkVgrzB67wpaCPSEV7vJeShdq7SI6LMDv2xFByvFr0LdXUSnJtqoCj/
SUtmQ99uiMIfv0lgOnahctAlZRDxBqqD6K1iCJBGnZuIoW4QPM0oh0MFB3ZbzkFInmUT7i6rBGoj
g24sDh3JGrl8d7CC6vbhNT0QQeZ6wsUAF7lLpQzGXZl/2o8Ju3L+iTdWL5fohMGb2X+Cm++ybOCI
ewvUn1nUuDZM5dieiByOjNJZP6Gc3kk7XqrcsLpfk/g6H2Ou0JWZ5tuLRXBttmwIts8eELZ/5C7A
Y3n1FNWLEqwvm3frif1MKSVGtRXodrYOy5Ww9Iht1eejv6L/HeuTudz+/34aeuaGlJ7aUtQTgJQ9
SjkvuVEpXoXIkW8GOQOF9DPUxmiZBqXJmmCNW48NnKt9lSD3AXPz65EocR7LnH4GTEsV3zDcaDVf
GiZT7aYK+xLQmXb2ndChvAVxhz+h4OrZPcyRq9VRIxMBr0nVxuzOttY6zF1GynjCH2aUn5DFWTkb
KL0lDFmwwGEuCSsEE+jYQRs6J1BN/2/2phQcJJTCqH5Nhkcg74rksDbyuF3klWvtTDEGzF4sW7PH
BbRVJp1Yu0macYnpb68cAvS77/u62XPjquQ2DBaFbgnaedhOcKGrLlgjHlKamsWwcpDZszAmULR9
mDjCUdr1IMp52J1Bocb+KnYtRIdH9ocu8ib0GcgY2ps18j2UHFQy3H3hrm5JFRJNyxjRLHEjjFWN
NXV8gRwK0+ntDiqJ9ol75vLZ6KpihFylr/Ldgwh6Jx60dc/IkXsEt6Ox2SYpmjwQ+dWMb6Uo19HB
ytTOMqxsll7oYboDry8PElSKkely7hdwBdbrlqceHffH/pH4v/kXi1bEKL0z66jeG4rr42h86Gml
7JI9kntDUFRvml2SGkmw3xzdbGaguxLsCYTWLWS+1xxm+gmPi5L4uRUzWzcpAEYLq+6fBN7ZJqSO
V+OnMA8OvFxzgT4RZ1ok1qjzKR312cfv+Yi7VX4U8zBMORnZYMooaxUgGNW5n5kBKBbmdCYI97fl
2b8HQSm8Gv38VTssUNWNZEvVA8O87OQjxacy+hePxZwrAhZ6ZRg2PVqPS3j4gVfsKz0uGOBJYkt6
eQbqSq0daDYMsYQH9/shkV9u6GrtBCu89sBHF5HMWwrNGl5Rw05daf1rQRMZaSppD3FJ+DIEgi5D
auTvehkZRTzjcl0QiCWjNM7RGb+QnFk00EW3cbtTLEHpMB5w55rQr3k1qxThMB+KJyD0dPtrID5F
MAz3irVNcxd1AMH/U7cCIj2ZJZ7Ms95wNfDFKtv9JlyKRDl8qk6YMr3XygWU7E4bOCZ8UWgyuNKO
+xKp4+pZCczFGAtqqxjpILeyQnVm5u6lb1coeQ/ivAmwdOUi0qQzoGDOUra0d5cjii88LhDNDFlc
Hvt4cQuzqE6ity2GZNL+yiQahrilmOM9zUJIirTdLShkurcvd/4gYSxOTjvumIIjfpxruYpwgHvg
a969zBW4IuLTbzw2aBmNS1q4ehz4Ew675KhdVjZL7F4A1xn0z/uC9TYi7x+tno8UIsocQGUA9ths
OoRhb85A87p+YrRryGsLn5pGmIxDGr0iVk1ZbadWL+6lRwvyNWXnyQUnrnMKCihZPA4K1j/N44g4
T2t9vTuVQKw2OnBfU14WLYq/jiYYdJl9Xs/mWvkhU0V87Sy+Tzr2G2FfEEGKvPDS5rpMlxokedAp
ab7gmzw/BARQSN62eqNC0wtHaS+KsPXvGIS+5PR6oGMbSb1JE+AhpY2YicXdtLmKzVGJUV+Kbob6
IImMNPHIUtdk06AZ0l3uiYPaWCOMSuBItYR8izb6+CIui+LDWlRSCzDwny3AKQs8B6nMZxoX07Ee
3jfTFLAn5gzX/pIkTroNjHECnWLN/pJ6zXAGhze18Dji8JTE0JF79FYH/JJ+OrB8GR6okk1xzMWh
Pa5gz77X7Ea84kY2JIpNYcYTsRgN+2/4I1awDfzsC7ivDkQ7J3yvVRFUl5l705mZiu08aEDb+gVw
MHclb4Pn+6F9ynrByqU/419UKK8CSToPITQ+m7m7uA9zTuN+mL8h7KYD2QEVHYmp29L7yhSZIZst
RD6OpVthqlWOqWy1Pil56lYqIpkzIwfqoNWLn0gKJwQbENU6vLL5f5DKJr+Ah0l97UyCpxLPaJPA
qzpnpdDfjioArnAiUaHEyuhJDRrMaPtIoVHLZDvl/JnZ0s61p06zGhnMqMvPYHqBPWakWJDzFeHs
apOqnYx1EQd2WJspqxxLlj3WPf/uMdHk1nn/PN76nWseIxlX07tzJHMrojonSaJdOfnT6mq9OXOK
3KGrw9FX/RzArREx9yy18RXuJpH1FzGxhPWcGPPzBkTrol6tGXlRsMvM9CkZw/t+3IGzgli/02Xj
pu9oz6XsCoVD6uxfDXkV2gk+Lnu2TijsuRVX00GTMDlZ2GlhUjUU7x5FEFcu9UPE1/47OK6N8fkJ
j6iIM2tP6gPlWUJkYKxi4sY23UeEmSa5g8bngc2Po/oODI5r+1ciysfChZKahMPjUjV7Pl03E5Q9
6gPXCsOiaEQmIS1wT9Bt7es8lJipuwVim9AFF5wA902zswu0gijvtweH/60/2UCsEnAuM7CpYkEc
uJ2Lj9HrAqbV5cuHJAJmW7KZ1ETH4J1ft+vmJ3wPcZUKidMJOeq8F+ZVugo8iKdyYQyFuv2/eFEO
CjRGYlDpgAEATznyNhckErmWEx++LQwZA+AupCfyLQieM4g8Ted6ne9k97VAwFOfzyKtVDI0GZSJ
BQkMAWdKU3lNKEWkMejXyNFtOiz7qnzFP6pUGfP7qO7+N99Vl04Uxr9pSXdWTZzvC78lAhY5eYxR
juvuS9VY8rkSQ3fr1cpm6QpA18qhuCGi4xh1ZxAZeBh2PGb6L8zmHdFU3wQAds2BksWcCNSubdI4
RryJ2F/sSqtt3nbFHV5Vo/lMtj+vP4AP7XS/0H7not8DwUHi8ugYqHPA26/YF0eLR1dhQyCR8Ka6
vvIbPydKrgb0eRlYuTcsPTbe2LjVSBkIEmnXfvCN3Hr40OgcYSUNupjY+7/JFU8ShTp3BKCD1aMX
btczFdkQBlioiAt3c16Sy101L/QbXjZQn+roYCt6zXis2vHAaZNOjLtAyfs5fVLoqr1sydnaoRBO
lMlHD3HMwI26LiIKk+AYnSn5VliyDn2rG08f59NbTEC7dRJY2ONeasJ749YetBQvQLE5mVHC2YpI
fQH1EBBS14PfPqPPz/8ixEHTkk++tyXT5UuTOBDkO735tREbFP1RssMlUz1XDfrqk15pVi5pFdOg
vNGmqF8CpUOmnLUlbNImEzYeXTpfYDODml7txoXN5KJzN69xilHbv2kVCrbXiY7TsogBVdGDY0h1
KFjJoRStuhhNyIh8m6PO7oNai++KtKLfb3Y7dFohethkT6/uKUqTTCWhgH4OmaYzcfpC9d3rI2cb
Wvhy26KUPsa2d+nJpURgoTWI8Z8sxCz5R8hcJPHYeAV7JZxkwbMxXDNbQVltEAAtOFaKfuU3dD4z
8fHCEQYgwLV0rXuBkZxD49QHZMyUIr18gImY+4wREQT+n4kzWyq2H6LHCDBVW0TmHyjzRZEy/SeM
ZDmrsBMH88JzaUsm8Hz0XBkHL7msQkBLAlmfzgghb1xh7YTxQSCm/zoQchToNLzvHt+Hufz4rGyw
ZkKiSwfJxDgoo4IRO59cdPB9BjwXr8C/FSdWIX0RakifrXxpB995VKR6qGOb166T9CWRk/+IjyZF
OCMFHBEPxUKp1pctxi7bqVl1rT6Did5tcql8UK2oKodtAOqt73FsrJg0DhY0E9VHWimmIrRtgemz
wgjDVLRajLfbLpOtWrqbNfR8dfCoTwzrqyP+F8e6jmLHHzxu5ukImCl0maf3UhVAberWZquDLcyq
1REVb/Cnk209/gpn7eo8hLD1CYsa6Leuaxaj/2PFWq6JwORFuKHSmHIMsmECeBBaV93MtOyUJYQ+
e3C6J7hGWrQ6tXRPvd+8eyaCJDV6lUdSzC32nLZk6eoSaICESTT3BVvWs1kII6wB0VwpAHvCed3S
44cabB0LUwJdKBYJz3H7wUC78Zhv/wFougTYyGAMp3fBQn+xgVyIb452OTWR4K1N7jGi/pZb6kal
KsEk5t7k6p/1PafTbrW5iszei8eNJh/a2vy8Jw9Ck1y6kLF6GbsuMtQBK2EnzQtwhjAs56Yt8+ge
dfbxURHj7+NKT0w8wqWmGYVEq6kVV87lGA98hBEuNu7bXEUhWwwQalzBTG4kRbECd6GNvgFXsejx
KlQE7c6eaaFiYGG1/MupJL/zB7FQkngdvDCozUVkNu12Io+kk/tcKnYFn/VXEcoaBA8qmla8xWdL
K7LborHXNtVVDSVANySJH3NNWXNsHIgP4VLQbcCQ+taLKW2Wl1iOFvPm6n74fdpG9DlYzJSbVGY0
esXeVKzZ0JDmk45yr9neS31EhegGy0aVOotAvCrH+5VQE2o+wPQM/2FdaCv8GZz2vnw7vhzS4b5w
QQPLYaVt+ubPmjbVtFPY6dN03YGwQY3h11XWwPULd8u88KLVeXROJnwSS+wqQjkxh8iZ7vCItvu5
660TNSnFxL1kTZ+fKD66bsNS8arO3AvMl5+Ja+f8YNXjrGeAn+96HZ+yt9vxOqiWuscOyUTFqEj0
TQBsVfmpeg7OhqcRjYLGALAvwtmUWWg+0XVFxnLZJ+pIFJfhenhCdGBIA/7vOZUguaScPYuEwqi4
SofPnp7PV4oEabinHUj3ASBr2WYujbckxfLX7FcDMmIjsfT+2BGiojoCVYY7dNdAS7VFxDGERa6w
EXYd09QqVQ2X9FKHU1D8B07tRcCmvekhdLWRpukwOBoOMOR9GaoYwxrOMXofmM03KgEBy942SMlW
NShJnieq1xVx7/CTuAZCmT8TLBy4e80+44aa5Blwlc+wmrv21VaFn/6vNu0sZ20rVkinTKQ9cdHt
8zlbPFEKCmqdZYHsTmhsnNGhbw+V3GTYfgA4uHjsreX8bWjWV8e2VWFaDayUjLyd2KT72CXLMsFO
cKWsO49DgyaBgVpx1Cfddl8Uh8C6zYdDOW9j6hyMaIVa1nsg9pcwf4Ta+oxGDRp0Z/WMCnDrz58x
MCaS6VONknm3pECj5qTUR3MQzv2hv3cCjRX0QAH2t4+U3FG8/d+5J828qJT2wMtVMvk9DBrkRVkq
zX57EKaqyZlniUeqCy615n8CjkJX2N70D3gxBh+P5sEXLty47XiNe9XK6MHeHvrBj3hGXRigQYq5
UwOBDC1xNOvEPuY3CdIElItWmCTTxDmGNNfLPl55rZqyhZ/zRqscvISqSa3lZd2AJWvPJM5L+6Xy
nXZRw1XvRXCAh0s8lAfEyaKd4RQ6EFZJTG0Yah0bpiBkTx9EqGcSfVwSGciMIoAdn+SGK+NyfCtR
wkfgFB00wC93jQiu6SLk+BUDvHa7hyO8zX5WZpo69XAEDZ1HeAL9N8tjcD3/YAkgT4bSsALn6Kl5
5CWXFVJ8iSzvkoQIVLuHX+iJuwPEj0L/iR7EcCG/4GhhFzlVyq6oZtxs4oRpm0Vq5Fc2g/bKa3q1
M9JfYKIRmf1lvosTLhMjD1MZ0FG3MigQrb+9995BPihfOZ+3mmYYUAGCR2ym8BUvoZMptNyZ8sml
eVafmI7M4XLDpHvhfy6r2FX1QA1He6sI2UcSf5YwQfUNMxxmvRs2pYTTPdnALELAeXwZXCjeB2z5
MONIvHA6wu33hqbExwibHAIXQyuUrvb+vVE21xmSS6KRsxABPnYodEzx7gHNJGMvk99dzXJXDDhH
bUlXkkzkUsDlx2sT6PzrWbt5B/JbJUpyqPOGEWSXFtNjrzHy1hapEW37H2efy7CCv6fl5Y7iulgo
YKdKNKyffMigG/vjVdHA86DDzs+2AnP0LiHsn/BjgHqEQfB9tTa1D18mgXUu2Bcj8oKnGvkBM9JN
OfrfvEhe0/CVe7vmF2+Uj92rPv1oL6JsQzGpcjHKuXq7mbmwOes5grCTan2cQHqbhie3k5gbDz5v
rPNJjif+YfhuME6hfBzHOR5C6ZH6cy0oxrCvR4YSVIudiSe4zA9aEVUngKENuGVHEhK5cG2uOJOG
10zrjf2rjCJtIh89AH0WQmXRMYOCOry5kykOtATLL9i7f/dRcIcUdHvQcqBiMalWKTIcYCM4Ydyo
Ne3a+4Vg5/cIu/usjCXTOLY49MOdEJDKztNqMk5AhLlQONA4G5c1EgVpsiof7vF3SGXAw1lePKxy
ezzCiAwbR3zA4oFMcven3Gr8mqZhFWSQNlT/qftPhmHbFHFt1et+ov13ubJ7kgepVYGfX59zWJJw
0JvWutHJFkhATRvYvUFziGDr7UBzhbyeMOJN78SpTYbCsMeKkxfSXe8AsOL/nE5EQqAhIZMCTSYD
RPDR3OQT0N4IRoZMLiZ6TIYiawOgiOkfwSmKOPDpErhga78gqCzpbhgrHpB1sCB+875RryjIxQUM
4zRKM5FSMxnOBzkazs6hV9BCVKJEfEz040KvhBmaW0nwvmezrC1GaP0P/xwM9xXcJaUSww8eEh5y
jPUJukQmfyDNpVjNHFe0fSBMzmI8Qgpt1hA9DjKkTrdHg6LHlLAMpsy7SytTPZrPUhpjtl3fLElt
LxkshQneYnZ5IBU5Wm67U5jI7+8FD4tbZDuKasCmZqk2TACGZ11iz6/4agFjygAwe+kCzScdGhzm
3y0N7gWpDABuqCCHRbyyQZDsjAP88Yh1Hazd7rSF/ANqmgmjqItuVMzvl4HaYc05z4U/h5b+GGCF
cuHJND5p8BttLBvza7v9qWuDYRa77nkJGtx8od3WzHDZJTpbkJPoiUVJAvHbBIn/fDjET7QVKn7z
g9gmFamtWtgetsyhFa2Vcc2CAt7rUR9Vo9MdJIfXB3nPNfUULICB1DRM131UtIfHHlJbZAoxCAgi
HiXVoIOGjBsnGI3SOdlWSI+8jsk0QQugVo3i+Jl6uzWMUCWfy2CTMdlB5gCls53PGhrhZOOQw6hB
PqB6kGKVZi0sFr+yIO8LZKw4y3SjgJwr0cmSqwRsQY6PRwguna4qZULSE0QpL9At8kN+RmVW0tQP
a1qOFBMZjkLFnT2k/BElFkXNgpJ7TbB2ChimMa+bjDPx5dxihXiTqFKWVmLJUjJd3OxVunDN08Xq
Yh40bqOwCHCtFgF7TYBLO//qOSEageTBfQMnY91IIsmJJ4eSwpDXXUSH8Thr8vioo6yQYB/JALl1
bIt9uhuchv2wQcIu09dWeS/KzvMcFuNZ2Qpj7PGPD+xacwYyxPZmWQxuHmc97dHtA19hRaLdbTqH
7g7gsDw/pI9m9G+tNadwUEiI+6cRobaX0TaIhsud1m8LHLm5rERGyIVYCanWLWN7eREmB0t6nNc4
pH7yuGVjU4t4mzSC+LgqBX2Lj52Er5P2McDWYXPuljFotyVOFpC5t5gcQuRvQxBhjVwJ3eMJxsRX
FsmIrSq6zh0iRePeYPTs8ZnMq5ANR+kakcme2U1SeIxXil8j10EicUTIdSn8HMGrLfLlS7XEec2L
xnH+YzsnmUH+Cf3gocfuEEm74XJCBy06kkbjTa71qc/iYg61Cg8woDZ++s3xsgH7/nsnReJCm8N/
Pt4b2d5CCgERxxjnuo81EvUPa5PPf8bc4Q6UXro30RQ4VqHGUMjmHKPHinwZVgqdEggm+8/LXfhj
uGqLqboS31fmqhq9OtUaxuZT4PW7MoZeEw6TACaoT1Ww+KuK4JKedFlJt+0sAC4JVODahGEabWsu
PIuaCS8PvTs4rP0ykr7QwZRvcFZLzHymeXq8ambSRKfn5EvuKhjqGcyqDZtfePOANfiycJ651dGS
XIxhocl/TN47kEf/+DJoHPiU07x+9Lv4aU5opgpvzs/pjnR4n0HoR3KYIy9tHn3Yk05TAEKZzrr9
Rb9rvhxiZkJC1rIJFOCVJKBxM/umMA1FxSCx+rDTsL4segWs8RTsWtx+eJYSUGbz6edCVTjxdAtC
4Cya4r1OQmyFBA1NCdiDbD3etbsb22m9sIjQ/TVlRveykScCp7dQFRtyZmCtnyO5XEYqFvumMOmu
CZx4wTCwTdbAwfGQ+zO45v/Jb0y41RnHkoPkizmhoeuYEU5xKrpH7spTvFjeYzhnfb2HwTXmzGyv
Mq4scLLsBdLoXPR873Td0NdL37LGUD/GwSGL8SvOx24Ht7UEobQoYNxWuQ1ClB/OoKBc2DSpDusq
h6mE4pIB9lOYf1XWRHZcBdNXwsf++c2LdM3v1268P5CxsDo9xs7f31IBBAQQ8uydhqGU/Ouhvn62
TsiXURsqj3exCoShKR2Uru4gdvR63DGTOQuOJq2dOHR+lhDnOcD18Bs1u+FAOeybS78pTJNFaiTD
A5pEMkBjCcOcBukaqKFWFJaU4IFGOzGwWWr5nDZsrLSKoXC1zomfLYNHDCl6PjYr78Bku7aVt7sN
0Si67aOpNFu/9bEidFCxXCVvJnDB0gcMxyfZIuKTp0qmk4EK6rYVEdFZ6UoBsU6dJTBCGuNUrbzF
2YLuhFkXvVPTmQvB8U68CNUtB2FbplZZfO6Lj3M/Gs8uGvdekvFWcgklMBuf215xU9hdWDdGfNH0
YdzEp1fIjnqS4LGH9h8TDqeiv3nuut0quWDVFt5PscpAisxTAhQL9QMpWmpjZvCxkUUNBOVWP8lg
0++PaKio8a3OBxpx8iTu+GlSFSfEuy6jlsGnfGA4/RoGprNL5JUDKSQ5WvZxl6aQ/4uQeHEdjnJi
9667dzMZCEAH7W9x8BhTm4g8iNQRzqZhZPlqz0ZR53ci/KgOVZ81usv31ELnoFOzA76aFmePo+8S
2Im/SXoQdAPvC6t5btHogHtavwfb74EeXKsjhSPTM/7bamfy2XErIMGfOje60hdStgLXIZZXF2fa
+4gGpvm2NmsRKS+41GdgHSlT+G6CfRKPNIVvmqYf0oZv1RqkjkxArw6Ehd64LQiPi4Km8PhMI0BG
5+kvt4BLOAq7pFPLK+Htj8O476Yq9bqLuXxMEfpF0GTt0Zmsd3hqd4mYM/RspME4o+I4u6lHuFkR
KW3GJZgzNM8CZsDN6TANxuYr1aQLf1UEu31TTX5WHR8gck5ion2/IkYFssMK9rS97nFBzmZm7AT1
30skJiWZN1oyN7F4aeJN44nu29O5DBTNzhilPYK7V/A1n+gpIWh+IuVpaZm84IWemLOEzGtYExa5
sQWjoflpwBIckm19VETmCVYdjoO409fJjST1B8soo197ghf3/NDxzcRsMrgyyYBh7SYBr4h+WpfA
8S5yDaEu+v+0SGOcbq7xcLjBVupvDCBc808uTIoYPjJiGFABLImYnabWTn7t1Ys4BqftXwP9+RaW
/bWNM+1lUFeIMv9fruYE8y76cQqXE9cg+CfL8vHsLM0a/jBVHowOyFU9bLPj/u6HeYK1XGkjC7Qz
holPz6yV2g5hcw/sSFw5TOsRpZmD8mjm+fuWC5+pYgPoFvVtv2CtuSzAMvqFKtSbyIAQf8MRyXqX
gyEelAmbOQVHGC8OGBFi2Gf/DVlN+gNXD5rJV/bD8G41YIB2sPkAQJV27uuuYBzgboJC68zD/zR4
dSi5vC+Anqo4vGvx8Ywz8enZ4qTOAAGlLp6Z1i7An4ZAAtUeVMOF8lUc3PoICJ/yXPcBwLMFu9E3
Z08h2Mx01wSQiyob7+cs9Ml0KaSOh9SKi/BXqHJ8Q9DouufB0O9AP5jpcK/3TA946HhOy34aKdP/
+3zbGVAT9+cEGIUUwpXWnfEmnuXpZw6lX+MZkpeAaEYls6EbBxRedrZIPR0DFnvq3NOaCr2vFD1d
gkJ8vMyaXRy8RVbJnHdfSxktkYA1a/bSDVAGD4FRY99XaH8w84hXgcFdXYm7bU6N8qrDX3QUAkrQ
rUovPJXaHQeyBgkjdBGkxwa6A/rmlq2s2rybKBUPa1vYObeU5oMcTYYj4hNb+8jHQgx5H5IRf/Qu
lqB1+mSv+rVXODnkUNx4e8lRmpMw35GgqUBi9rLsgd6VeAQX8MaEyPWZsGR7lo4beCH71vdcZrFw
6N+fCk8e8yMaG95Vzjs7fQyl6EEktPpij1kSNIK4eGNwwEHy+mH1dU0mhpbxvzGrmvtVwhmUiV/W
jg3eU1f0crUYekftFMZR8qn31dCdtKGX9fgq3dJHtsLRtqxGTiRDwoPXeJyLXPCwFXh+/e0hLIV7
/6Y/RTbYuY7MydyFsDB5YO9Xu1PLSK/L/GxINiK11B2NxUEZSImq8rUEbDhsn92ortl+n53/5gBg
Dmogtf9wGRI+6fyqEapTy80k4VSgCVjcaeX6WPoLSURnd8kS6ZBoprx15Mcws8gg+ubEYs8oXIoD
bea3l5rWlml7j3DKE61A7UcVY3eucR3+pBnUbAtcARBxNCUud/ffAZLKXOzdCDc9i3F9T8Y7BTIF
rSf55KqkJpM5OnQMyyqRu+axttYHu7bEpNDPLFX5kMxpGoZBn1zgNRH6v54WYGB2fchAEnl/Nk9I
2Mx09zdilGr4VdEUvGr6k3dFqNCRtcP8rFv/Zsiycgp0hHFjhDC9noAGhb7td6tDgXxAFy1hBNvE
EUAITRuWG1M46WuJGOpEjM7fk9HKaJX6iqTgqhteVjCeWnX7omRAcacaOBNczzKJ6D6mIoI+2uQh
ezE+NQDH8OLRsrZCwyfDI8ZvG9kmvIro6oZMQyj0+Xe+0Qik5rGwoBxEn1GJo81nH2VnbOJuf8/Y
TSL52/Kv2z7uykJQrlahRPo1Zc6ykPog991YuKhtIUhN1ZGhOYtoi6w8/bSKYnohjSfL7SRHMhX1
01iuIjNf1gkEP2Js9JUmtXcB6ZZ14iipWdjWN/uL3Sr7Ra6nGX4jH4J6KvJZTV3k/WDmLepY2Knj
HnjC1V2dVm3UCGWm00v5Zzh0/IzqIJvBGMqDSEXlNw2g3RXOaRTjSOOVfVY+c/0ujaLlJyJAqVgx
HlfpLh6DkHEiUr14zHDewhipfNV5ZFpsWI69blaWg/KPRZX+UXi95v+Bxn79ZNWrE9eoltoUPcWJ
q53XnGgE2UFO68T1zjvbB8dcwM8x4KsbWkwgWbIq2Kowqwb8udhdSPi+eH3jya42kY019vzKX+lZ
bRJwe/R2MdfyWdMbH6IU9rIHTOQVsYjJtq2G4K8b9qBfnGxC+Uy9rfGDqD8k6jl0rhM7koGQkW9d
b62tW9e2lx+yZesr7zGm30p1/bOun705iO5faOUTyPGDDwffUz/l3eeQGd5EArqXrPCJQBniveSM
A378mPY8yUlPaIfzyJB4IiFINicezEAmsqHLs8ZXB73W4yyNxy7KDZpCRxcUaoB+aj9YTVLOh66u
WPzfyAXN+UNqAvQ/z4JTxcNTbD/VeUombkbAVn6H33QUJTGN7K519+MXuWqcmPQYBvtI+S4QMe3J
ptmQu8X86HoYI4YdtDC69yOddpUHgYIBppMCwigcDNb4vJmMk+oOPzNoz7RizumNBK5oXYyhyCyE
DSju8JnLV6lSYp40YlVXLssIY9rSnCA9fnAe29PcNGvFUoBTy5RpgCWEXkiOeF0TCnTidXsUzuyc
d1Cgsv1mUok6F2oWDKA9dMejAADcmTaMwuxyI0XNOXs8QbkLuxvbOliSbsuPiExXKreYlDZyUvGQ
4iI00qvbb0yMO9akm2agR/63/5uBQRi68fcnE/5XSt1Dy2fv7KaSzyq3AgKUVAXh/axxyEUpJGHX
JoRpZRoyWeKHFWEoQPWIRsO7SpZwrKSXuAUO37dMeDleajIzRTmLzHLSOel8mPMuxB083hn7vUIJ
VnMF+EQDOYL27H8crxKNVIg4u96e1EESgCMg6K2R6pvW3TbPcULJfrIWFryFqfcsuEIK863ahcO3
9jYls7gAevWyPVyRdBLmMvPYr0PWf73nPdWV5mqwPBORfN2PMzPUL+5Eb+9dPJVvin4kuogyJMNv
+jIU+ujhQzecU0Eu4zEo2pSLYlRaRovWEmeNTihQkFmbBKZHKCHJHE+04Y4mAI3hhc1lBXtUNxD3
9Uu1g9bHDPyIZsjuZ7+k9UETADr2qOZTWbGv4KE16aZmomgwEUM1lnRudfJrmfgRIsEqzWbOpasv
aAt/qTHHwMcqPpeQ5T0u2bNcaePgkWk1ByIp7ZuGkJ1NEb4ZB7tm8NSrBRj8DYqTJoiQJZ1oZ0bo
vS9fp8e6Chx2kXix2GWPupa9n4vwP7ynFJSZFR82sd/kP+UH0HYvzkrQBNzdouBItoLTajCAHIln
fnqN/MlEN24dyhg2M+XoI6XxPSRmIYkj1bTmczakZwDiYMo83vE/S3WLUWeeGv0gUTuE56tIb39v
l2UgxcLZw0WK4ZRLaWFkg1UBK6AZpM/CUtmEVYRdT1J2pO75XHD3KUhmjM4A8XbIjvvsa5ZrjBDM
J6ReJHm8V/2axI2fAjP7RlrxsA8gm6sh8eD7iuYVgRjMMdxbyej49ajunxf9YRTVgvF8xPPJo/cm
VT21bnG1f9YY1XXps7ztQaiqytVpa5bf8TjEeBFVVBIvgvTVd7BVdM3I9Au9linXhv40YydT5A8A
uIHGi8wz1frJFbuO4IBm6ux0cRyaR4FYVdamaz7etMgshJLOifhROctfjXeB1eksCaF32cqspdM0
XQaiD0GeDOaXKgTm74+MRvMTrVSnSxY6Z6F4zsc6m0R2qxd+uRsrXSvTBUjYg2gkpiPCyYdZYz5J
+ak1Jfmiot4kAqESQZT/PrEnc03ffbV3Vyn+7oHBpk8KtBk7nqa4YBFYx/aPihF9WOYYvoVMAa46
p6LWaz72NZWznIlxsMdzZzkPnOj4bzXrIVoOLeQVRAYtc1/XL1zFcK2VKT3Qj/zboMdjZTJsRqCy
d/VgtW/yWqxyCZkr06NGIK4tKWmtawcGwskFFOPTJSCjAj2a2lOsI4lQYbUXWt0uwDTbGld/xdBb
6smrQfYRPATIEW19wkXoxFDIFx9Yb43c10boV7d2fbdtZ+Z8AE/JB5gGBrg3iHfyvEqc92IO8P6h
NMTHsWYEZ9VNJaLluvASfWOwqSDjujs21Rp5KJ4g7S0qpfBUtO/5JOU/5nC0LvK0kNWPB3au8CF4
MYxR9Zc++pJRDS9zZ/UCNAubRBdClpxR7k+cackqC4MSXokpLmDYYxzabAsay4C2+TLqe0myZk3a
BDDSPcUWdV75/zcrjlkSJNFLWUGCBPmgPZ2aoEjvLJN37yDUFV9WZLZuQ4lEPPedYK1T7+8QmD/L
Tj4cbuGeP/9XhL4Zlh12QL5KKi8lMXmpC6WE5Kb2ugkI+CVse6ltscbcrMf8HOGo+FqVnmjapO2+
/efDRxcR94F+WEughFDjBbo8nwDOSSYLRpW6HbTHZoSmVLn1bSifh7CU6pfHU7SMzHfh+q/zFQn0
fGetcKikQ2ieES3LMh60xN9XTiwYQ8BiEptsgkIVym5uKbXdJsvncWTjUrHKLkq2uVHWQgDMzMWR
3iFH2ct4m9hwzDV2ESaxr+adAIVV4Hj3gcJ3zK+BFZ8lJ7HEJK0xZVeo/lxsMooF65xOUUuVuOcM
hrLBm5CiqDPju8XSsunlPW57nB/BAa514E5T1jGiXdAXuccwvUCcCR2A/nO4dBRAwnxyIPTlk6jA
uTkSK5lisY83T68a+M66SHnA569THVgp+UwF5GMaxspiW5ANpNYIUSFXJwoSihc0aVOxYK6QV85F
UfJTMAgJOWGBvJlplJZoCbbleqDLwnAoMnSpK4R3gmeJ28EhmESznRHleTcrHqkyngBUMqXJMeL9
w3nt6Y3OFs06zA06B6YMz2eiMgSjKJgiJtNBbPXQlp7js7wcDlZdBIFkHB+mfCdwuCbOuJZ8qoYm
1FQgaGwytAeSP4QLLIvCTrfyOG4pWfuYpqnFAWV7RZ520c13sDSRVH24BysQRUUEWa7Gxt3pjjtA
81+dPpE1OLRbYOU5F7Mhzz5R0pU3I08v3auIzfQKM4+QjR0itg8G7q5i+JRBcR4Y5t73OHotLjLV
g8+4bgB3YmQswWBG51VYgCAtOTvLgRXGTucJdfpQC4vLQ6hFPFvEt6fv4szBwF6LIX2iIkEvyE24
mPa+MiELWI0srbrFKwh7r9jehHlqq2unc+DK9xMTRUfkaQUlFzDDiy1RY2pH1omT8lrheYnMN1tO
OKNobbfMxnoaQiVbTfI1zEvcjImNiTO8SqiBvmVUbA7WhOiNaB77hfo0PrFbL8PT+ofhwIrkvt3d
ITrtcK2GCkA9pMR1TAS4HcE3TzSDaKl66OH02HsCaK18WAl9j1kJ9AxJkZF8R3plODHZdRCTBCxI
noBdvXiQU6b0MzkqIw5MbX5x4CnCjovvB1E/8/YE4EuoEkdivMg4ayAkkmyPDzqlrGhhUEzSezdd
BcJd+m7IPRGFlhgmoKf/8BCYBJj5cDoV6T/mdrU1rLL+FzB3/i4UsvJAns4OuDXY7Cux0uRmhYMB
jmNR/d1k7B71jPnxWZcHn8EQmw1BCEtQdWuXCkfw1FxpniGiIedbLpQPr8OgnC+uFVIOBwFRewFo
2DUK/4gXMF1hrsUzF1yDCpxEsmcIgzo8WwhDcwgMIWrrAge9YX3no+/JHMCbPftVTWhy2LxpZJV9
zouqNPmSW/v4vHhYF0E8ezNrUastqKbxPGZk6ly1Lk3vytsAQRtub+z0d1Bcwsn8IPOgZOPdKl6v
0jIqQzcE0ZSLmbJy4lHiYhZ6svUFVazmvw6IUdYHsJfIk+RXywB74CnVSYwOmXrjPHhEWvTJvdIF
hXveSWUP8TSp1rSWu1fhPZ5iAy6ZHeooSJN6W7yQe9GrJu0MMW+7k2wHawQxdXQmoJtmQbtxabty
zLYGtRnlU+daooDZwp9m1m1BxtBT6I7h8G9KJ+UQf6GHwnUzuM03QZwKR6BGl9xIvUQ45R7o9MCU
jnVjpzUmz5QrxrHXqpT5CdKyBwB1DbJBKtjUUSwvy6blUCVAD/hmsqzqNaNqdZ+e2W6JYH563aHX
QA1GpeYeG4QlT4eRUhURSnYhPkVHjfVITKI8zOBEW88DgwpA8RDEkh8OS+cTMKB+FI+AKvcQBPRJ
y7vaeZhGYqTRDziKAALDBWeErSwMRNZOjsuGB8X78tsJ8dyzovQkyy3lV53hSqoWtf8ynBJD/1PH
b/cxIjKjtFKaHinhcHIzUcH62uy8wD2P8/QVREdBQZ+IKC+MHOokSNS7pvBFw3TtO5pewuvYvtBa
RwOiM8OWkeQhP8xuC8MK0Kj2TsYQQOxyR1zUkoIEB5u3RrFLjYUsfh+NftthGDchp7tDp2q/M8oj
SPTm8/M2qD31tZ5bHv975QnFeyEIk23NEfuetIa8Zb69StmP36QTXa/tMBFJ4taOj1GQn3Ze61FV
eRyxIdtV/UqpYkTi4eaFtqamUMegmmu+ZL9hyVAs7GLl7GUQxZKTdzrSRrYtipdKpeEG1fpzzuIR
ZOvgoAaAGQh04qKLViIPZ+yi1c5eQ1XjD61UEpz2n46tP6aUhZFo4fWx+tGOONjcw/uzSl82JRZI
qnCg/QLVnDHWBwjH1bKYefgmhAKMxSjgbYgEtlf9bw4oiRJnMZFHph37ePMWYaf+JuGnRzUmUkuZ
+QBlktuwwER9/dllHzSOA9H+xDv3rsCP44HLI+b4meAy+0epvHP+uPjPmPgDU6viNKGUrZ8L54iO
YtSWMtU8LbsirJcYcXPWXQ6ADQ/9gBXQV2X7/pWTarkRxJAIt6puhDg7Fg/Tyu/Ck5zVoNuKn9LN
ASLMkNc4ciml04YlJ0+1S+OicaVDzV/KbZ01+d8xKb4IxmFHLOixm/lvXRn4gPG9ERG4Go0f21gv
7BmG52PHE+VlH1DPM690W5p42DC828Vjsm8F4X39kjjinVK1SfNhJHsNslZS9Y4jiXnuZsQeOO9M
Wq72p33aPL9UpA7cqqrA5Jvx5JvZj0TbTHTzTU7Dw9GvwwgkvJZ5ULS8PzcJN/xXaZUW5McEQZis
vc4tUv2msIu3009Z1mgDlZrUrrHe9up7hRDuNhYC8SWPmsHOq+FJcrffnZD2mGdkP1UIYdVeXbVn
+oSSP//39p6tG+eUd+ZMrNeQZC7yBrlGSq8LByTMhHDPnxNbHXpviKN29dPA30zVGYH8N5KKd7Ff
vfLz4HhBPGz3BZyTXVfHfzxl3zxo6QIlgWWMgfY/L+Ti491hpc7W78wvdSxvmQhuDTdeyzqHJW2b
H8zQ21k9TtarZ+qAQokjI0xj5DwUr8wffjz1aZB6HcBLtaCRBypMG16y6j5NeTMxmdrMZaZqd+Ut
8hqI3zSIApnA9+asAzrsKRE1xb3pN/hNOsrLYOfSx5jiNljEXT6w6IWTW1k8tnjo/QJnxMmLgq56
QUZwapi7gB3EY0zIhU762HEM5MYGSF5V9nHFRNSgnU9uFyt6VmGha3a+RyMrfKUJWJEWzSxCmMT+
EJP5XwqqUNjw+w+OnrZqziSTMnOuNYi7FGTDx/89IA0JZxVq6Fbe1v7iBGKJT+mFg6J+r3TFTB/n
bdNK9sxQU3jujoP4Zr1ljBvJ+WsEtlN49H/z3C5FlQ1wGzuAEmSUMTDxj/j0aB+IsdY00uMhbuF8
aAl7lN5pUPAMQCHOcDLeQgN4yyv1B9nvt9c3YsUezN+UfF5y5AYNofqbu8r8yWc+USqrwc22wFvg
8fW+LKN/rWNNk0G3OpcLPf/M72CT4HzeywBs4c410jDyvjDnrf/RXpiFNfen42AgiPOMOmkEar2v
55eZxC8F+RLy95W4NgMYN9NgXYLgcx1mV7kqLQD+0elflmGt7OAGTmyjVt40yTa6uhg8mVG9X8bO
59wIUOjtcBjX5pm42vxIgkdYfinWdFytSUUxu4rxsWGol2LGJQlJlVENQ6+MOzHYWBTMDbI9/mLD
QWx1ZLyhQCRLyQMcZyE2YH4h8Q9iYFbJw5sjg5xSM8pGY8RTNIGBloJYVaRIHcXYQz/LhUAUDNGH
/Avh067vZw59dZHVfTBVDS+TV11dbVsM2BtQnHLiquDx/UZaoQt9hKVC9K2WcBeJttOUzfCkZBJh
u7s/WwiVLP/3H+ATTocUFKjNY8Oov64v+9sBBkSwftp4HmoPFHzjD8QSN/Shd0VlY0UTj0bbm8Bd
MB/GTJfkiwVwVv9Y3Q1K+8WV3Uv7uEYf9A67kP1daMaiMvRVn+e8aeMRO/4ExSSEUevntMVPew2x
Z5eVTSLKg+32lrVdxQF0QoxSJu6LUguttWRNOXETumPjOCypsm2Ls9NH0UfUt5a7LQ9B5SS5f6B2
Q87YlqEZQ54vhL4ieI4nhrsk0Q6L8QSdmTm+1DfVuuZ7q/PDWYF1AeWhvCHZXc6Od9q6DJmyJbOG
HG55tNm9m9tp4qXgRWtc/R3/yNrwQ2ibqA9Lf9vwdxwqv33DtkYXhlY6/oIvShUbQ0HwiCp2pq/6
KXYXga9yA1hvalv6IcpuXqd6HqXo1fVD2Ww4MkHmkJfT2Y1NEWlDCnHXITrhvKtFDBVN0aJYYnjF
vGv58/suFPTmzu4LrAvONVyAX3p+BvFE8SPAJNgU1wILgyTu2/ED9qZPeOjQSKB0vsElWPj7vOQ0
N/g9nqmtt2CvcEsSDv6OrhBu28RqmujeallySznkM6Gj47i1zO6ElA32eaz2LtrLKuTjT3ps0FXw
Evr7hknzeZPwQSmXEAboPFrjqyJzSVuH4z3zKThHrewxrTyRyGvJQlCEBo3L5Uk91kF9OEcoBplT
wTBdpY4LEGUWz6C31YqZXAkdXCU2qzjFOqA73W0JCyZwG5k5YY2UC/FPPkFAx79WB6z1ydpgm2fu
L5CkmdmytnuCKYW98aKn/MuTdrIcB6OLpVmc7+BJSxbmSCiGU+B9LydEN+AnaViIp+TpQ669uL7v
Lq1lHFcgqUIbuYqPf0oYZ4ailL2j6FgB+jMjaaPwXzmUd+o/3BOt+QdxA21/S6F4MfGhTdzWepVf
kmL1u+1ngfmCLTNoKvj4GmuAcNgKFXGfMft99p3u1C1maqjya8Ug7S2Lu3WD7N9pnY+TSO03t2NI
8EBdIx8GUnxt0/14Tr+eGwuEV7vCLim31A8Giz+WyJNZaxCMs/oIk8wsYgDNSkSCbiGKd4S3tT4/
z14KZzPWfAmtLjxtQbJFGc0J2J1GE+sI7kQnK/D5szjS89o4l+olx2danQfo5zq9lMRmx/QdxI45
+uxpUJkdVC6R9LmjIC5IiVc9j/ajQlBgo0kI/2eaByMr22I73MxNl3FPv4ZIJcxEDAL1FEzGeJhc
IJxwM9Cl4BKY2Rgm33DLoAU4Z47pHiAP8W+06mtV2lqHo4lxIP1o2M8ACXi9DX5oYV4ey6HLgvQu
g5AfsBuYG+RyQN5yJ4xRUXUavBExkxT1QDwWxTL9Om10MYJ6xHpbEi6iCypgengekxCfqcRHuygm
sew608APfJamkI2/xYAV5FAfbIFpWQCEZ2FP7cWTc592PtbBVtI1Y9AK+5o5qqB6UCPq464tc8yU
HfULz7FVWU8U9Ra315Ik2FcYe/CgT0sVV/13NzgMzgj5u6FqAtqF6vd0P8QWa3aIAPko/EdqVgab
0Ld06UBa1v+Kh0mzZ0w0vEn9hL4eKxxZUWvGl+UVUVtovDrUyxeYEFzGBUC3j55nEI7Put/5zhkE
U8s7OuffHtjKgVHmRl09bSovhM4t/LBtA7tqGpQMogks74P1T7Mjs4/jcRFJRM2vNgvmrEa1bvxG
+mvk3iw1C0yFUsKuApu0iweoI6jhC+BwCeyBBg0dAQE89F3QOyP6nak4sSy0GLUPxtkWAqa4JaqY
3WG7d4isI2WAYn3MO0HW6RmJ48Xt6dHvBvpsb9eyCXn+wCa7wSnjXZ5VjGvb4QHbR0Z1bEvubgMw
6a+QLI37d3KwB59wG9+FSSsTtkrlbASD9KDt6sMaYsgC/QBTNxmjyQcsmJ2I+NzVitv8pwUPIxPL
kVT5nORxrjeRzRS/NKbYgWMTIPrdwW19arRbmX7dAQSyUM701R60T7nSKKBfPOlI/QIJ1pwf+A/e
SjBOrrkkKxRBLgqUQi9l2ezBQuoeOCER6366/vejBs4lG746mGok4QmVhs4HU9Fm86T1Zj9j0F/8
83GRgVE0/ylcZJI8FFzIkgtTBEi4iV/JnqPDmjoUYNnhjYtqgwDPDFzV2JGEtXBMPiacl/gqC+3e
qmLGCXSJEtM3JL3VD6bskmT3p8hBBy+2+gwQcNHR2V4Ep8SE9+rBuj5ZJtkQO7SdRYlxY5ejEUpU
J1iy83iUFww4Eu7QprKhghkFwbkZ+N+sXdI3bejL6OgkzCILDun6vAkoNr9h+5ZS/BnRnYHAZ5n5
A8hDYRLQsCJc725wQmYRdQzcN6Vh+COYI31Lh7+f3r4TxbFuPk063wSXyNYWlwavk632d4Qw8NJR
M9amsuFvlNJHkV1Vhg+FjarAdwtMq4BaHhZu/OJY0PJymbXinYcXlHeZXBrOOxXyWtVo1wf+FQ02
aY/kxyT3ta4rO2S26UT5/rh1yXt4mTHd/i/AAJR6YeqWM8xw6N/3ogvYzO73DhwyhvAA3dadeEjm
rpa+Y0261bD/s/oEQFxqXjisjkIDNsHphOhW5m18Rh7KTEw2XzsXIfFrUkAU+cKwVwIkdkzRLNgD
rPKj057Xx0a6YCEzbTfsKVCnrsRSnFIZk+Qqur56B23eyFGiERk5iOOx/kj1Jvbl+dfifJaQUzxd
myu6I0QG7KXmUTfyGeqzkUq5fqOxU+eg2rHZRjJ0zAoo7eokOe4bVAeOY2Du6uvCKMTISJ7TREbF
x0IdpAe0BepZQ+sL4w4bSwtt1p2faCi1ZHdFtaauSQ2un9rIQgaJ0YLYpprN0xQxy8SyHhf5f/wf
FKsmCfS5s8GWyypoHVz3v/hQV15rL161Tx625CY0JDwjotxFHrmzBcjKFu7puGC6VGJ9rDqEPrXt
wugRp0FJuJCKYm5PssKt6sIHPhn3vF3fUwbvc5tJWXufSo16QiGem4aJ2CuWEFKFec2oIfJaZvWz
KvcQI8VG8MKoRwhz0/RQ1Q4qLxH282CVwtTLF23T8CzigbqozjU1xYT2ZcCYyr51wF+OjOMfpDxS
J9W5CJY/wGhVXCGcfW8+x1N/EfySiDrJ2cx+RPYLBEHZ/5HEcRskZqgkp6zuGJgQERWQhGtx6mJE
o1H7Oj+uJiDMXmuhgLOkSnRh7H036DTaOkWcPDoGCTjcLGx5t6jtDd1fliJpKTnmL/gQCK9zzJhk
jnfPeii29ngblhiPz4dEDbjXUyHIgUYcBDhyVJNGQQk1t2G44Qia2SrsqgEeJjuafcmSifdRBiqz
lmmzWkZmFmgCscsDZHTsOxZwiofnc405tD2dJIzEgEoo2bQqhq0g3UkJzivLJnQaiTSOGbjl7jYr
W4ZyMWRB3AdjKyKbUP2NFrTLNsJxZoOlqJxxW1PD73V1iwudzxCOugAbMdnuFtLPEAPIBgrUF+PP
GwFMGBQCXI6EULRjk2sNlPiWR/NUF8SJ9i1nYjWe/Ef1tdUuzjN8R3hjwl1SvG4jaLeNqKYzjAdI
aQa7jIBin1D6QdCwXaOqcW5YATICat7Pxkjg08XKNh15cN1Ocy2FjeZC6X+W8TsHLPr/Irixdc8u
ozVOQnF2BNQnYUm8urN824HAUet2RWRqr3q/LztGDD7qCRn97/anEjyz688Zj4LaXbuJZm67534X
ZXrMldi73whpyhEwdlsyyNFAiGaoGbsXr9k1oWZIYrMP3TSzoykgC3nd5q46RfvA34P3hkXiGQql
HqhenbCXEbu7gGCPFIvHmULBsV+DHdxKCocIvu/NPP61qhnANL2GHsXRieXhwAPySWaU+Oj2mT7F
h3vIZeZtydy/vpq+OBKDN+rSaieB5BfDU8c1YCBApvYHVHXpjLcX9DrsWdJo8XTx4/PD25Z5ctCS
Gx4hm89ZgeWmZXc2pLGT3VGHIAYs4fRTPANErf9NmfIUAIt1COMBynDtd0q1zXn3pBxTSaPkw2t3
lsGbxS8kK8NXr/zb7c27h6DTmV9huB//A5l5EDkvOCKOzFkETSZ9sGE0FAmCjAq/K6h6rkxoI222
Axs15rD0PvnmFPGPMKey1uevcyxQgGDos0r391AdajEG0lxwepNc6AY/G7MpLfDW0JIsSHEUUn7o
eOxwmY+64doNGVL0Nkx9hRbS7db55f/vO4ltMaZDz0Ghm8MYX+waI5zVHqzb5TXQMv493qmcOjZz
MNYsKSB6p4nK9X8var/boIP7ADi6m1ZyBSQtUnZA01Li6HZ1rEv9uDTrHEkM8isAQgKWKKm8qdNC
kZVhXulg+csFSBQpE8z9KzwUErNpFU0IMBtOpIc3GdovKmMkLUpb7Kevq+lgU+5T9QxyBzVbILZQ
bx7AzOy1aFn4O4kfF1/H3/a55/2qO+1GIpisvv1B8errr9JHDaEB6YnjXyrcCCVX1X4alv8R/3g2
JxNglf4BPkZ+TTglM0x7xwgSDfDvCFr4OUK6ajq9fyfnU6RDVlM2FUy3nLYsNNGFI6//XCZw0d3e
1p/5t6SAR6aEdshAoZC4/KePAt3HIhviNCGxsaMNNwdOrJ7ySFHIe6+pgHQUWF1yW01aerUNynok
Pz3yxaKkCAFk/yz/N25taA1MdWbunxyoUdslO93lBuJiDFPZfDuFLVndp5ZNYGF2lWPJ1ZTMWKiQ
24zcH0s87LJnR4GX0XIZgaD98HU22cNVXmi8C3DCtJfVjIyx8WvF9fD3Z9k03qSF78XYPn57EBJw
PC/VVUDcxCgl4k0lyFx/BaHfbsZmaRIzLInMDI1AjPGUzCm7lukgL3sZrffuog68+XyuU/jlVnew
lZpDjOOuOB5pq+LkbHdMYgTGeR3ELPFhnWMSEltj0ow/eVulCOTu3ZxS4MHiDYJzUYb9e6KN91Ib
j/PQgIggCUfkyB3F2UpZJEIvtnbbwl35lHGNYfWlfaa2NN4RZFpaZcYTpsKaKxcmMIAvKADD/kpF
y80+dtSQwE5nHmKuvhrut3zbdpu94ooNiEll77Mr53x5GS2jKYWjGt2f8bynaWsus4B6icqlTrzP
vvbCPobec7+wzSLr1HU6X2q2UbjAJy8gqO4KEdVPU1ShjGLRFUM7P0flh6hS4f5R3H8+zFCXfhlw
P54A2CiljKO/rbCXpz34LM0DnZQQ7g070q+0Y3SgHn/LDppD98g1nUIKcSBacQoH2we/kVNhQIfV
d1TbUJ5ptmO8zly2Pd3LHO7iZUSgl+O7GUdVAwWLqQCm56zIvHUPv4d8kDSwlmUq85yHbqLeYFEt
XIfxWOzO29BPhPHW+W01N1Jz0X/sALIzAIEGfTVWvFv6uEPayCl1oTVd6FxzLaxEcLhfyt6YP8oe
mbo8lQpDbLDB05oVgKE5MH12GPhLrbxXyZ5+ltnmjyUmnYIr2gV8zl6JNLJuYn/kuByAN6QxapTE
YWxWFMfSF/9DBJbnE8RUrpxheJq91RQd5bvxFccRU6jjUoYU//rA0rX+IE3nk/rXyvZCsN4sKcWg
VHzN69gPcQNXCt0AnLWP7LtoYGbVIwTu8KvUy8AIxVCegF/Gy59YvWd0LQOl3khp/kjgMrmWvdhn
bWgfYoLk+UnbpLfLMklRETthBqPmJQqywXUj8TbWju+54dgbPwqsfpEIVDn9orQ9tYv/q43q331P
fjZDZNaYAnI3HiUnA/ksMmuHlcb5M4QB7igHULSPd/98vksFCj837/5vGlxs4KZ3rRIYkdAQvuMd
rr48uLY37mJEVGD5wTNrBlNjZW2Qc/lfjb7AL6hdjnWRJW7x0aE1o6o24biba/SXs6LitUep7wQl
nENmeY+uOVpGwyhaExdxVEno2iVPkjjFUHlqcSHstfRmN77JX/Ja2Lr8YbGgXm2FHt7gs+qJSMEp
Y25zrgYKGn6RWmvDf9A9I786iZ5yIoFGThz6jzN0TBOxZBigsQH+4nVwHdF2Ltf2sUGc2QNGWjlm
DRqszUE1c+nv0KavAcb6xXjpFL8gQND/HgZjPfg/MDDG2yvbMMig6hK+yu3GCRpcrHwgEBi9YrZF
O4sR2Fk9MuSfg1A+UEjd9VCh0C1mIY2qPhyVOTSrzNNciWCkdsNpcDkut3Nf6fxyAvmqiOCBN8XH
FvCdhkn8ztJ5q/+AqQdjxEWfVSu8wIq4qJ6faMoDcyQF9i6fRYbYPnZ6qs0mCAAc/GW5e2JKdBpe
v1vmTtXtD3KxBFJeIr4qFMX+8GBVp7xP9ZX6qUSPSRrUfFb1Z47O2nqPyBREc1L8qal7adoZ8bdP
REi2JCxnaCLUaSFIxHHeymJbzrAXBMgtG82SA3YXEq92CbH+yezwTzqKL7v/BoduGDfIGrMCVKqe
sirx4dsO4+OLWfPmiDDzHReoM1JD0En8R9erIiOfOKzJSbBqFzYt5RGy2yTphY4SsZSEwvGAskk1
N/kc4xoO97P2X/plAr2n2m/YL3GbfUXnnRTwvIDXeHP07lK/XrYgLrFdUbQJf9CtVTOj8fL9XYuK
LD/hTsuGu+lMKmscE09oVmGGws+bQisvfG1TI31FnQJcx3OdJdvMmYcrEYLWEblM5lV7pg+4Ic5T
9nCYHH1pluAwpOgYkcZn+fFKdNt3s1Ikzafofs4yRMkwRr48KvK/X5FIWCSus08/r47Jjdyxkdu9
7O5oZfPy0dDF+ZMF665E/itRG2JP3yBj7t9QBIdPEa6V7M2uSmkIl+pe6fH2VNK2Cn0C3OqH0skV
BxJia9yFLvwKe611MWELO0mQQkLFcEsdZDNZjx3KZ9t4nCZcemV3pXJNIJFhlwVbhGgvhu/MjbyE
yoaN8mNwS7UkKMcyZF2EpIaq6Vo+bUMIW7qQmExOiCk/W4QE3TxmqPkNm4FVkHrC+ZegnGaquDoL
VdOEpRWrjSajxay0jSt2Z/mOdlSsMfkNcuWkbOFmD1QY1FIsmTi+pV0XeYWYeMm7Ew3vj60UW8PV
co4MXmblHmirsmRyWxJdxEX+sKJ0UEL0YDZvFi5VmO5NBkIG8huFoirD7wff4Msl3kETP+6QsP/0
n0a/+zhUoMFechLvJElwv16lwCJeG+srAZgO88PevSUWh2tOy8anzSzrxU7/d6iHf3Lj+RzCpV0o
8MyV9ZkTLWQqd0ROPFITRFMPpAav6lGvMWtKVqulAJS1blbZORCPa4bthQS6hl2OmTe0PUPjlLa8
Yi3boayFZdMmaVx1nnV2nepc4d0gSyMT9zzPmW6txYz11N4+HWexAxmq4AmzEGnR87b1Hotad8Hk
eUHoVcUqXyWntNrDaYAPhBBryOBL6NsFUmj8PP1T5zUcgFevJiWqYBQWoIb5eoQPM8D+uatjIfDt
JVW9vyhza9t552+3aajuNt63zUhzg54umee9RwI/xGy0CH7zz1O8dHol6Mv64xQuHf8Cff+DVY6w
V2INQ5tPbmzZDRVIDDERDFNS5Ql0FACFpmdl8FrGTN9A9Xgv5y9U7eJKerx5QCmAWUTV2VscreEU
LqFfPMDMUyLoxUa8aT+4SD3IWj5GI0xj3TzP4vRLwvGK0In1/OqBWgJ9Rfy4vbdqaXhZZxPDxzoK
lQILZVtN4VA1NWRkf+Ss/J1LwjPnhIKQPivfFLbyAHzN2LvKDMP0Hd4wAxJCK+6hRtzVtiROiBc0
RNAOt4Lm5EyiV4ne5F1yPzDCnVvIBW35fbJAtAKmsf550aSi8UwVf5HlWkUnOcTlGXGtMum5uPl0
FNCyeJ7nctq//NgNqzwmYsossLEtP8nGIRpPKXLdvMHJBBPeEpyyF6xv9lcBiG1gZeWqjqhUMGbB
jNlFxrzGqrJfzyfoAwg6ozm09YDJXjrAFFZrBpZI9lfiMKk+E0lq9SiJrMzjbfDQnDAwaYNj6QGK
iXXXIb/npvJRGj3L738wF8kklg4YGIwK19MmhZISDJ9r1ErO/D65b7DH4atTPHZRTU7WoojCC5sU
FROWz5B/wZi8a0yJI/8daiFOOOIJBG1tgmGyU/vmsvnJcOGHkpO4sDGtkoB4yRTh8MmRJmDae5SZ
jAKUMtdUBMAm41kZMwrs7+f0Q+J7RS6xxgNVd7/YNzSECbHXCJrAXkzAwZWLCJRP0XtRCvcG4bpW
gjCLGIEe7ovzO9AdN+a2WP4tvIZTc9B5FvIuHiBtS33PYNRZ+5aZHumNfuayPsXE9OwbCM+ksHgo
JxjIgk2ZnjfU8Q+eshMNY8jfs4cYllHpHmElaPzmWWz7W8Vg+5mj0AzhmO/R2axZMijJPX+ZmccY
pvwRJPyBcxjZW4NX0ziKS5r/eClHTiSImeMVAkED6AmDR3YzOSR0ubJOqEWVdS73RQYj63l6D764
p13dgCC33z+lv7nS+Xmtt2d+N9tgtMFGXS3pU4CzYB91ImqSDn9Z7fQkQ8QWR3JGUbIiudRpoRcZ
fDSDHdIVjLK1lLDDQqW1izMN+lJqxqm9aG4gVw+E9zGaoPAQR2v2Iy7901pBV860HQ4p+UMVbVB1
hGRpHqmb5kr757oPAgS2Vp/kl5/DZKFVgQpzTHb6LTFXbVg7N8GB4nD3LG9p3X3gQwguoueZ2WXM
kc59g0whZxTv/CiTBYn8nr+kx5aALvtIWzUIgzqI8he3mQzYRBZxMDbczyoGkObbqdp/X+bT1CXd
3DVQS+Esx2YE8+qjUDtpKN7tyfdDXkTLOigL7fdfU4CYju0Sj4DhnAZPeJMPKtFTnvEQK3BoWvo/
ntC7DnMPUw8ZbSK6OgktiiY2RHHUQnVDuSCLYKm0Dx6FnMmCUQg+q075GNTl1uwDhmuj/P3ScnNr
i4q87gcLeJmPhS+RAjT+WtQAW/ZpKWLayF1VHBNKt37sBthI0rYwjVKs8jgW8LumoqKGAuRvHT9b
ImyLHqHnmY+DjSsHgyDa3IEKdo6Vah/hXCyyP4vdR/dFzCqWtEpzYeoNXACvVrGhUABODijZnKxX
iuqhcru4eUYE381ciKyW/iOoGSJRwBej16L/VCbuU7Fnz/qIuwe+HdIgVUONkl1uj6qtSrOHlIyc
34feadI3yXQdwkRED8eLO7lqQpxBBH1fZ5czq2YTlRFlST7cUcaxI79zjhOBEhr4PXfwBGBnkkc6
PlAV7sHpJtEcqRJVT6NEwjFlcX9qFuep/y8OqTMtHQAo7LaXcC7j9sUEWvxBYrmpsr7oDIXJbg5D
8LA8DFIS8+nAD54Q0P+AihyKn8Pb7ZR6kKAcJZgHSj7ZrW0+TcBGItXgy9UIxBVTsaRHCmfEtMj2
+CB3514dCWlp45fhlcMXx07gt/DwAYErm5tat2vWF4b+u68hWnivOj2dXlZFMaU8+4IyPtNkIYmw
NszC+grsv1ePz3qBaNWC8Pg3hVyHO+aPME/Wn/I5y6ImeUit1o7iMHc8qJm6oVDB6UuHZn0vm0m5
Vm9FAQ7a6Mka/weMgwZc3bT9YahWkt/+ajt3mM5G8Bp6rg/QTR9EWnhRqoqKjKcuAIzXTTJc7dE1
wZiOO0Z1cvwqfn/9kJvzinFuvyTVMeqKV0d6tqY61Kr8D2cnqHsB3jt0/wS6Ccx6YSPMld33GUPQ
gxqovES59xdiWXFQTSMJgV5/i3SDcSxhBrvWvkdMk/h/5Tmi+5STRsGppR2VVnFS8GSqR9u94YDJ
wrmYZw8AZcpYURPc+5u2rD96XSHhWPTXMqyo8/ByD2jCHIUpIR2dIjZP8izUDM88A7EjvMwlXOxM
CmiXxAPdvKrEnJPrlF2s2+PNlrijt0o9bNz9YhIRDMTiRnEfDl7lj2DMQXMvKGg7x1jhztm4zJ2E
rErHhApDBSYkmkLoTyxQo2xSvKm6i3ej/uB6rybUr+8yFCHEl/QjX4Sn1wUetf5Dqjfuh/NhIcbO
l3E3dPU92b33JFNegidVXYX+p864WJ7x1W/cYcY1gsnLtFNasbWu6eJDFqDCeq7ol+cJnQG2prUx
dDbF0KPDdkfvQnT1dEyexKeszJ1hsVYLr63CvzcjbfK/+qe5GwZWZRm7Wuu+z/Rt6DRxBZXOg4Li
4BaU6/FRJR9nu1Wh82lV7vvTXq+ljxllb3IECm7RYGrY8Q8H/3aBWccjbLzbiK72iCk8hlnw360K
L9xguVNKY092NoIPrE46szP2p9cvvVLhs5RQ+El7QsXGxd2489xMW1pk2iiYQTRZ7cHXun5TLPRi
aVLsL2U+Y0JSAzSwX5xI80pcBc3vxFfn13+CH0vcih8ZFwzdN64H6+mKzVU9qoGFznb0qiGvYNTc
ME+1lPQdiGySWnFv/gJLUbQ5jyVa7Ec/9ZK8xJ0NUlRpIIZ31J+jVhVi2tUzA5/9Nlz/WpubpMx0
pDGWEt/6LHVnG/HHtsnIkbE4nV18npSRrEvnHCeanmPP0E9LZYQ6IsmhsfJdoyvtNDXMeFpHiZDi
L6/g0IMgFEPE49n0Y2rfE0OtRExv/mfcbm2rIpyRV+tfN0BjLRDHpbAEqRp3CJSqsDBxWJGA8XXb
8SxgpT2v5EBP4RC83EQMx+lscCBEvh22zmdOwKt8FpWs5s/bH0MevWWE1wgmtyIiBek3Z1OI8YhK
40c9a5YwOkoxq1TLCaAlWOCesP2BjSzcRx8hoN0kp0ylROhDTp93WbQQJlw0oEe1fkyKIF3OTiFw
p/lDRHEXmuNlAyAZBF//7iWOnif6QG0O5FSSmPl+0AU6vk6c/IWEIduWLiPWO1rntGXCIjB23/ZT
nLKPYg6XdjK+L6nHSSjTNmTLLZPjiqbGz4MPsajnyBkMFErKXIS4qACqu1T8zjLG72XJ1wGeF9fg
YMmeJRJ/bHjYxarjvFZg2jCFzFylFJfIjSISyPMl54QbKiR0MOfQ6jbppyXSYMgTFb0AhWQqeV3r
0f57VPqOR1Owc5Q0IEkkOlTlqqWIKnaAB+1hcp0TA/lI/nTd7gxxmeg7shrH3mGwzThTjo6dg1e8
hwMi53otCmdujfeppUyKB72oVJPPE0AlxzjukQLdykxOXoLoCh+A7UX6piMWFJ+gc5nRHKALaSdT
yNAayxwt7aLP/O0WIJd2bwpavn+FjgWEDU2qJjpbAQ1k10e/xIU50pjYgCz6UjDpADR8qov4F3WF
AQ/N7/oJIVndx3I9S2MrY5nYuHo6NrHKMweqRf43cw8Mq1cuUBUXUUQyVObU78bvdzJRwz4FhSex
2dWUXQDIZfzUwt9aWqvLlxqT6i3dqu2XP98rlDDmVuWGSUREMecxy5NRsmNlk1MXLiaKUvv3X47w
3FtD6Ds4RU/2Cuh3hVPFfhKE47WTfFv7FubfVy1+OLvAGB5dYFcZYKS97a853Ld9FLYgjdVfXRaD
ZejO/W6gQYX3CW+VCQLcf6L5+HoV+Y0XGs/xsVvFm+lL0UHh95bHe6H3Aj5cRT6DWhrNT0fXx2TB
HAQAFuVGS1TJLypfb//RjxWDLcrGPJM8rpgYDQ8Wd5YucYitI8ESjU1x/ukAaqj+vIpsy/hi2som
uWi/MqXk86wMwMA5HWIK5jmQBLEap7sLaNu9koMAUr9CKdPEnuZUVuKbCC+n+d2sZsFJjKL8TN1V
FACQ8yqg8WwGlcyj7t+y0IG64wXYO3tbYYaD2cq5+mXDO7j5OessyJtgj5GfX7wqLfScsGsv/xfC
uO5M5R0Jt6FMSELpjfZt/Rg3+ToByUXLjwx3iwBerNcnUflAkbxf5lltBaV3OgsqEfcgVMQgVSzJ
HdQ9eL2ArJBnlLWAPVE9tXqeD4eY3JNN4mZHiG/BhTmbo5OWbrKaPtOsHbNOi8+nKScIuFLLA6er
Q73ZOXSz/VKAmu/jllMe84OpZ/81kGJHDViG7e7/TD30UnmnMtc2ctfj1lx1X7i/XTY6UqO114w/
R1TpC5h3X+6Hm40z+bgaHQP5BT2oCn/p7suBAG4WBmfMJyM3480ARGRdvyFVrio+XnxYn4kvNXlE
v+dq3zXP1ru2wvDBfAGhBBR3n+Ve/fmo4x1ntFipQYotjyia0WbGa5H49eebOQDtYNUUPh4yp88v
tjiL6OSjRP+Z88O6wm/4mIGz6Br722JRJbqe+c3tSs+mqEpuOMlPJtfQ/rZOAL0vGZ3vKBRvPsHw
dVtCtn5WjOd+EURFigSRR8VWMNvrbfFhiczMxbo1ueRJib+CvvxiUfvvoKKhx49qiJRznqAoUzh4
MfYoH7QterfTnG+N0srgTnQpmIY8GoFbzuDidLb3GHO8T6DUCJStO2lav6OheP1fOwC+coQBfiEa
ygu1B/Cz5qhF9NtcfLMluTEC4d7JrzGO56ZSH0P/q/svN/PX+p/rF7v+ly2SQPuYXxFcvis6ILPT
yjAaM0EY0iGnpx8Yiz0EdC6GpTdexK9rc7qBwhT93LlM3/Bn6TOyba5pF7h4O20JYCPafabB5umg
M/xCzfL9HHJim5ldjZZq/B0WHSrXC7JbkKW+VaeJgklyyH26iNEZJX8Ye8k1tb7SWJiwxvEJ3GPY
bFMZittyMGYyZoMB/ozjcaUUWyvhCbjSJ4ZfnILqKiD8Gh+KmEMMfu2TeOTu3u+e03oDLxKvwxie
x7tKQBgJLt04sBZByDT41CNPV5CI8J8GBCuSk+CHS6AzPRRPfkeK3ZO/MG9x5PNFZhO4r3/PF8vf
WVQfvA8REWeAior/uCP90m/wyLMChVthNxd+J1asDDDGRaeYOm8W5HSoIOlRhrsaCcGx6Aqu5Mbg
odHMPO1A2YNEWof5D1j9gkRoQYtM/lzPcPLBxMjRmz6ckwrs5gkAl6254YlfOBcCRy7U+h/9ndta
h5qWg+eNNG3PF4i3g3HcfPHRrCRXgzVj0HzuKsNPGxloxoQlBdcIlIcqCJgeUGD4JQkDVCKycDub
SHBEVeCvj/2kyZ8ZHhd2iPQC+iiH2UDHsbo51ZPSEjBdgNFd8wWQTMl5oGDei88LLRWGEQi9u0Ke
iByZ16s12YuwuoHBGGh/nKHtvATOxmyjh6wOTiIi800T45OeFMdjmoGYjy1cWRopP7ZuX/ys7fWq
4/7Yf13rDS0HNElc52YEnbWPZc1cdVeAoGIObyjwvf0rld85vor+CrA4FCKPWBcFXmqFcVgi+Z6D
nfD/2YjI1GWr/HfB2y6wnhQIqPdB9ZZroGD+WdsIUZuj03Z80Xjms/YyXpkFrXLNiq+krrsAM+VW
AR63MWKVqYFBcKQxNKaTN9O8WCTsEVbsD1AzhG+pW6PRe4LTMKqNiPX6eOTkr4MsNGdTSDj98E4i
PDEnboH7uONT8hzQT+tKMpYZYJ+pbW1o6tINEqXBY58LhETL+0BkiwlenwoZVM1PPdCJtKPCqykr
s6FNDBaB74h6gHv2Mqls/SE6k6et/oHp7QfYqylypcc1JBtm1KzvG/yvsOXXApy5lp5ptWgJY2/h
6jfaqi73bhTh1XqOZug5NAMtp1ZhJKrDULirSP7IvbBz51UFxCtsP58nd9HZrAs/nXJdInL/GDqy
Nms2cyfJF9W7uPGbe2ZiLHQly81PwqN8WAwIuJBUjiGh0BMpa29nVFdxMKr3K4KotcxxAFtojvl2
HYXRHFOL5okFM2jVZTJCNL3L1H0sJUGJpzbCgmfKtPK1iB5sNEu5ykOujYai7dq/aA/pb/rgbR/+
3C55EppYm8WZ+NoAyGXUecrrxnSoV34y39Vfddx1mBSQEtnMdp+j1ii5zo5Rk+8908yreqp5+KtJ
fxkLRgxKL/CnwCOKClcNbxE7A2TmY7BxNdvn9vRNpAbetx4pCV9653l8nUmiJ2y3Hc54pT3EgWV2
5RnSalHQWpqXzZuGvmw3gE705CAS258z4IxQb/8/bpMnUYcPcih6cokbrasknxyznIMehAR7srgJ
e5RDgRX9QT4nYRplHg5HJklQpgy6ASW9cZUJToOrKFXhQxREzVBN0zEMROMOicUM16B4Q1vUHX/T
IsjM/KWprQ63zZ1psNWo6238s1Gt/9pylcqtUsh0jzV6iBWbyvShKJXpDa14sot1Rl27WYOZ4dJA
JAICQG6BqQVRl7vB5vJbOgyRHGt9uuq8lq/51rZuWsLh/dY5AAFPf+4mwrHyFxEqVHdTQrdZgFoN
5Zs8CvaCJ4WZEN22+n96PwNA1anhA4h/fhEIIX5TVzf/74CzMJPXoS3G3eZIoUScFItDYmF+EID3
nRAVO3xIMIQAxS5jfF7ff8VwzaW9vH3eUVcPwSpMclXt5zf9wLmMqB1Tk2fRSY5/v++dDHU7ROJG
61cB2K9GgYo6ge6oRQvSYjfinHvftC6/Sd8M8gst4beVgedptsX2mWmzEaoxbJ2XNvlDeNxBQhqS
P6iyg/QLhkH8D8k8HPN2OqULALhHgSu+LF7Cq34hEwLw0TAtMOYzoZvQbfoxlt2ka7pwGt3dG4tV
xY3zTUa/BoH/kZlcrShD++8rPxCjWedgTxhVkg2X5y9M6Dn0oXaJg2yFpvSXiKrjT4tO1ejrAtVV
GNVDVjXBjBlk3H2ZsRMUcm3cszXP01cDImrg6LnZMAcCkcHLYGaxtXIClX2eNSZhhPqfad+HarHL
yNWmqD2sdl3tOZTE60DPmRlZSPdl/Nbmtg2Fp2AQpTFjkwRQ6Sd7ChchbabP0d0pabR+abAQ/DQp
3MrWalPFyLVN0y936rvbV/VbxxDpzVX7/XFXrJcjKgZicfOYL98meaHQTcyLW4Xs5jx+/+egudGE
xxM66+s7ia2DG3uAc7VPDByKljc2f64SiCAoZtdNeP8jeNEwlvSSRJ0z8mhi55gr/ZFD/rFtxykr
OuI0Tf5WEppr5HAg9/UrDw9QMis4uIMqh+7xbB7GO2LGIb0eOb4SactG25mW213t0iUh7ohYOk5T
z3G7TetOEyJZsKsoJxa7yoQghQaKKLHq3jERCcPPybS7sDhhz8tQ5qJbcAKO59xHWaLlB/hjJFPx
cZAWDYy/loR52xmiCkjVjHJrsBPwZzTFk8eY/wTIGrWcB0dJ94EFdRWiqFRiTaYVczjvoO/5diKk
OIAtmvgiUURKP8FSCb1oCRQIIf8wI4OXgQ6ADmIDRWa0jjfayW5o5iMtMIndrnHTwgyBCZ4qYGqL
O+XU7zdrokCa2awQnEIitZye1NRdMbh0/CsgIMzZ3+M5EbFE4atLRLV7vKInAvuAVnqLg07c+/5Q
iCRrs9zyEYGXZ2ka41l/eFBvesT9/pezvA5brzWZsMOaphMYaSL0E2im69/uR8VWNLvf9OKWL8+Z
VFJsSLLeJoec2R6WqQTd6LIa3Y892cfnzXLQSRqfc6rKoUZ9LKFHC3TSVv1+HWYfW2erWXoAMdoF
g6ZAPYoAQ0vpmiXVnt7RXVFnuywJML7Q/E8pmfpkpZ0cZNK1pb1z1q3XD12nfOU/SO8x1tbZQ0H0
Viql5YVWqZ0Xd45szSvpnlDYIMyvAPXy8f2KHnkeiev6M8aRMa5Q6nzZ45HoiRzxUASgB8o6vQaY
pG4j7Av5bJ/6RjqvsJsRwpBxHdJFDaJa08SIyJxZTKEM0H2y/0sEoPKLCTAfQBWjyVeOYKaFs+rh
C//3Q2pMdWyDubUHW6ua43rFsjt0WGDlqNB6+HQmA7aJ3kz/AP54DUxprqbSqvV96uAeoGDKXDxr
PX/BEFxdWVQU9H5lrPBa7XHH3BYYhB3ZOKpc5vL8QjL67oKAto4Q+MXXBafgPSVGN2v5KdOHe3Rs
bl6EH3d+BwhoV4jWK9IbcmmZYxZ/ew48GaDdub7BNN84Jx5F7sy2tdY1WzxyOZ4sOwy46m6gMsho
Uob/KF02ZWdBOagHdjUNoUPN2MN4fiJae+vCV0b5/2RYbpzP04QY+ni2I59/9oBRt6gKzCC/s5yL
CiV2FnX2PbcpYLVewRsR6duz3grGzW3ZxcOW16yyr3DMrxHwwwS7ektDAOC6umE0127CgDvvLHtN
jK3R/lAVo5iP+P1uh52wyYJRfngs0gB2Jo7dxgv615IzfzSgMLxmBUdF+OCRQN4yngrMimMhLzES
FcCE/rbfKBtd7GKC7N3CvQAHUVsreqsHbk6fio7uBqRhmSYS6fw46hyIBJnPgQkn/ePhs7c9D7mR
iQnFYboyvl6nxOwM2JQCyiYIaVO98lLFv+sX6pXl8CKEn9Q0s9ZC+fsREx00nqt11sF9l3apJ3G0
vb1JL5LTyBFWQ0xg9KOc3vCQxDt0jkf5HyKZEfgvDAOqm8awtWU2PLwFbS/7eFVFhgtQe5fU0Xbz
gC2ceuMXHFfIOz1fTY8zshv+162FLetPmivzveCmMl43dQ7iDEXDGzBZehD48DMggeYDVZGdEBy4
utOarTlm97JqoxLGejwInf73eVd89XlK7io+SFuKjNQWHq4YIThtAJGJxhu3NoNOZEbPKnt/Em+O
/SBvqLZ5qZt677vBrxoWCWg4u+sZ13SnH0KuipgZWr2CfN/BckUhj5+kTcflBIl61Q9cO3FKWe+k
ZjlFMkA0wWouv/BPxH6G26W3GoanKxwr6fRdouE7R4cX2VWiudsEx2Z+F849gKaE9d9lHFu1C/so
jVI479OfJKp3u7yMS9UgciGcZXPNUg8b4IfbwLtLdQvlH3X0lfqdSXjRreEUOM8GwgX74BI1IA14
SA53WnR+pBkbegxOwc0fsF4krAElanNV85wZfGYx73Ab5KV0HgJkY+62/CsuCcd1rAfE0V5esUih
EMIpl1XH8xctU5A03ZrGtKoL8S5N79l64kWqKv+r464L5Zb5cMLdhwH0eBGyZBboW55SY2ZYNjce
jLJE9o9hFun6FUL1K9ciXl1nKCU8mk/xGvhCojVWDj3FkNeTyvB9l0PD0QD2wptJZuHBgQD4HKsq
TPdQOhml5bRGFifr9ghowbUoOz7MFYFqvViTnjjoYQ396gdil92PKq/9igh8PnKzcsTSSBVzi3GN
0K/bqIQP/ZN7WGCDJ7rE3JeG4LUaW/Fria25GMGPsEzrpoIThjlWy/cIqnbWruKhtH4PcneS5696
y9ZKlB5Dw0v7zt02wTuGFJjUMEbQW7GYi4TIqexELIrPRPcot9Ot9dIWjt5W4nm+N2b0siZ6PFAv
k+1+quKfrFeokFd6AIUSx9xFhFuJBCR3Ebv4G0Ag21xp9njmhEMNvMslgPWdN4soQ+Eqh+Q3EYWi
4h1Gh6EKkqGqRk1irL/erHA0pFdCXEGqerXw/qilbxGCrftI9WBRDLZZCrlk9f1LPqfT/oRXVLds
Z/1KfX7YcYRUKCOVr769Z1LuIUStKZ0vvyynBey2Tu54Or/tS9Xz023K8JI7GbuXdtYKxyHWanGw
ooifBdxmX3j9C7FdUKm2jZfatJd+U+1QeeofCCdx9Ghu/klasaxFJ1IikefLJvOWyhH1TYZ9odJJ
YHJfFwYDho/5MajFsH1GMHhcOcIEWbdJWJOuDyaL/oXCaXlpjr22l9VyFGPxurxr3Cc6q5JR4ea0
nXKe/sfST95U6qqJHvHvTWyVgaj5dX6kD2PmAHRhKQNw0Vk/QBUbc3NsoXIJkApwFfNlvZaM3Ndy
FxN7qRCPk2j/DDKAJAeaqGMW5v9lT1+xqs7AEPSzh/on+mHnFEqwTS4+qNje1G42anhtGvEo07nf
2AEunVHLubPBD7lJ+yDd+1/gRPwF+8O9E/miayq1VW39nlCy6vx7cdRrFqhoIE3a1tNzauOHz6WB
y/7Fgow7FbLpWYCVd/MvXyn5+CSEmlhI9mQeWBJl1Tcb8ss9dLPmNJg8mbAxeYyiU8w7IIuhbnJX
c/K1VhSOYIdgbfDmGPDA43WkmJD7tAj8pZSIlyPCTPE7XS6ytfkCxu+Co5iYJ5i9/fhU0ngyzxz4
0BHgw4oCllocaohwZ+fMqReiJb9MCPfP+WB4nZgr0qimlzd/wlxbxbJZNRvW7JjXfwdoddR27Smd
ZDrE+YZTgruHomRwojtT67OidytfAD3LHGLMyeJa7to1UN+5lSYVK4BbG+GJZN4wwHYutQagjtXV
UBuZ4O916+mu2RxOBWQ2FhlO0j/slQE9acpX//bfqiFQ7w5E18JOhG/9PYzmNmYR9VbzraIiWoFn
sPbPHN1ctb6w8n8LtIP/X3Z8NHthC6kfn0F9vX5b5zGyrOa8RlzZC3T6DBDWn+vE+dwUxHMsWOEf
nrYDGJaYOMKwLHTlZc8Ab0Ry7qdNbSYRv3KbUD4dWFpMiCdJqjTH3QkUXP+WXwewxOY9owD2pF7k
x/KE64/ePo4x+0t1Hrydc5tIgX5kC/Tzo8RLg95rcwte6dLKw8SJqApajK3UdkpUTaHiKEsMLavX
ZqPQPSMfhUojdPx0CPsdbE5tXqUE8G3jVoMM3imoqWRtK9eaDAtaZasKB5/qSa1Wul+6h61FLB6C
MGmsCvs9aGMb915AQae8HO+t1zdWvasr1fbwgzTCfSzx+szHNh0EtcVhlwGTKht68HgYRMgxj2UJ
DKQ/WzLbYiJDxoDiWin7IPVrGmjdeETgaSIiQFwrdUgpUfa/Kx8FOXAo9uNf+exMOmwtgT4Var1t
lrrWMOp5F6tEhoiavcsp/4315G/grXyobzhAbf7QAFqfrxyhYFcnr4xidKEjnOC52uYWuNQkUJIb
Y5OpmRmjcXFR6afFyCyncsJA+se8lM8lVaiHmRZass+K8aKIfeN8OOW5hYKWiD41qpjUMbgVQEPU
/52BCZqxpJJUo99SIIbpzY8/BNhYR0iPW74pgatjkKMZpCtIf7fJCiytTQqmWLwgQfdl1tIVRnZG
hHhmsSI0+pso9ahYs77/xdHvnQ8Uhk1+2eQpIQdTgpxCfi5vh/bq/TygBPQoOe3a9BI49xoiiMb+
vyZFyiWX5ujdZ4HrGXPaHjwG3NTrpWK6+9ogHnWzmVSippUN5CqdiuTTAlr8XpYNXp92LMVV2koQ
3vFC/hkvQ6WIyvTVUTVusHbIGaSs6bYQxIpKcEXnjOyaqFhWmx/xONC7WDmGLsYoE7IPo9wUT1gV
shUJSXuOikAirwsQGJRxyaYMgIsNluMFRbpFmXqLRNw1uysbbHnkXew0rT2vYCrEdYxga7mUDLvk
IP4+hDY71F3yvQvwaw8nwhzUY7hRJW0nKSXmH0yql/Bk6n5obiM/a26ZG3B1jr5nv4Pk23SddDHX
TvYPCX6SYEwx9LsJSFMPOGTgYdfqQlsCfPgQMLyaH033Lp55myeKJsUuuOy6Am33Tot6PLIn5qPv
yZTPNA1kNR2ad3dG803lXdw0sEpTRvK+oK56+EeYywrXoPheNY4guR6db501DVUFrP6jctxAsdwM
44yCSo3gTf2G9ueKRLlkQ2Neb6zfTUTsf5K2+7hNQOa/LBMBgBL1EToldX6TDOMEt74G7yQr2/HG
3qxza1poUFMMzKPK403tHCypI5oWWQv8zkYu4klVWPqdWVfsSOVd+O5T2oZn6MCLElt6MlTRtG2V
0h2rV/OWL2EyG0iMpm3wjJFpH1p3uLjfNcE4I9KyUpi0NLagAjgyzjrDAgWeINc/bt7jlP8XClAr
zrbw4VxIj+OVQxYZQhUDWys0ISkbE6ujrW0sFxENsLyjn4cLYnCYF1N9313MhHKNGZQqtHMp3wu+
m5QkIa5HuY3sT44bAz+xie1zPOWF26lLP3d6GM4dNyzRP4KlmMUdtDqh9jly0Gv9zZZvfh8L3Zcj
KSKEeezyqxIq5ccNfFsvVpNZSTvAi0ihLb9IhecKkOpX2WJ73swtoEhZ3ZrmKXUnRmxJeEtkpnXp
kH0mOMrHiNWPL+SpM2vJsWive8bjkKI1Ch1LMSs7cYG0JSeQC1x46G0paa0yB4vq9ypBgL/+9LRC
iJMXEt7kBWw/GjRB42ngRHkCpnqP2Zcpu/jT1YccZjcydg88Qd4GWc7kOQtSDldKiTrTXTKGIcuY
m29TWa0kF8tDxOEMXsxhCL41t77OcnSU+l2vQWJPA3ObrK4OK7hbPbj8vQealpv8U+PSWk9zdYyX
mNxXsByDSvy55+Vr6+nhhXq5dVcM+JKe3VYPgVCg1E95z9TJ4fhKNF1mRCr9gpUxFMgq4Jg0BTLm
r6AWZbwPr9Bp3pePlS7szhH4hC3DENg4rTJcYzRlBAF0YHacIsNhSC786oCbgbPxY9HyRsV0dgWd
wmQ2LUTAGsqK07sPypxHNWb9lDsWfyGkqk2ls8+pHAq4ikA4cPZ3jwBgUEtLLL6BgH+kSxlyVWsl
LgBIScEdmHdabs5r7y4QpVcOa7+pfa3HrRI2rvTo4k+3Oh6ak9aKWYWXNdhJR6eeY55f6mAZLZRT
jU5vDUfYWv6p3j8WidaRZOUu/N7YlWMOh7cgKPJWLycbGOvOsS/hTaz7LFFH1wSDttnJcCZCjn3U
1V+u1Mz/XOa0sONEZbOphTL4dGvCBuMwdmqQXcbT0l30mPJ2+9jUgGRquTfPTQd9XZM5AQKg9GC3
BKGK3elfDQ0FMyK38XlZuh/Drc+B5ZXnLl3lfrSQZfIxrtcs8M9pMmmhyEoEsD27quA0Y+XZg56m
+OAPTk92PUf3HVv7TnIklhAuFBNRyJlvljGFPmWDWzbRlnqfsr84XaxXH49W/F1fTvKoI5npXCkA
EJMp8+k0hiwr6kgXUrJLeOrHZpvLkciKJZ0d1ArCndWZlN3w+4tKWILWu+BxZl3ZF0dWMabozEs6
Bdjzs8U4aPcQMms2fwZe4QKll9GkOAEY15TG9BoqyT4IM0b6MC3n5I1QgLxXi9dQFGv1ahjl8m4s
FqHGc+0fp9YWU/JvhhX+MWyQeXlp3afsarNqqz70dmUjPUdW5B1dkG+CcbvUjSnLTIxyz9bDvzHs
wBAGWY888rBoCJL73s+0TMOK/8QZDNlwGCQ95JgwfXJ4fCXt1GU43LEZ9xcXG6hgTvWBhbfpMz5I
mcOBeO9xH6Bc8niezyOMxlJuH5tCIjKcrr+K3x7r61jMEjslovwJbDLNnVxZHFreHzhUf5svPD0N
rUDE27jakyUZBkBu69ebUQsumQLE6zoRHO6TcExfchJeLhZJpT8AN5+8NqwR1lNMaT8tUVlwTh5L
7ajhe8TCp1q89A8BaZJr3w8QH1hCuxLNhaRGn9bzk/27xhOROEag9/y7GIwwQkKbu/BmoqrDt2P0
5QkTdEL+ALU72pmB2EzywkFJZSxUjBrAx5RlntDFXdDcSUG8dh8CrdHjk8nkZbNhhkWQYI98HzTI
VRdxJVojixkzGbq8AuI03omRG735+j1ANgm/di4vqHdsqxZvpDD7z6UmA55NuCFtQCog/kKbXQOG
/RtLOueCgtrwWfmRBkX7R/LA5SIhGrOINe5KVObPHr9QW+7XHYbHNXRTVxeeQB1DO/AcX/sxh7BN
q/ZKWOyQswFjwEcQJWKkZE6TzIuwyGXs15xbQjFTf8ELNAeGU9yefDWujSEyPWu7BO9UW4iJCLYm
wAaYeYvbHdv/s0y5xc2b6oxlPU9Ixp9kHUSQy7mPkhETKj5uZOMhCioIsblltS5N4dah+vfi61Qy
aw8+h8r7P+UK/KUKrNwdxWHXCqQzsaBCSBQao/PDj3+hnM3inYOzlxBXsFJxZqgKC9S5ytHJdZ31
03aN4qYqDu6H7xfGSmysshacLZR2xprMQjg1OQaBeT4HITpb55KcFQDdiIPUEzlc6Coldixs2fXt
+RqFRp6gSzGI1Aufm8tgOW3RiFPb4O0GgJx38kfsN8z56Yk1dKzH0PENftdPxmXTVHD1AXjDw7yw
B5caFxvX6dYcmAz7noaFMcZWVtgp63jzn33n6s3CxhJlJzUx5wdDWnFlwFv3L4iQCzMQ3zLMn0Us
lrdn5g/u6ut86pSU7smcyQ5+pi3ZKEMeLlhJjUmxI29fRHcUc/J9625z9qBykb9mNOBqwUjIdatl
8R0yLt3AVoVYSi2V3mpBzzYKSRO+MpamofvlVNWyz/FXu+5pyBsf8xHqYa+7dMWTSAuqUX2NNQC6
NL6+x+vXuQ8BH5NMOx77CwQSlX+fX9pz1mnMrx8KxN63xrosSzSemaU4PqPdh11HSReB0PCCO5Rn
on53uW5r7i+Ju68sl0AEjHGSFyLQM6orHcuMfagf7c2tqpgmwRZKumDqP/TlzTbRiyEBLDYaQq3O
QqtIM3QOm+Vi1SmFI8wewUnm75LM+ieMxKRI8GKtIx4e1sH3sQTJU41/2BPoELxzktY0PEU2JmP5
fUEffQr67wYSvhC3JB6ZlKovCNHU+3BHyM76oJVloZHy1HRnn94/zRpiA8YyHfKf4IxELTY+twfb
WdwKQjfVmXhzWYaXEhANkGCH3bPdTJLgctVx/bLS+3AaaO1NnPU2e4+djBB/Qn3CZfhIXEXJgot8
not5jM1ENp7VyYEmHFujSgv20QHxHEqPGx5y+d5/nzC68D+VsnXKAPVGe4dPvBAaOJV+Q54WI117
GG9V9jR7Ul1FmHnvEyl/6+bPWV5EzUIE6QHBjog5mL650ID1qzvcHB/phMgH6NlVGQ1MsoKEVEWf
pTgU0y+3qsU8VwigmA36xgcxt1AcnGj06IsEOOqptF6xUhPr2IH2nWnSGjNCJZyphtvNByHVvdHr
il2PVXHAS5fNDTrKLEQ8U9jlaREbD8YfQeuX80ybFgCKcg8GHSOqsgrTyRCKKfIKtgpKE5Y6uZPp
SlYKXdFQFJ01WQ2LxdDkIhM4hN7DMf2126wUIuupEgXk5C25R0wJZIj8vpstdXmciSF6lm+tI42R
SbKonmP8q7ZK/vyVgDdUixhXuhJoh+RyXYuOHNlmIpze606A/z8eBPp1b4J0YfOFYBXwNp004Dso
GyqoBca+iZ9/ytXDESaKBA3lTYTV9Qgcfcx66RVlC6KrDarZo+J3IEiHaXRA+q7oivbG9sAosymN
cpV27n9GXvHBEBcBPc/I03YC7i99hEuM/aJ8LXoNFqXnXSfZLJU6T7K7up8zZqZpYgDoun9Lup+P
Q7GYJXSsDx9w7zL2Xg1jSC8V8a1yny0kfjY/2zqQr1jPg9n13Vs+eR/TtYK6EJT2fHIUt6pAIBqC
kKROT5fFsU9QlQVbQY28j+pKkLqpq7DR+PhWtxWwYEvp5pxrhYoRIRyvm8dvvQ12DbdvZfTrEZCb
RVuIGN09LhQuMuZKrxN3LxkKM7igPSLsfIrU4FJK30/u3lnRq44IlgI0zmB2JfM9o4LouOOlA1W2
YHcMECKd+piZm6B7q3c5EVAfsCed486uSVMZ95x1fu2Hr6WwONHvr/wXveLNoQ1SPim7KDD1uoVP
/yc7fJE6vkj9PR1UAweaMjCUveuzB5hq40oazsVP4X9AGeZzgKdSYkWv0ZphLVDxCQhiyO+XlNbg
4lQQDdkDbmkwOnXGUL8nR3TEoMKns3cGZao+OPiE4WtdSXJieukd+y5D/EZt+jxK90sp7iWd0f/J
HpA+g48s8yPLIoRmjCflWI9CaxVhH8BE3xWylFlqT7Nwy+tJ2PIHQfvWy3t0snk3V9DVqIeD9zL6
IUbLMxnZ9dYnk2xpYjpDyGagEeuDU76A/YphsDGSQP89IbsNygisH/kDg/PdKfY/T7SFBmK/Bhp8
KbkYHsJE4MR9LuQ5+TZIcizCZkrzwQXSH3jH2sbKrOGki3JlMBwBuNiEgeiVpGklBS5OVu/odluO
TunYfFdfdmjR/Y4Zu9p41EDEAW0Hgjo0syoYd9iHj9pQaEkCa/BIDZlVx/IFyHczW4uPX68nLoOY
Cyndrc5RSQ/J3os/LKTfhxidQLB3iIO+Jtrk3hdWMLwJpSSdLccI9kYfnlDxhQ0ezzgJwwA75+tT
ZBjyT8tHcGu1fonPWHePXeqOnk6r/82C+Y9lrqG0QYagYlL9KIMCKW8L6LkqLb52kas7PLrn6akf
dcI0oXWrC0BX974aRPFvJJaqcpiLa0Ir3cEKeFH2P/uLszKA4Rese9l+AnJc8sMoQ8A5dLICTviE
kRa4qMXidYdTwcFYWmssClNnRy+ilo86u809gzi7D1dhAWiUV8SU0mZqdmrX4/1upOHlrOT+zdgu
UQaNYdiPKYyDH3PlEMKbEGy83wwr7kRRKXW724RJAmSKKxOTWszmOHirU7U9iKMViL1lRHQ0uBal
Iv/jSl5WRPrErrHvcVQXhy4pYLOGP8bE3srAji44w1fP0sBkzf7acx1CXlzX9G2LaLfjgS66tJ+o
A0Guld7w3MfL1vtvkWwlY04lAs+HGKBAmLaOsyi77ev41+3Ky/OOMLULJ6LHtDe0KA1V6MiDBuGf
V1wzNQP7GuaWBjsaUdhm9OuWqRgetjHd2uGZUBQlFtpsy2+0XBzmXDZbrKdqnKAc9xtJJ1HYLbPd
15T5bfwnfuA8BidMDbF/f5HATCi85Z6uZdX8DY1cavuDXA845WdIJ/lpByQFPQL5Ga64M/sF74eH
ICxnAd8H9Ru4cGyTUBfxgw5DkrT5BassU4RyNP3yZu8TYxBxlxtNNvfUzBbhxnAvfFRyave0gCmW
Apw8q0jbHjV4Bwd6fYXcg60z9KYIG2QS7fXm+XHR9msNGUTF/WU8HG1pp1qhU+liMCCmRD9v0Z+e
EkXsYr/mHvPznHr8uScp1wnHVInyTZ58qgBMvhvQ616XcVVcHLYXrx/BvpS57qJXrZRHmOdX9tqY
rlcj6tFupDmGx7FXgxeWNxu2nvWknUh65oLJycg+XntXd5vNc46pg6MOI3GoM9MP4M8mipsWwk4d
itef5T2aS/V+cJDl3WayBHF4cliSjyxyxkDSI8aTpM3EhaX5QSUX/SkvJ60mdK5Y5wzn5i5Zi6zu
S6YjA0Hx1XiNXlQ5xWmrRuYJyJTF6Vj0wzlcRoj7oQim43y/wNjtgrmH3iqnpefgOFyDb/vA6d/G
MLnx+sz7L26bvb1CA2i/G10kzIdSVWudQqzqIVR0JzEDQ6VflQO2FXY16wBP05TZ12maDy0f+WO6
pBYa8+b3JY3pUHPf3c+WKNuExDZ4Ktx6rkZOyKCkzMkWA8rk790MSjmvpHkOv+IF33rjgb/xfKcN
hCDbQtvW7+9rRZ6tViza/m1Is9cBDfLHV0h7UcD4qmYO4nOC/uuLhewNDsejWWSyqRGIRWQdsjTl
Os4ASnan5+q3U7ayXQEr5dYY+V3azoK+aYfGsoUYgdV96a2naEKjD80EmvNxZXnNWn4o2YuvLrNY
Aehr7TeSoFZH4lFvPY8kqJpyMDjyEIGpS5inULA+Qk8mcgu825RvVJG2AAoUYQR5nm1Bgc62Eb6Z
EjrAg+DGgo712b/Nll3unY/9CVZ3ofjkdOhoBc7uQis2Kfnssn8ECvVpI/ZPdaW0uSV9MBbTdplM
kLGhqRXv+7c9A1UuC17Eg03pp1Wb0IojIeYF//w62DTwjj6sjSSjBWRzDPHyE6lp9cNXKSa/ve6E
kmeWR56eqlaj2bIQ6HJ58gqwHv/D5g0ig7OBlmMTxzwiqGO8POEIwuDwIBVTv0p8XonK4FfrXweh
GR1xdR4INZr8mKpBwIGoGzZALO5zmZZoFIVN399MngFQmCCb8DG0ZmcX2mAP+8ZXYM3KF7Ol0P/m
8DyOdgK++QghWe1OKwojcc8kUdW78fnS9p9d2Anj2mkhBdlxWd6c8wZCvVqcWS2kfzysX7uYGdjD
gKuOtk3ITMezBk+smWzPFh1Y8MKIHB8+cQWtARqLa2cPS5xzQnhBgbo3IgT5KHPpBwwARFVJa9Wg
B/lDQ0xhSAsI+qp9RzJeKy8pEEI14+SOU5Ng87bKT5ho4WmmVpdENFqqR6SQRhPjOQt+uo8SGJZZ
qcS2pTjmxghdFQ8Fq5ed7p+dlh9vJ9mfTespaW8Y9dkiGgTrLlOXa/u/7jOBTw7XfChisqEsWAE9
I2qUfPhXNfoMT7ZpU23KZJQPm8WrMCZ/5HqOJOpAgflsQNS8Ex81slPU2gargtuZtDXIJ7sgmxhc
f6OkgSXhToR4AS+TFCklzr8SzAtV4oCCe8bjPwhtYY9bvM2SiGTEZKA44hw+c149b3UryIJLKTbU
NXA3LDm1zlVuD6abjY8FMQejKgiKDWjvWThfFY56wjL6t7dtRyp90l2KOF5+zcDsBj/V9waZVj/K
qPLc7GjaUj5jKWQ/FRDW8lUxgSSx5XPKycimUfUu70Q7AnahP5fU7fC0VztRmjH4afg43lrIwaY4
TFiT+vTGd97SOOfZNxJ9FOuTBZDVc9L5TlBnAReg2Tsl8VJCMqyXY4S/eT5Wwi9GVOMuTemhFT3z
8U/7d1GQbGHr70N666E215inxzwqCkNiJxCvPgvOGY2ag8qwHENgCHhCc6j7RBOIa4zAl28hSbJ9
MLnbRQ4OaQq1b3W/s3e5GK7yAgGykaHlba6DvnLs8c0J71vsbxS/bg9Nhx8DVjHDraTmomHFTH2p
yaHnZTpP8AXJo+SwRO991tlseA9tVAZkR+xs3oPZa3bQue+QXbNdgbKhekyCdu+NNNvvrxYWpbfJ
R9qZ/U8qIuq5PV49GrJUHdYByJVrdZYAYhxrPRbXx1T/nvk4f1k4/cPWIg81dLda4x6+o6zyqdYD
MnTHAPyn+z0ZlOlqDv/AzUHfUMO4MqUD/PFC88PE6uFtrnAS+f+N41UOUogclZX+e2JPlNZY/L3/
kg7Ox93IuI056xz8sfU56Au/mI066Mn1HRi7lPW7UiehUpxJ1UopOGGG0HbJEDDMrONvPKQfRAyG
t0RghA2vXdaTZFCi6EzV/IcoeSX8MNwplj46yMuxdaGezdzTiOajA+Myxm7/s+/Q3i7GzBYDw+TZ
t684bjX+0sue0yZ88ss5/drQIeYn14iBdp6Mx3NKjGbT9awu0g84PQLsDm+RvYRZjT7wPf2Lv7Rp
msB9uuRcnAzj6rY7V8gmacqYOL3STY4EaNWgzkoF3vynO7LOeOlDLJ2X66eCodT5vt413Mvx899c
lfQPO9OZGjQp4X6RY+iZBKGTPBgsk2Q1UCWXtJZpw0y/YLj2uZm4qBd/fIyN3Xia2NrkkeyzY050
tcglVnI5ibGlmk0mU7nNsp79As8dAyZ6wc8ZtbAHWC4GTrzLgOCReHtywt8imo5P90UDpMSF12Ci
Grc6OGJTO6yUfRnzC0THCmkgkS26ubZii+5ivBHrO9ey2znSqGJwvE89yhE/z8KYk7b8IIjBJSDD
sbvwZ509+Gg1jQnRUINDjw5zzYqmGjQDghwwCvCIeReNBJ4AvwIMblQg7liWQwcafCYHSzFnByPE
zKKEolOgCwLhdAdFWviQ5avW8PnzTV1G8SfhTZAevKxT+a6BzFHW9GPI/qWabAAHcLu3TpkWy86N
AL11F4e+4jGKbpgGPROuEeXyou32F5HlsJwruRsLLzs4f563qAVJBtugQ0YnUlaCsvQdzu2yx9HV
ixLG7ZU1IDPhwBmnqnJ8ja/XZSVnzwV5uP7WM50PS3+JB/Vl9PhZSDiVhrGU3RMpSs4A1YQabqwL
bcuE55lE0xeEtHBGMXsyLBj4VX45m1byfqsJ6mQj5wnunq/ySo4rRkzMBOA7ByfqZUX/tV7yYyhB
1BUvX9ijcALw5ecO+cR6E2/5Xj+SuNm4kaaSuWwwBBsZBe4xF9c9C6U54QeL3htJa3AjCUA6kEri
1JmjtvTa2TJuCCOIKSDx1Ejmyyd2CREXL+1qL4tETaHvvWYHW4Y1lttT+d6prZjbFLOinSOnfZRl
DwjhRHYCEXtaRDL8z8WEqBKJbIb73gGNT3thvY64jI6wgaXYCiQIhJD5enOuSYroGex6jLPU82do
xsjt/HceB/xfuBcF0VXXI/HyfP/4i/81cN884BbjUAuoxDwe/rVAuBUi+P3pIf2kdyJ9nR8TSDD+
/MczQh+A7ChjilB0Xzjl6F9S3Pz0U+qcQ9fbrrSub7IVeb6jbY+5ZKJ2s7z2wZMpqX1+f4niUqqN
+bmqsHJBzpR2ko6+IssnA48uEJIvecJgtLsuzvQ3ANJoc2MxrXpbHiq0YZWBPNDv1AJ2B6A6IZh4
m+SwGW4gELfg129L+7vy0xhXjLbMCSKniMdI9rsCffPUkZWSpeEHfn0Iosc3szY5PjLG8bMK6oa9
RayAAGLRLeg4atN6kfpj2wBddK8Da9Jw1RPbDNDT0Ki7/pYyYOUgfCUfCRbQq3fwYi0df/VIZhtF
x571pA0lVZTby7Lxh5p7hzTFRhSElAaNFQv1Hhzs+iPTUCghs92vCDsbicz4bNg0f8NERFJBGS++
EOKXHjPsE491RKL6uc4SBvAIAPhVhnzkp6biY+Ptg4xkeZV56073ihV9x//wIvBQQp1Kuj9HPRtZ
wh2ceZ6AjdPLMGkwOGtpnmDSx1UiwSz6sMEyqHhPA5WUavge0WHTOXiC5Xj2OBhPMUpAzLitSws/
xKxY+KTZ1CbEIZqOfz2YxK0nfk1vGG1gBaFuaYFuoDUhsdr54ZFOy8bujefv2X3s7eJhFrlxD4/s
U7/NBVNY0Osi/xOPNHm9agqFiQLlsSn4X4A9Vt/UKSQ2YXb8Y1FRQYVi0mqb94eOA4bGi7URa9Ar
nycs/XDLi1sBlGp8F4ecRq/2QvxNBJZn9ko1MVeVjJxm3LYc18+9kGL7oWud7YqW8I/tKRhsG4Jx
AuGwwVMVyir7S9nx/C2V6+ySpNMxt0FAQ4DNQ/Px5qT26jO+FVmRSwlWdB3ZQl3WDlDDVjBV/i9B
gECJNZBYrLzhEHY2NZP3b+KmQb2WsUxHRBMgXdwbxGIjxT+zJd5aMk6sVf3zLCXI4kIcWD72aJPs
DEedTMmqsU5LKccovVl29874ktS5A6A83fHjbdeVhOHa63n4Q7n9efKAFS+Uj+Y3bXupSxC9XaXB
3ZtQS7XbX8lwTbv/jhITO54X/iVrH7cNx/SDuB7AS+juNvZy3TiRTU81kJUjJ0ve6sipbb/6XXo3
As218U5gf9/2VOJiQtGujYbWrGTpk9ao5YPmAkJE0xMyWeDUOfuOd3ss6QBG2I1Z9w6ZnWPI4sDz
rZWZFsukGv2V8CjCIfn7hCNRNZEKo7a2/nLBHB5WIBgkZKhpJ88uHACHl/NOJkKBQDAagUteF/i8
k/fl8Oc5zVBc2gVwROOEa0tPDVfQQ+mYXZY7yCAPZdPSesr9jENRjvmk76hmX/SztT9MYsbhHOG3
gyytsUgswmYtDPhqbIc70tFaXwTBN2F8EHp71WlNN904LA+yTYUz1iTdI0Ww+eF8TanVBJ0Wl/za
bZaCkVaUHgJVAdrPypssVL+dX5GnVUA7P539Kv/ODhFoEosBy4/Tz//LwCmoC9BuXk6ZM1EMFIU2
WbV68bFS6RP4U1TMT5/K8NYtD25lATOnAMLvgbi+YMtUTpMyq77/67dvfeoraR0qpunHAvOYXRXE
CRrpBwPjuKBMsnrOoTqcsUqUFuVGi22Pp9vtfnTY1t3sNesp3YeY9HFj2o03yecpVgPUOaR1g/8w
RXwpcOz2jne7a4FrKQMMfAXp9bAKd4fQW/MYuIVb/A3XenqWrDQsByxC590ncs0MPIpE7P2KqA/2
4fr6thNbBCSIlGzQ4cjn2UtJTGp0mn8wELr50bTP0VKLYgzchcQ6wN3DeB3Sah7NmwhoJTRU+dmd
fu+ohB8SLOs/xLTP8C4IiLrubq+q2hScNCiOfyR7EfNCG8ffjDUyTBJO7fw/anSNISSZITHfTp7+
baDidf5HwZZHzCOSSYecwC7YJ4NgVgHUxOE1frYImdss2CedH69RJkdFwtiEtEI6c1f+7F8VQn3e
vgJ7b4uJOai1QlQWjCV4X3pxFYGH5qyecF6lMdpUeqouXltgHAOoZEm5mkZmzdvdAaEd40Ar99S+
bdGknJG8kMQmoG16qV806hivB2FSxtRvwtDUg82k3sr1N9xHxOiUEwNlHMEMwAWOGBB4yql3JdTD
mMaM5xvZjAhjJLRQVo2Oi/G489rLqlVdSDSHSW4vabI0MtG2Mu6ueh+uv7gdFbB3qfsYxuygqnmv
UvkyUZ5TgbDpUhJyXHsyi9jHa1kJImjvRz7h0EH1+IsfI2K00j9X0Ifmluij+jhBoM4LKWwmX5Rh
FPoJpDj+ruoNKb0h3yL2LvDf277gYYQOsWCX92IjkohoDJMAxsy4prl0YYukvh0AA8yLvrh3vgnG
nyxvdyNhD53R6i5n+Y2c+ML32aod+3T57aCSvs0O7lkSbCGu/0M4vuphTvvX37ZPM4SSS9mdaDjP
2xFhgezwS5iMK8wxeXQMjkBtcyhyTjkGitKf+2eKXamCDKJMYByeYmCk55psr76cUdSblALRIYxF
zTQER5GQoxfuzPAwsfBU/PGhXqHG+vWiF6cAJdIvWUdS18c/WYoaldIG340dCTVzn/LSo0w6V7U5
i7R3D2lUAv6tJU9pyJx/yBxh6hytJqGQVeYmwlYPOqX74MiH36hQ+KK3QAImy6VO6fAFJD1FSSH0
syD++dcEoWTjAQHGzx7kdh2m2NojPsicP7I0gSm7/0SNrXd29hhyJhH5QHDZ1zFMriw633vx7EoV
jR1ZWvKh3hUg0rUi2MA9BThsEfSRdYneTnsOnqTP+BOpS6C3GW2bqWMPwriMjZoZoM4WPD8uQPme
8s5dhwMUS5bqVfia0BuTugc7f2fN+8V9hsAm/RWFqKKNGZZ2i6c85nKmncdO/6lS4bHzLgpY7V9G
sj3uM8RWUpwShXec10xhsot1EmIDp2n5YZpHpj8roL3S2imfzp873DfSj3Jk5y6w4+7foK3ZKCoB
KI/sNO1ejqW1+To8iG2QoESt1YU1hPZpM8yURYDZH07x7Mq192kk8kD+rpdk2kFN+Z8usvvYkESb
VKbMZ+YY/E80SrD8+akCive9wJkSjUi/INTSsA8E+DQnWjcMqRdoqzc8psWZdS1FjAAfVLqBFQo8
mW63TiHXgMfFR0KaloLWDaDE6FTElxgK2ysWynth9B3n77E1UgjVN01E4F1pKgyjpf3dAmRFDBeu
llVNqsS4EOjNIwMXv2efmfkYbs+xogaqk+1GFU6VFqKeczJQNq4Y+NlMWtjhjuJixp+p8uLF4PAY
hhcNsppiUYxz55odhSVCTCH0Rr0Q+Mc3sDw7xPGkEMjH9kGwgB3i6PgkuAbOmcR/HIbKX+751t/R
nWD9ZTYOtKZ3FPxizaju38c9mnq+AD1I+sjmxatTKOVQMWT2R/VmkqCzPl+cjbXYbzmCNUUNfYdB
+hwR+LNtzAgbbeR/aZLAFZEoKiS3TXJw5l8evbJcuOZt0rbTvqMNQu8INWBLkOuSHPrE81qKiCXV
TEkDi7wMmLfrihWJsjaY4vOK69RTuxeSGScRqSDJvYNXvrb9kn3agmsrwjUtlhOI6H+UInHoivb1
B6S47oG9U6A8EFFCzhnA2UVCIRhTWS5tnWcWswVZtWG49WesEZasE5hBfFCfnF6SI/cZAXZ3xt4B
b8G3+lNjdeBEvcVqu5h9jQYSgJqL4cKhMCJI4qgf+CmUKOJSp9Vp3hklzFFRGjQFFNpUXs99hlLD
8MRpMF09vjCM/5AL7FObLtP1d8Epqa07Ta6AwbHFzEpZLriLIqC8VOZxCaqmv66IabcwB0CZV0d9
4eaz8VxWunnVylRKhtS+8gJ/yQVBNDZtTkGcXZ69A40UB1Ml5B7qJ08nRSyZVOq9JJ7fXeGy6E8m
5ugg/1SQedPTj9dybBekoH5w1vQI85znh24kvrFh7vs/mmufq/oJUF1kApc1+e7cA3OsqcIFvTGI
LINitwqjPRG5ZNNGXHlIg06XWXA8RGKtS/Cho8m71tu9MaCH2CWsFUTHhPd+XpZdY19Q9qQxCbpR
N4/nwMsGLjKrXnA5+IYfWjWX7EUbN03eKn2j9wyc7VA6E71xTEfrOSRxUGIe+HeAlr4TSn0YVh61
7zmjutiVaGLlItCmL6Ua8I0a5B9yehYQaWTKhgq6wuHE/WvVrlbi5sQwrLb9Po3w9wQFMbOhVXm5
Rt1RMceBDtb+vW/zLuOEBXZksRe1OVrAHZfMMfxZNH2uX5KjjsicTCbb+MCt7KT17tZmDR02MBzl
h6C1yC82S4NU4V/PbxKD2QXvw6S9Jrvn1axxO93T+GI5ettFjAbAD1Uh5DOYbRNMDRJwPkJJE0BT
cHd3AmHHb8PmbJvC4JgkDtwuMHru8oQoOinRVA1bF/erBkZCfaZBTIlrJ0PviLrlBz5cZrDZno5O
/Etm/yi0mB63xYoei9hicOkcjTaloGMuWzlPLsKQb6R4128aVeE0CmRB4OQocS+DSAREdycBOaYD
Bypp74q1qKD8fg0og5ZtqGZoWk2bv9WLER5/JQfDxMdkuBrRgwpeLRES1LH6XCXk6eozrmKNeH1g
7Kampabxoy5KwDYgACjaSIJFKSt9fU4okCcBXaubl7JQYhDHRnMakikQtUSUTswFLqmr7iaAKFq/
KoqnCUgdrLaqfBr/4P5cf3eOuznnOBJK85zxNPeodJm6gQfCcH5yb4zVde2wcq79jNXrQQ6Xmo+g
lm39Gd91hSN9i9EZMQYoJlHKPahcfrOnEEOk38Bu8rEp4cyk8tB/UQqqChDYhJIjW4ncZ+izZEiO
13pLV47OA+ZoRRNFwQACFEB1p/CFmrD7oR0gUl0gVWFZuaWzKw5rT0VKCRsAPqPyX1gw0bHXHWCW
fzFCDjgcEasvHzoR9H6a8NtbA5T7KSJ0tAXqjAbCSZWPSuvOtZun6w2ybI1s5t9AOuVqKYWl3ejz
1+i4rt6ySaS10xnChWRZD84RvZDPg95VmLj/lKNQHHuRgadzQCRXqQUo7qWTPR5z9VzMPqeo0I0N
4Mrrj42jWk3BulWAEVWF8sgKrdliBufjh1iDf13j8fKVEhfJNjiXZ5WZgUBEyDurMw+1G4vpkyAL
3lgTEeL2NLKJtOFpHf7SFzuJOXvjANw9tvXHYo42w0wykFu95mUoGoZX0z2rMDnkzxbVIXz3wdrB
h9lYJ9Fy6RD4vPyutAfvLDK44T6/OKk2b1zJ6ijII9xJWm6FusizyFN4EvRESXSfLswYwzOuYSWc
R6JpwdeMayeeS6b4d9kLg+XsLyYy6DCoGviiUuYTtF9vmbpvIRGnzjG96JIEWi7JFsSR9HW992di
91nYC0VLznEbxxS6nl6KXCpUCUpAGR4u1N46M6WYIcUIwY2Whu/OlBMwG7zuEF9y0+cJHPPaoWtO
lJ6+xDWz9YefGPT2JkbavfBR9P6gc6BZb+HDvvtoq6KbI/huKuscZ4mrnfYmNLwkX13ncoqExEmB
wprV9zBu9ycOP9HDTBWTReln2whNn40ZYaUNBzRsR8jqM+wQz4ETfPoTCjCfcjelUl+ENBNJKGzN
+MsqT8+Xkj8WZWitbT3dWDoLy+tHohoAKaj4wMDucqV4aiB5vDV1ndbFTovsbwyRtMgSq6Zfd0ab
NZ6Sa9zDMl5ttXAyHiCHAfNIAdaQW5JpniTdxJZghKPDBN3g8l72UI8gczI/93w1TahHWEMy68fe
o3sfY2cSMag/+Bj9ieh81iDl9QEC52ZbnnRMSnrC5KfOjWOFKBmy+U0CF3Tf6iTFJ+B2BvV3lqal
ltQLhin63UTPyxZ3QOCtx0WPMBEVMZ85LvxUH9CJ+OTNmjUgKP5KBCZ2TKqlvQIV7o2eBpRQRfiN
U3mt/VyOBrZe3QBYJd+BQHXKjkceLpkTAe4dALnYop2toHAcwwfPZijdLHfiqavZW6wD0yVcyNgG
ccX8hgC29pN3EvTEy4OCqxHLElG3eVKnMQmwGTZrqlday1f79LRNxlo8sUsQpNESc4zHjMWwdRGA
+QG4p39EFTTBrsfdNFr/3vv/vQWQrK5P3RLBXqmSZOJxhm2shahxEYr45fUIm9/DsX5JpQCFTdOC
kv69pIrVAbrPAT+NLxyNkjaoe/ev6bh79MqMVYSZJVi9SBANU4Evarr7b7tPBdZ3dqzwAvHPFRqo
tC2sx0wNhWUJJiGUsc5/AxWdv/Y0tuh9aKfhNxC6gw3ZIJqAj4p1IbmaN0BF/JZhnHjlgNPV1ZHP
3R91Nwe2zt3/1khIWDeRH1vYUFlPYqGk0BGCgrURW5O8PiJMmgJCANpC/4wzBq/EonrBeR3Kc2BV
HubqvUsZjWD4i4pZHvROTRbwnqIyXKX16AvQQ0NfBT6S3LZB1mf2bmYeC/OsnWHQN8lW9WdFX0XL
xFTX3zbyRcPfWAmKjxObu+ITtnNU7t/jENvgtEm/n3KUoTFEm083h1PsctTF2fY7baL9efQhuZPQ
/cEn5LpdIb8XphT31uD/qF11kytLx6KSRnLOZqGN/q5U6ztkkHUaKCxs2+HF+PBRknF3k5dW6aQU
K0Fp22V0hM0iLZyG1O77o0ntDMReJqeh7yj7XDzhlkEIHsOW018+5EDRnixLXQIsx3rjWMtCQfOd
KuxM0GfPsR58Bc84yLzuPOtIeNkoXz6OrFsDeVtsAcP/mxtD2gmNGaw41frRTaih2/IIu2tFlkY2
QAZCJkbv+xoGSDmr1PnTEHzsM/apyIxjha6S1jwlcaR8ylSNO7Rp/ZyPPUb1BLaABs6ggyL6cABW
NKFhTsSO+f33vOvDVcj+o2nbmI3ZvkTVFnNvL1pO8k931h+b8bJcunL6B8UltAe0SV+BYGcmgIBa
l7zOgQoscAlXe+6ExfBBOQrh8mknBVOgDzukbWn2LKwftsYyqboaiNGE2qM8o2DLgDnDDN2HHYEJ
Bq9HCvx+Xu+whJWVhi6RN9gZldtzmXwOrAHD/Iq/bwnv4mhQ2ou515rarGmIBexYAXtaYSV4yROG
NzuAVIgnJJ1a9Bp4C7YkTS7MfPgM6RGXX7ZbQvSwQ0q6R4Int3Kc0nlAgPuPC/rg9viwOieMpVvR
CcvyWw3Ooq9j5HPBPGG3lydBSjdCEJpT2mbcA2alP43xUyOqy7gXEmciC6uVk+3fVb6jqSz1OQH2
oiWwJpsMNW7oYfHGQTeUYLr9PgT28z/T96mKsrVXmwM/2QA5+bUqFnDkyeNCsobBzO7qBH1sefLP
Svlnl7HzmcmUFMc72DE/+8gSuX4guOqxj+aBtXdxWchqh9oq6CI2zybwxFYYWeob+5PoRfSOGgy6
TmdNKYdRlBeF48UjixKO/V/MBCoQJRUEzi8g4mePxcFbU71Cx/pINr0RAiGfGgOtwZHsPvrCs2YU
hlCPa+0AAr8SAuLay7XoC4Mj9gBY6CrW2LBGpu3vSKwMZGSGLHnFsbq8cD4RvuA79bPCoGBCAQu2
Fz1d/QcrL1pXbK/ihnIMy0MG2AObz8iDvFydP2eWQSIYomyyNxNbhOI4+FFpXToMtEK/Fz/8f99b
ZEo0ky0usjcVGnCHDT8dGFPzYjYaLru0Odop+Xtf0tk1ujEMqCzBsy0x95LTGfgPGoXKaqHt1+pj
yOCyYiOiqaagzad7BdtB/qsizEfEwBDGfz5xTlJjAmhDmoTTV7lARISP4yST5JvrIoV/lRoEsqbr
nI10s9ab/fShQ7QrPM00QThEzKd2pZ1mHOri1ujZVu8aVKlx+vjFdP6EI5vsTCT+XyTMsXKfNnCd
0WNQ0z/DGpwLFzL3rlfzMdNeL2IcReb57tyT9+vx6OM1e3cQeB3XlwjlFQU2QqOJbaZkAu4fmwLm
WoRxovnrZgQJxBx1fuQmGCFs5hDaQ4eB4v4+RQnR5o/euLKCsWcwQZBPT99E+UhO8XYzmi+V/nX9
eUgnFrK3K2H1MXl7yYL2FopPYUNR/pU7HT7kk6oaKqyLYrMGB0l8nE20N01GDiTkQYxmNdHGxcRB
XieNDYTif7Vl/JBQX84+7j9ff001ZBj3853nulsRv//F7lkFXVGrtvs3n0HF4qoU5pwGWNZUnxYa
PUnqvgJw10WSQ22v4KaKw622TA4A0TGzdf/YkhXIt2zfAXHJe8nOALhTCNoZ7dRNA6LzZDPqNn9G
Q0iS43OoTo6fuCvlaWdFKpxVdNJ3qVJbJcs6nhpfqEMVZZjshXlQZ8ZKCzypsPToFPV/6JQL6PNX
eTa7dGS75vTjvHB5PrfiDnBaV25n6VFnngPoZme9BFPg4Q0W/wE5jL6QbllldlmodJklgE16boBn
ouxQib30MFLBANt/Q1sqQJfbq/MNuyVR4SJKQ6ooh3tqcN1z2XuYPuIqkqcrGNvQb+Ys3aTkoozP
PwobaZIDS6vAol2hQCcrzlfhFVfXAcoIdjIhZqFLBnB3czipoDEwbZOMpOEUtmFdTEUGk2Cy3HZP
avxL2AKpT2JfsZIxC/vNGOXeBty65NHd0v2mncLHrZ3Krx4Z7dMpgxAut1ZOnmxR+Ut6+EufyjI7
RPM75DGCjJ/2ubyf6JEp4Wyd3OI8QFd0h1c803BfJDDnU83KpVlE+eFVN89CUh5FDjVHjlTbpxy8
ImDR/t+2yZcUmer+s9aU2JRxIMYBdqVGubRvPACKE0DMP8iPplKQYUYhoB8JHqz3j3GqWIDZLMPD
YqquubaPuXO439lBLsTQYeMGZvWl38wtuPOcEbHwQ7RvDdZgQbXCygi9diZ3TdeQRIRngv9G5xAv
TIsVVVILBK+D4HAIeG/OAIMsFBe2LFmhUAf1k9sR65oTh8W9yZMc56OdV2H2F26Wz8DTVeKWB+e0
bMYVYYpRyx+Q292QhcG/Pc+xZEF6Aq61bqO8Cvoc3XHwXwA3kB6xBjmmMeSDCUFlXyNSh17hicpw
qkULqcRDGeDjxu9rAZmyyeXiDcvD13drTEat/pfz0O3JBIZSVQNFIxHsW8dNFpDCSzSoaqiPatVD
hAfqQTdorjPnuMrkUSoZF0ptPs/HLCan4evCxoU34JpNacgNZ6+kjVvUh81F27aP1E8N6AxouZYI
IaFAp+FQw7WAfP6PM/7l4pFTR3DNC8g84ElokCsh6/NRVM29f0vZr33PRU++X3suGk2RbWsZd7yB
tkW4WT5+7EgMIWgcrna3Mh6dAlO3W1XAvMlazkknUtoqJrkt9B7+pU7KFLEMYBObZb0Do/egJPhs
qVDhRtgZ79QVkGOyNlxq3QFSn2NGGyxRIpmpzhKUTBKwzEvY8hZIZnd0YHb1Agrz55hpCUxIpcrK
wyz+8QHg6bS7gSUwAiYvhRBkfZBN10W3jFOTgqAw/HJ9iBWG0dwBkIzdD8ycKHs+mY+V5GSjF5+0
fhgrpZ+gr8t1renmC4vObq+Lv3KT2xyaLJCHvHw4CxjPxZAygDVhU2xTYAXSMM6XStazYaILBGiS
Zq99ANDIbAkMPPoR0p4u2JkSzRbUrSpH4kDtRxYzVUMIXGJ2bkvSW70LShZNSpdKtjPNmlFl5W7R
IYVMKjR1MVGNiHFonv6jAReiu6j2/oCnlvT3xlHAzExlRRHySN8NNxnF9mrP9oDKtQVsqUhTIPyL
jKnV0s49VueyQjg6Y9oQQwZkrbUjY+sLWHQni84Y7vOraCMZtvorODsxJWLSIpVx6TIUSToNIYaP
7GY0svKmCKf3blNPscmykNO9Ue2xUOrhgnhMrQP0N0ZbqNzLbAXjARaA+9sf/AvbdQpHX90KZ5dh
V04TnWR1TBwX1wa5fR7Orqht1rC234j0c1poKTV4IW+VsuWW4CjCD2/3F0fCph0U+2PM5acl0QDU
dOPt6FB1UVIVrE9PaApFTXOI++wpuKjIgbYm0w7oHAb4y0T0+MdNPziK2Df1f+jg2l+9H00mQWzZ
6tw4iGgWbfzgBWjiTu8D810XJLbJk3CvkwlhwvTle9fOqtAJ+KHfuX9S3w1q4ARBIzlBHxunmq5c
zaTdxtnE6viGg4W0zIqggZT9pT3eVcWGEZRVlm8DyedOHR8Hu2YQgqQlmzItdlkcF9llGokX9edq
tlrkIjmDLY7ggFH0d7EFbeCQE81XL4vuMjLLy70l7iN2iqYFTiNyruVgRvRPgRlMmyCP4I7kF2UP
I2GuA+sU0m3Axe1F2zZkd4ZDW2/Lhy+vOefHl7lQaB4h2N5Z4/qca4CRDaASDzZXRk+E1bbFJLl3
7/M4d2ClEemphX7Jbnq6sA6fRLZFyVuuseBh9Blxf/MfgTVvEz2evT3L1388YMkEuPcxwrIRN9bv
3ga2IeP9QS6if9am4RnY4A0W56HO9BbH1YE9NauuoWX/Ul3pu3XuHWIp0ekC8ZW6URnDcHI7yHqy
aR5736llr+p5Y6kOe7W5ULEC2n4YHWQaJO9KnuSY9sLtHd55+eNgbo3dXlB4ZRdPt41uYUK5rqW2
okXysLj8OpToem56o88pMqeJ+A3KJFrEuk15I6UuYn/28fXmP+kJ5PMlZVQTSJv9FZtGSp6qzK0v
n5CzTsm5TmNw1VE9AXrrM6x7RuXx8rjwN6oOpl9sJ5C2B8K4QM+ZnT8xVQa5oHZcxyY3BL8XHjjl
57oYUgRillXeS13OQ+GUk9gZjjC9mQ9Ba0ERnv3VpmG+7TgcT/etVbdXpYeQYM75b4RLfWmn4cqg
n3J4d5PpWDJ2HibfNUAvxFRKZ2s+Ymf0yrvnWNOppzMVp9wWrHp2uudoyIW72y5eM0MmcMABJuQS
qyGndyNrbFRImAkI0SQFOCyGt0Y0St8hoYz5BaBc+RSYZ4nIm2cyKKWDc+Ao0QHrJC5/uEcy5Nta
NIghfMTuB5Nnr2UIBxy9plV5qD6TqOJqxFRKzDACmSNNBOq1SSqi4pXSyAWYZR8iSHXlfCnQmP6y
n9dnO04B9HdJUbSQse4oHCT6IVq+fK8rfmBVj2/NEk521q8QSgzN4QpoNA4VqMNLZsLMUs4Z3eF4
zdpfhQb1wMZGRsWcYTCTQdpeyJtGBU4hws7DZ8TByVWrX+QR6mjR6nVs2gj5G1YMitafDK7eZD5C
Mz+Ynq96JeULqklgN8v51gOlRIF1hDAN0IHdbPtH7gUs4TQjVmRX2UHAq8xDy7ocNvPhV1haOZQG
3chWHrDOCHStxXE2DgmexcDGiCPpkI+qJToxKJtbZB3p5PTv56GUzFK+Sb90DAoTFdj5+9afOHLQ
T5l9zDWAPdYS1PfHdpi8TZeYNfMgORp05w08NQh8wQDAUqWVv3OfBsCFNMfL6EMRbaJb+2fxbu6r
GKbOOdfBxm+PcYQAbV1QpGdFFfb7m2W9V49MNNj3YXZIhd1zscV72Xf9t7Te5hwQM2qOg3hKaX+K
ODtY+6clKq3FCIlsKem8G2btJutn59soYsw6lr0Jz/iVjB0Ji8u6SKhIaW8kRKQhUgIh6UXjTzwx
SkECbWrKW4R65LYAZ/3F5rJ+qAKSJgw5dtNQ5dYG/JDNcxBzHO/iPn9et3hMkRQD+F4Q6PmHu3A/
0ihtVFrqXkWLhzp0Dkea9O/pPFmZed0eRJYdesj0WN45U1Ot4Y+ryPCQQM5i1Mb/QfLbXGlvuoul
K9Ofq7OYwXjHkih95JO1AvKTmS7evXmCRbVub/WoSYf7QaalxQtUNhrRlpollT6b406P3cHqV889
Y8V2MYQVnOJ1UgSvxr0nex9XTumWPlWnozbnfA8ikhUpTnEW9P9dXkmgeXSv5CPlvAowoUhXIqu8
nzMF1pdTrvV7g262bSnM6glJBLeYXYXMqkWXbC18pcPYdbcjGaEgrj7bpbRJ7qW0aks/zRKOtVME
PDME25ubPJkSOSwl4GZue4JDFTkLB9moRro0aK3EAdzm7+MtIW5+dFcmFl5MK4tRogwjXtgCHAss
xRv2pDf690g6syvMTJwHVk4hcrCuuy6emhhIy54r+pFB9GvRm4Suw3NWp0zCF+8G+fWx6AnwoDip
MaoneATkwm2ZeaW9XCuLemihOaOreq4E2NlPTGbYXdmd/KFSouS1o+ANFlCog9rs3zYPqElGiz6H
nQlYCKLGNBuZI7Zv2vTIxZW8dyaGWIcJTwVw5lbdhLQhAOGDhvdeybgWV4w6Sg6KtR8H0YIxc9Ml
CFWRGfpQhWLQJWU49mYe8Klk4xiQnYfUV/xiOhrENDYQrynB3q7kT/YvEbjWGnSS7xlTHULMRkHM
eVpCqKVXBLpUcofJJ4vx8neJit6Htc/xz7xN7B09ErfgIOoaeiD5D4S0QE32XQh81z8V7klCXdl0
bkuJuC8H63il9RN0ORkSdziqRT8d0fuvj79RFrLre53DfOA9LkBAUdPaNd+Fsl3b4Y3gQ2ah+wNv
fTBeDvjjxPFBR4cJXbGS9TsKFEuMZYeFOAeLD7V4xsJywxS4xX1zsi2DbbXf0qz96olJRCX6+xZM
JEfA+BvmjvGqnPy1/EIiqV4mKMSopRfzHnwb1JHhK0c5JCoNHO/GAUsW3dQ+khUBcUzY3OTdvrZL
zon03JJbpuic5pnUezH/a4pzba8KdYbCrd7BdgxRras/aoFkJOHJgiLsaY+Ebn6tCI9+sSC6xbsp
yTJkOhe8wAhSzPsMS7IJZ0hVsMvDzeCg6bDUOarLjQinUoEi733Bwfa8qLjz7k/BH5TXVx8XAL3k
+Kgo4b+Obsjc+njSUgfI3nXD1KPU03WQ6JJLRIQdYRZK2/8lJk00SajpBP62LmobBFbFR3oXSCDo
S1wMxgJ1yCUS2GVnQNLTXuUyg7bOzPCOi8f8tzAlJSgME4TCfPlkUHacNn62uR67j9/qDhJRv85a
PkCCwVV5UeeMpfmZZFPwwWCHWdcNEVWJDEKfkM6TWE/ZBsAGrUg1oI83D/Crt0jsj4He9M7TopJV
L5kYaxNh0UuyjPXUBzGh5XRnXrekc/nbUeknXhxxMdVXvJQdCg8cSR5CV9fSeWYMvYeCSZeNnZIn
NtqxsgV9Qo26aVydGhbDs/WXEAOZyB9Zbpxakt22Yq6a4SsCbO4uMjy0PcL94268+wNCUxXK8TT1
DYDQAdn+j1PSKmM6XjKT4+cGI4eB4mopAJZDbGhlLPaP+ykTzHv4ZowlbZ1P2NLqaOa4jtaBDa4I
GESoSQ69Z+IGQ/f/FmW/jXTOtifIPIBjsZXbaddBuuHAaJzktF+jHdrcUyFsUVf8b98QkBzNKTCT
gqpaEl/xwndkyu2zkd5vxLVHQ6lNxo7rSCCHhcE3TbaDJhMCcryIpDIctCBbRKjVIMS+2JHhwBV2
pVbtuqbPh+l3jBzwoTjSdMs5h5NdM2xCoLGC8yTrTfQguqn1JbGhisKpH4r+k3c7p4rClCcXqrl/
Pz+3GtC1pawmiw1IBtc0OkjPbeo13ee93+Yq7+sNy3yBo2yM2dyO9XqtoIYRD5T3ohazVtQHdOBN
UZxWSpSt9BWKSnORYSAbQPghmZCIFXCgtWbuuGX8dPOCw4Sp04gy1s3yMkHELtCSE+79vp4vfbCm
DP9CiVeiMTYvl0ousNoHJcQjrawAH2lR+buDJPJ+ySfoN+F4hvogFz6VCIcwAlh74oDNjCjvlEwt
0s4098R67dL+/9y/82X5dznDeApzavPU9vQvsYI8PYJUbSkPOKkg1SKNOzwhq49NhWKGnSzxOmwB
LuLguQ/mZsHziQpZTC4NPKcWVl5ApQG+6xfEs+ycqTi4T+QEbrNdpVu8r1f9+k5JkiJkiGjHN+52
pKc9sQz9TK0dNSv/tYtrDW+1I6qniHfh6zS2gunnTxbuzWcpZ0tPdTAYpBOX8xIsuwySxMCb4SZA
I2AJt3shRZxTT5b6KSzq4lWfVN+CSFBq1N2QL9IvdVasnMrV4cabmuMbhCWlWkzCwk6DdAIXuZBR
IufCUS7TNbwdmhBxzI4ySJNL+kzdujhZpnKXWBVIh5nMNYKhImw4Ks/FGCTpkSLkReSHUtBR0Z0j
E0ISfKJS77KL1z4FVAmCywPAJ3fv7pUkb9WtymPblZppTF4I56+hHZWxeLcLT8+p45a7m/i3kldL
XGzuC5hJUqlSB/NSgDD0EJtfseOw5MOfqs/Ll902Pbf+psPjjunHJsCGyZDAk5Xnm5UbyIFrU5T2
zF7Cda3MudhoxtFhst6Z5Xjd1ym9ijCVYuJ8TpByKV7GU4OSWyRmWu21ZLB/DByC0OwKIy+n/lNb
BfRa0e47FlP1c86vn2lvKe2c4SLNlvzfC9e5PG/MDjSgbc7vo54r3+cwhEjo+cTujrptdxR4gIgE
GT22bAyP7zIOjK4FLYmgrNMyNbEx6xdIqm4ctPulZKW9oY002QLFa10PYxQ0W3aII9p4VPa2hIga
XpwJdeTeZMIxfy5gmnCUGu7z0cYk2W7cG9byAOiGP+PZg0KMcIh3wX/nrMRoDlTOmS1+PX1caB3C
ZcW7lTXCnQMtlKUJhH6NzCOab6BWXPvTO87tBdcWunUPkvuv5H865S9xdtNGw4lD0+H1fkr+86gk
E2V+bZw455IErxlAUgRFFi4+o+bSjnbJo5G6RZ/uedoKqY5l+gdur6N33UxOVG4i9KPldARpswLB
8nOyPGwJUSbfR3OsdRddwrfQc36VwA3sTYsZhhEuVx/pMEwLjUGtRgKMb9oSuykQkdR+Tn5gmJC8
bG/Lmihnl/5iI41C9hPJsyo9y6tUQYk6AFATWUZjdn/bQQ5MjVWp2wXN+BxVHfx0pQtdQzRbppoN
oY8tR14Vrl1wrMNPoNeLp8CRh3C+blRXuLdWFKOyd0Bxisa0+YzlV4aPtR4pE7bD1qIWODuVqUxU
L/Rb/TtLGFimXJquYtMbbHM6NG0Qn2UVDqOxzTGOlE3pi89sKyxeEPYziPvNMVXuvfVL1sFHIhq5
/5/C9GFYDhr8kharpCMi/QOumxW5eSJ4AirUV9YbDvOV8XRWV6XzD5GHOxnqHaobBuPuH3ZZ3VkQ
OXFE/SBUH5nKUNkmZdyZgJdOOaFvZq/fQqaZ5+wXPDlJW41oJrux7BLh1ij6ikJjOKTfZ4YTAswB
Sjlb3j1ii2Jta4nmGTGfcnKVfW6EYVHyWd8/+CZgxUDAJy9dI7OwpyGvoW1Bx5kFR6sBMHD0rydB
h98cxeO7iv5rjU4vb5M2/TkKB/e/lyH96Auow29jGQN+DWIZp+mc9jSYOaYPR8fgdZknvwjFU4j7
c0csVVJ1F/2cwjcjFe+fUw0bbbaLQQvvas8JAdwmdFiwSXtZqWrT7KtIJt0u/N8AJnwm9R226NfN
EmuWdEkDqrKXsDQqDOxHlc2RfQSsvPNxDnulnmsrMxYRyX/zdR1VYn7v0fqfiShRBpYcCgp4KXKT
RD09xPKnMRiwS/NbkWEO8/wtqdlsK3tSIYfF1kgJ6wX3wnYjgqGpw6jLemN4T0BZsp7YY/Xo069Q
hoFBF5PSmi7lFf4Ejgm5kg0A4/mhfdIe2O5DEQ3UlZdjf8jfTWlXiNlZ+tYCayPIrYPGgRI6s/0E
DM+ZcKeS9TRpriNCHEYuc4CdX9i++6zOwWZDNQdiZp7MlRXECOiIAJiMKrN25MG9i3ZB1BNYHc4F
z1XFFaJ4IkPaaTZfhviD3TgLWUeHF2SVHpu+5eU+Xk6i2PyTxEx9ZphIh7Gr/GkRz4HXnfQUquZj
k4X0O3cfKgOCc4Prq6o3foUaCJfVkiRq7as81RXxrxTVd5wmgPrLTTWuWuq9QE+cjdmh049nSTJY
N1TS1W2Ux4Cwg3eACVQrEuTTxrIBukP4PUkdp+grPJ4Qpu7u+qxXValTuSnurERp2GXdAzeIbqY2
GCaKclklg4xYUjeEMd75KOwgoY3/n/zuffjuTWA1ux16LlMjtHpC2sANnwKKc0D447oX+gk3cnVt
q6jb/HVBcF9Rm0POqghVSQgkqN5gelduyQmlIxPufPncy6Z06YrKKArfFp/Or6lnHqXa70GXaZ6k
PkLUiSVz03qaU05hRKiFnvB+hj8TQUQgpjyKELfN69CSJoS5x8RnuPSIHz4ivXFDivBElg5DVgxg
qyZQsK90FWwZikZXoosp0DDUmQO+yY+65Dm1ZI8LbSz24Lh0bsTZClGflD0+TnHhY/ZB3+pVVEwN
JsycbB7FPKWUoHjcBlDhHHYycfQR4uJD4XtEbJ/MD6GrXDNOsTRpGdcw8YIYiO+DXTeSNq0FV8KF
TUrPmXJb7oVelSMAmx4tUbdy73WW9rrCyti97VfEg7yTGn+lWW5ZHZ4iLPdxiuEHugCPetkIZ8LF
wrpTFZfT0J4/r8cY2WDvFqLNeoxOSMyqB9Jfh0XK6wV/3jBC8pJO4mcE+E7OOPdaSlm3PyIL6Sg3
8wZlHvnkHghaJvqOBPqltY/LsDYsSRmXCTdW7Rm2q/NLZpoanSRUT9LN1V9wkY/Ru1ABQxEpR5PS
4DWj/XVYHDw/3nyo2N1j8Sf7MUft6/1mifxgkXe1yiyzz95n10UlM6pIsGEdIZk5CEd9gWoYAwdv
Uj8OiR0w8FkGv6LH4nuMEdveSFvC2+WwqiF/JGTUNAHgaK7XXTHuTKcSiJklDmJOxObNopJbH2wl
0sxC7mjLCysCqBBR8FwZVuRdwQrF2dGeT/KTqJecWE/d5dxXpycZ6IAL7wJtn94g1NAl/gGiwT5M
5VCwecYjp68zhwTTA9M9fsgNTW3+zB96rHKCRJ47HtMtkGArFPuauVJ59ETp1PjhAGDrKmSMETV2
xmxG6CbuP3wjk01gIY7KkZLBoxfBtThCww4wMwJ/nyN5kwbErIFlnUs9Q66qlTJ7IKtuOMdF/ctQ
0KqSaS577Ti1mRsdORhQuYZbWsbGlKkuLfIte+LzkP8140fSfn46Ip7rPrCbhug32yMSelBLl30V
+5uctkn2w3tALLvUb6YyeJWf+vf/cr+W5ilyXu9BM3fSsxYKjT70XyNumGQFzUnT74EeUbeFd/7z
tb1sRQrtU0MtBDNavcCR6RnKoR0nlXGtANjXAnmYncOg39LPCuEVAObdstGk3UREv8M0Sx8XePQc
D+HdmUmkcshKM6ypgh5PaSjdK/L+39CAJuK87cDOe1qzobop1IDxEz00czlDMo0Z5QDgDm7sQOAD
pfzj4mP8P/hooyAzyJTLDnLc1RvmgxHz+OMSDzTuD6WI2Ae+CN5KK+8PwxdOTThETIdaGk0Y77MT
LL/zCEaoqxRzvuKjEIf3KDQvIp8GyEaCDaRAWJAeHrdNruixEyPzf0tfWhKf9gKFH5UXAbr1+ouY
VEqIzmb3OSCZMnWCr59LuC/Dsc2bxvj2+SAW0SdS+yASEiz/+ag5ZL7R79DzfcR6BKCnXnH8nGrq
j3PMXl+wJvPzmmV2saZywvBUYn/Xa8p1M4kuIUTp6kyGAMI4rv2Ue8q0cl7idkyecdKBIPeKO0NQ
lJteRvebpNaRuInNNYffqCcjAwV1RhqF37uBkTHAfsBrpFUeqeLSo4k1XQ5vowj3P7NqXl31QSII
rxedMsWR9FQA+BfcR/bRKIQPO7Jo/driSDCGhlaeO3bHoLew9dllo4jw4Fby26S1a0x99Hdc9DVZ
pO5pzGMaV3HlS18LsRgTbrvrs2tb/irU9HgaH4HzZnMPjBGbSH9z+a2FwHdisWzVv5yssSulOWmV
FvJ8WaLLvKemAazo/rwBEmTz6P+vPtDQerQz7/tFp0+2zQjDnhqoj92AmbQm6fQLPoIBLoD3hSxL
zztCbbgFcz1O6JPF4JB4Qefg1neTVKFUXo40Yd3sEIJINK0C7EweVUY7NjHKRQSdBh9WgOd2bs6C
+DIrWBx8o/Suxmb8e1kTSXUWF8DF19b6c6dT+rHnCi4GUo70dJ4j2XgACGZtnfbAgaBquIxiwNox
t9E8NLWr8SWJsfEsKVMT56aURO0Lm9gb1EJ3U0Kk2oaDNfOmjacr+voEXp8L2ZLChnAejUQ21HLi
zZrfw1U4zwCw2zwr2e4ALnup61NdD5uTNVvG3lf7BUHW8idhDR1CTIeuIvmyXONwQ1alj2ec8qRG
KJs9GI5R8kdNhoC+/uu1EoXWippxFUBZw/SiHxtpGtI1ICrsW8ZEao6b9bmddcyeVBxUGnFf9dj9
d8kM924JA3MWooJf8cbv42W98XmqQMWX2YdUOt4w4/E5S9f4skRxdxl53FRkQf3Cbjg8KYbJ+9sR
xT8Hsmh8N2EHEhjanE/7S+8kFRnOZONJyqtxab0fe/6toSvZDGtYkOKvSJH5xHXPl9/EjXrODJpw
GwdrswyluKkearWYPqy8iXAhpOnZxZwwC3Qu5/26vg2JU9qB2WzOh5zrGtQTOSNgqBqDONA3xxP/
/pU8IoviPwRp9aT4Djwg4TqY1iKc/4gdVh2ZD/xoTIXH6hOjxfZRYPskT7MS64h7Zt1O7ByIInjR
rN3ytKKS+At2qV/3/f/gJV2B5Y+pkJph52OLvBG6IFLVUQ5CkUI7QXZ/ry2pG+Vbsd7JksvTABiE
T6jgUw24E5sE4nRM1QES+qs7gd4Bprvwd8GLefuYbd4qANdKhRPUwZzQc2ulOdlNvq93tFmcnTh0
D2hQJaRqzEtSxEEXT59d2us0a5vsqAo/o+llfAEUFlUEIYX6KhEdaq7WtP8IuPxj0OZ7BCNrHk0P
Lvu50pREuT8CE9qbh+T4agNEFWB3dIyYhOvdtwAa36lKZ5IRJsm+Tz5ZScaQEy4IRftX4JFWPiuZ
UPNtd5zxSXVCJkGeqPxN17fME8ijbHYzE+2ljWKaLwR342TjLGPw+v9fZ3Smvgim/yTTNXjy/SBn
lU+6B/WLkAK9/sKxYxCCXzghxsUKZM7o6ND7fTvrYXgx+i84DD2xc1+t7uZJt15LoRJzAFd8CJ0l
XcZl2NySY9pmGFoPFTIZ6juuu25qWIip4ZONiRGvzndkNW0tPCirWHuTqttwZmV1MhC7shvoqKyU
55Ip9C5GlP1DYwXI0wRFOCqzSNUuoSRd2IMzisR0RYI+tPDpi8ygdexfszMxGmmHb9CdpxekxTPu
itm+awbeXez/3L3c0/wwSdO2nt6bME1xFUK1Bk6NSwZmZJyRgaSFaTcpwdeOCQhnmyxMFW1WjFtY
1dWG8FAm2TDv/Tek2wXx6GVuJVPRVAiM3+j7peTQegoXYUjoVxntXGYv9UtaWlF9Ki4BT59mJpWF
RQaGGDvMz25rlXIMRdjwX3QFN+6IJZJbnp/3YkY+wp/+yrNnPidT9D+/MC9bLIIDJrW+PtBDu0KC
a+0qRAqUgedc9CDkzZt6OSrxbr8iFqwjaxY+qnIK8Xl8QPfo2RgQ5w7FKraUdDAzbZpeFdfGMb8D
eaUV0+Zq65blcCAXPI06KaeTO8GMX+SyL52eEa6C87DJ8wVfkcxHqpc7KjKVeICnRrI4joaT379v
HkYxU757y1xam3fk/6XlcKRDj6B2p7E+8EmlympCx/LN1CdZeuhlJC7Tphz9JmesSjEpaZ2bjRNJ
bSyzKNGiYPT3mzuXeB3++XR16LIXM1gWQNH9MG/ku0T1SsyMmsBSBmwuw/0tOzoZKRPRZVMfrBhv
+VQej0PzP3EpEzfLYh7Drqyznckf0j2NXYqRX9ewIEVIFlxKLNijd699TPaOZFf2g+oVNHYyhUyf
Jbt3qrN79DpQKGw3IZsiN8fy8PuSy7747cnYduRvOZ+z8xC2pOSAyujR+2CEh8HOeQVD1SjjgUmh
Chv5UlkiG2na/BQRxI6Hvj+Z/zBR015UVVJprGFvEASjrUWAhLnysgrTWxPEXX8COwR7V3zEo3gt
UOMDXLQTG0PlpApvmDcNExG68ILML2r4k8fQfXcpSTZHdeIBUGEZwWOnSCmdv+5Ivj84K74mZpyt
X0k5l1fD9z5sh/wvZ5BsraaGmf4L2lxbWuJP3MO3O4Bh/TEbpF6NqxbEyAwhh3ADmISQ7aSfCJD1
dTKsOFjKq7u1jcLxUTqitiqXTSC11/6rSSAUwyuLnYT4czRr3o+R+dZEnGEr6zd1zRtMd8+mt4OI
BIWW/af/Ck8na1hLMXpS2v+xH8PJpa2BgrhReft3U2igVLW5+MPWjJjrLQOterPjfsdSvdqmiYR2
11c+kU5EwEnoJCWJDnW++9tWrxtjZotXdsTRmZZ0fhI+KfUpf2v2fqoA8YoAzTYxJFHSmohnj8O9
KjKZjMJo83ia9mt5HvMTE0z4ohvUk2JT37+0apraPqeX9RiSBr113V8H8PxIzUcYeniJHeMKfCV5
2NWiYxwemskYFlzUoB4vxURTdmrjv4394OtuzWC8skASH3HKJypOfFXNzjq1l35oTGAZEhHKFnZh
yTJQLCPj5gdaHGhwACz+EjL44og0WdXb8n96oWQgmP/4Ml6LrLIEA1zTJjb2YAY2e4oQOmk2os2G
IzHVqjWKyheOKpi42uRsRDciu0DibQbqrKm9/pLWWGAYC5mQgZAf6bX6ZIknoSWvHqhPNNoC7Kkp
1SSnJRfGdr0GVC+PdM92B3KpCbr/Z+umiheJ4S+jp8Z125CHOR3494IKcvdLhjV/8m/MTo+VAiXW
mA2qERCw0Atq+Vy2VFhD/HZ72kdmxOLY1gPmteqIPxg+UwiGXsyS8xtbNB6hzGPCPHw7XE0H7gfQ
vvM1iG2pm4faIWrCCn2ilSfxtqjP3rrvaaG3869mgu7SzcZRgwRGhlI0VIA7FnIdolq0awO2CBhU
5f58Ye8Up6k70IxyE+5pCWt0Mv0M1uooM+yhV1hfzhGmrI6ASv6ZcqFSyEaS3iPH8Pp8R8lxfXSF
rtq4xLNxtWcX5KFudcDFaxLX3PwHoyTzWtSteJmgPa1gephRJH9qoCWYeL8iXKUCLXOIH+1zG8VU
UAC2vclPAAfNSFUSmUqMYRRTGHtYl1/IxwVkGyL9mGZ0a6EAoER7kknB/bdGrznakk+S7/iVB+Sh
OljnWABXdIDQ7RGcHtX0bOnodqpIjsl6SSQmZMd6mm1Vlux9u1g2t7HzBILYn1o8g4I4oOukrIns
HSeLCyK/SAoak37DOituIldwS7G7wUm28c56wHqUyQvhVTjGx2E+q461HwR0EVEgf/i0jjvXoj6K
QpYLbOdYqH0o0+zjcX7c8EIQGBR8zE82+75nW//f4iZtQOZVe/yHed0uvrvES40nzRV1cDm/nlNc
s+zHpZgLwjOE2Bc9b/FcwOyHd1Nj8EGRQ1jR1umXradJIrBBQz9MYd35tZv07dLop8K/rR/XqoDB
TtmREOVmFh2b6Ik9WdvFF6r1BvIZp19JfQVsK7k5iHLKfaMOMKgeyPYIrPHmD9BPNVUB9BBFxEGe
q8DC3uJsozFPAuHA2jhcZiyexfetNzst7m1JjiWIFn3SaSiEUkSGYEF4AhvdaKtfMi6Z0ezKeVbA
V99aMrtbGF/FfLR2nBW2G/k4ofWDlHh2H+rxxXdmfxx9PL3G9xO3NdNk+wL10++Zmkpb1y+2yY+l
haht1j2NUb3kP+PdZFqlrFbwM+3G0yAxY/ecCKR1MgQqToWd1zFG30cpuwhGcEW2MOMUNITThXvB
plzCizRCdpCwr+VsmpT1FEMHVxSl5maAx9D/8o/KM3WPjVrxeRH9GpP/fmpQwxTIDetYuEqE8NKA
y6T7Ucreujb2H3aUJwiVY9PX1QL2c16fsXml94Wy2Ca0kpkLwUGf9qYVgsCqMfDOhBy2yspSF/5j
0dCeSNMNhp2lFZvYH4skR7qLzVwq2TFV64FIDSa8V31H3si0NfIvurXMeGNyNJF0h85d2jsRZ4R/
ohIx9BSWBC3oQyxEkS9vB7s9F+a2GMTGojUmW/vunPw77rQzLUTwxpukXPEBwDKPs0f1JRlBTqmf
x+yvmkYjeYn8J+9G4htu9JjbyV0ZsAF+DPb7eCpN1LSA7j/eTvkNpkLa5AXrGLCHxDmeAuHLNWIB
wc/2zYGRSvTRyC23Rfi89TLK50FBOggtYbe0SyKIn/yvD30n1KYA1FXEZOpUhWPf3sPG2wSEBWRp
R2R4228g+DfZsMaWdId0OqfYUG4ODax4cpF69Joep917soKjrXpijtjZdZQTe+JTqhLPUUXAMy6i
CtipqL82JtC+FBFk3AZ0DZWbLAW3r4+fGAIwSUt/SWX/S1GaiXIb+Uk+PM3sBhhdAmjjIu4LQtTb
kuc3agU5Jhdbcqx544niCtA7xBvV0WvYIJXdlyEy6mK7IDcprasjcVN9Lm5+yDUjIqLTDLLJ/U8U
bPdxwukgR7vL61QeLfscXAK4ASkoWmIGYTmMv6ZinIJY11Bz7AKfP5TbcTz+iKqkeWT12eFOEJFH
ypYmbBXw3dVzRvW4lPaB9aVZlmXx56Pl0CNTNs1gQm3PKfhWTbSgXGzT+2UF/6eUYg15XICCjOiI
867b2raKCtCc+mv7CWDI1Q8IC4yE8CJ7c/IXEGl3+9uA43KzNnJkMuSDhy3TNb7kYBMhbC4kMbgM
qnVC7TXuLxyrC7Vu1FnbDHqt7mcinbNQmyimB6+kTXl27nV057d0u7jD7YMeO2xxoWSTjrosF0Zq
SLZXljOtUa37qCgYRoCk8Ii72M1XZWvlSWE9o5vucbD9ygrKDQg7rpp3VyvNOOuDC7jBJZjJ8f4T
U8YR8obl1kXjqmRvgHOkWjqwuQJMteiRSv1ODHl9YKAtzzLZAUiE2mBa6nAoU1C/+DciKei53i22
208eiMR7N6oFQhirzStq6a/e3xUvYIcQbASiDfzzrEFKuGtJr+C53SADUuBmWpHrNqVE5t67axRB
/Jp+kTAkrzse6u6V7XnhJXAnzkM5Kt7Y6rybLTD+Pft8zObc3F6wd3rVqitd9rIfljLrT6wTSCkY
rG5oZHOwJdrN967gTXR8CIqFI5iXFyAWqYGbXo7eATPwygmXMzkLIDMeahcABrt7M4inD+NnngbE
jNOv2qSA6OQBAiDPp5SIh3vgGLwewmGEnISEQKJku49usNO5zjRz23iF4CG5snHPKUZ4LVXLdFPS
tRbWucWOPvijW9kW/dLubz7wUMF9hv3qx8lM+091nbKa2GKyn42izastP4YSL373AJj1FJb8LXDA
qwjx82OZ2A+AtGKxrzfvPUrWmREKiKe/YiSpGoko7ndFqj0JpbBrkEQTorD1Z2S3dO3UoPjm4vgK
EmpUXZq5Wv0OazQB9X3sBeoyjvZ6iha7fdmnkC2lWnDvyID9UXSMEBB7ZkKFC9FOrU2dHFcjpKGD
6bcJowpJ3Q+I7J6WLYg2FrjJuYIbnMkknBqcrquAxTZxEIWw5H6cKcnTzsWhqaThj9PpFbjn4ZJn
VkP6nDMiX6LL46BtPW55k+o24vvEeOr65pr2llS92KW2Rcz9xEjDmhUVkDDmiR71vZDCIgRavI98
G44pZo/TrX9POdHFUUvUzbL3TLRnKb/wbQJHQCZ36wPquL3JzmoYyVs2AUlIfoJdxrZ6/CLX9kGd
x7CsvMDgA1+7S553oD8xhgHHlOX2h3FtbjeD45peIQuGkn8jOdPAUqQ9M72c6V9FRpy/PQbNvPjx
rBdxk8Ncpxip7q02B7GOMGORUTGgKHsJYkpmz7HhaYk6G84iaoF6GXLifSiJ/FUbY3TotFxjrZDU
9F7kh8+w2s/4x4wY6lbuCxEzfyN0vRSWnWU5tbhG70lzAnneBXvCOpwIwbYWkBUMx9gb0gZcGufy
V3G50S9Zj6W4M4ZGiVf+G960q6BYuhFaeesVedT/Ff40qcwNKuYneOJK0g4ktONrt3jmHTnlL9kk
avhzujzcQxC42Ms7hbdhnsxKgY+XG2FQEpNo5WAUBfWz789j3MydMRUPw8W/Dn+M74IIf3gX7rqK
i4uMztIbINDWdUxKWEqEent/krubDxlfSqvCVzE0bIMSYw6/c4Yoj8isxxRaQiKXDNPyiYKqcEDp
J4J5wBXmmqB0D2cUyRh4VKD4L0b2Zw+QM8nqpRR0DZ3RiapqnNe6/tGFpyEs5E1ZqfcufmaoCyx7
rYEW8DPpAASNnsMpa2fv0NF6LdiyZAAWTcXdUpnteX6hV0dmf3Z7JJMcOzRlrPW0iaXCU/gs1ImQ
U73cyOO7gvx+uINQKT/w7DWpz8jafFhax0JiYXPBkl4aZlTk9BSMFygFk7NnbH5t5e/yvMQ6kwu8
/aA66MG/4s4uK8JdZFBplcvuuQUSyay7lF4MDncRjmWtex4SJc2FT1bIKYbftm389JrO5AE2/yxo
XUfSRVBZ3Dh6AJ21ptsezw+tldZuSnh//g31JVGJfVdd1vrDoFCdTy1TQJx9iTyhd0xUs2uO3pCv
zAn4jurwJM8Hf4tNfh+i29thPivSeGQ2lc0v5WGzqwn7uJ1itSVOTltkTYk1EC6/T/Xb81xXNGvn
isvAeoAqWyklNr7MaaoDbdAt50b03KT9PEMLryIodbK7F5SssTphWDyHZglf8La13V0ek3LqK9U9
ngDzOwgncmfg/hNtbWRisZlYBUmsF6hB0QLXJrzWRW/y2o62PSlfK+0mEr0PdS3JXkkHFw69syjv
twJsERIcJmTmt10n0Vc011U6h6axtbvMRmUzLi9hzOkV1ntEYiYVZbNDUhJ63uMMFkvSl5Ja9oEi
ET22F+tFfIwMLl1z4RRichH4sjV3uTfK18QQ9nLPqoBmkH4itFPXDl2GhlbDQI/xceQbRL5cbYWN
DVXTavSJ+7hynD0kmj9xP5qGf0ZEYbYdH+NMojXtCm0hlDDf0MR7ivmtpXQnCaU11McX1hGqIJHh
+sSdgdvBI5izce2jR3Bf960fCmQ15IQwYiAvT/iepvKak0Xil0dXyvcLb+elX2YK9bC3zreNj2ss
Z/XFm9hDjAQUdU7vrQC0V89tUt4gMxX+LBWUmovNET1zSve4zEi/gVI6wI4IkWoUlR8WTPisJRtP
WPRL8Agc2NBwuIS9fSAGDyZXUE2F2pfQPFPMA6MUiNKyb3AEd4g6Dpz6UWPf5PzIhUESAzevjc5b
TLnM++COKH6d6LvoqSHp35ocXekSaAGbVVwWkshG3/61fvUFNNIKy4vVnt8gupzY2puvJ9ofgmHB
ovc0LHXxgafPJYwch/e7p/ld07KgIoBJqwCHgXLm9vtY08F2hxpVA0mpa4oTYtoZNiPglBtFlfCi
9osMZkB8P7YiluWUJq/daryzXvtHjgPHXEMepE8T0Pi5TsO9vSAdm2005IF//YwyJPXJLstwlfQ2
QI+uXaqPV9rpUEuOiAPn4jiy+yLFWvYiIPk4nDAj1eSW18zyQCWhRyda/vbYYYX05ElgLYLcFmQq
XrRGsz9tiOAHjQkJ9McQqWzDyHdD7VK9UEKHcxU8yLegV+PIZxXAzYC/WY3UdumPOJ4fvk2pxxJB
hNmOPxlDdd2SM6DOhfdM0PosMX+YbGS11p6BMK0pXuOyxu9VmWMdzfUtl3gye/pl6AUKf1SXOpZG
zj3qpM/ItvFdoaQY3byQ3lCW4LmPk+Dye8ZdUV3EWwQKIW1eFeZ5RgN2zdDZkZUkkkkeBXC4nhhG
WMsd42HANmbb6iwGFDnC0KNSrWiBoklA+7SUyJn2/DoFBbFzAWNhNvtSD5Zfj3opdLp+O802cqRJ
U3jAOMKz4ZS6A3/+rRknTFKCxUwxnkRtwAu7ldnkEp7oUuKXq/4Iy5vKadCKMWXw7JQbwC0RbaVM
T554K218pdMRXPCsPBLTsYL98zks2+5F5qF2MwlUf+l7YI1xLBvlvZzlwfkvoeLF0l/cOnjTAZ/O
Y40Y/lSOAlAP19Zzk1nvq7uJwu2zHAwCdD3E0Msn1LIKfB+Wm3JxeQ02sV6mVD8WllcdRy+AMRjx
6zZys4xiJOA8faPYassMPBzCDAxqipb40b9/oa944W6XErk7He4vXoKPuYVZbVmkUy7d+DbDlEwD
F1DKH4z7YBLCoKrqyfb56CnRyZch945gK75iQO6o8BLSMFlxhkPaAv9Wm5l72dnj/M8hon+Qpwds
ZbONP8kuzhDmoCIqjDIU/7XeoPUVhBharzFS4ooZQ6A7UgsYz6FFwL/de3yYMY3D/GlqYcIYYJDY
ikpELBK1CR6vd72V8ynlZ2gRPzaUCU696NVtGRrR8vKSjk4uBZxhZV5hRTIPQKCnXFDFkmwflHmJ
gKiB1MCStkC+V2RvfKpqUihHUTq6O0iJ/QnNtv2QKNpWq9gOEdcQB1xXJNgODgsMfXte1HH5eS8Y
TmRLZm3yD/YkW+UHGMNBpi2RlpDCqrCEUxY6AXboBrfm6NHwD8INqoNS2dBHpA9doIIjkem+f2f9
pMTuQZzNHZM2uvvWY1Tqn0JCUMNfT/wvBlgbARtVS30V53gJw8rbWLJbp7a7b6lZJBoAoSgqsD1n
/zkpJ+kOyxGPusX+wtK8OslghoPUuq6XfZqoDYkwwoDSweuiN6qiBNEE3c1CtiGsQxH02Irw1/fk
0g4ZrakEn6U+Tb2DLYr0tewS1dTXL7sVwG4HOoIud0OC7hKfNmCI2MyaH5yZDj8J0TCmwFUxW/t+
UJJ1OAdBGJWmcfcjbwi1bauPrViwOIBdSpDXiDj4gpYy+aZR0aaUwni98MGkLXZqcTbVjoINH3Y7
iWFetm/Cq6ygS/wmalF2gTK0HsX6MwF2Y0MJjJIQcbwZHFIYs7wOYaufWPZGb6Drq9UweyBote5q
V9iw5/z8eRo2ve5Aqk717RCwGCSeLQaW0Xx0zwQ0Jp56UFiO1C/4kQQEK9sGfXWXlVgu6m0gbe4L
vr5/2o94OeDjKXWADDMnKtHb/KWvji8ct9UHiYLKTP98qcBQPyoSY94zMkj404TOpVxKBSUdUBUx
bNhKkvPanZ1bGJv3fimpmW8wSbgc9nHg+LrhcsYH3l7FX4YRFRUzxhC/24VmIjZTV8mA4LzT4o8A
CqhHDN30RXST9+YUkvacTyCuTz22gbvsDgFXOLAiuV/DTNznWUMHfaE2MN4QJg5ZwOjoMfpNUYQq
QeetMeeJMImX0TFjH90B/eEyAKPbhaoDQy/0azSF8z5eRlXdiW71Z/9jypNWH/x8nVes9ij+5qzj
nkrjGYBxo+aK8cTlBeaUg0f5wHFFFCPFPD5DyzKrnj2R6mrAoQlI6wOPiomWe33L0P2Si95l/Mlw
2HFYezlUN0PocT93lD5nfxdYkAL8cgYSDzOvK828nAFDLBOnBX0axKQakFh12J3KhftU3ijZHiim
Jlrws5RlqdL3bbAjl0m2MD9xGymufLA7uoJH3R2oiH70uwmWonvesqfApxJ6NDbEgLrqbZLco7aH
IwNU3d3T3GSrr6b9dbCqXJnDooFgiwj+jLBdOKvVHojsiST5WU36QE21lDbo48HtvJGBKlbIW19T
VwEdT/3xqHx3+x/HAqWCM2mmBkdrPlQhjK/ub1n1JYGurBqemnHsmz5HyPklJhr5G0fUhOmZ5T5G
wZCeu+vbVcZxOQMcR0Nhtr3PwChCSalFU9vEtlr6RV00iY8cE59rUWoC0tZFwJftAyKtgchUds4g
Bkis4W5nFdD5c8ElvgzDe/jHIlBXkoj3sha/usfqhq5nuamzp6blQUlV/q8kqCU3GVU7Wlo+uhFP
FJtT4EUdGYp5xOZTRAFJHrRdBxJL8Q1XRV4iB1LIIbjGY/qwGiXEHfLcOswlvR7ihtrg94wjaSeQ
HVqqoNl68LuPqXKNlgpasX7RDabXZr533GGdqQAi7ZOO7+jy/8BNNpfkH5Gea07pt/G0qfy5KYSV
G01KsqzqBtwnOaofWZlEcqJ0BIAKXvu5WNP2S4tCLcoLn5VSxlTMExl3nNEhZmfF+pnjkWdMJcQB
fvwUe70XOUP67OJb/WIw6i2JB0KNdjNhBf3Ia1PXri94ZJLg64jpMNix+WvEYLp01Qqu4ZkG32fP
moxo68kDV0avsGgFAG/hmoxoOJZwXIhxADhKb25LmvfLkXBDMGb0BgcUidmG7OkArb+lKKs4Qleo
580TxAkGixwV8VP+yYqlIad0NgpuPyWAV3lCATXauWjpIqnTgqNg1fcZhRfG5zMZuYjLT1S17T+0
49WuoqGDE6DngWjCM5tKJN58RVGNfn7XvXn5cCiMb8HIgHz1KayTL4+CsqyEDIxy0dRhjHmJ58V5
rTvH/UVmdMp3EdRogCgIugVPn7PaupseFOavSrT5D+w0+abeCAbXTsJd0DCOLOci0webxWNaVaHz
GYx3hGmtltEizBDD/FCZRVmYSdQHdcMp3FuPxxD+O1kGbbJzzhT+mLNwn9l5N0pQxoqjd9Z3xmW5
O2eY8/CN33AWHkx+uSDvUojEF0TpDV5ceQhrXbjGuJzzyRU/OGysxsXl8gNkeTODLk9mdrDx7zL3
j/6MieSdf55CmwOFZDiw1I7gD3ObqU0BDwecTybFc0DY9g6JPHeFblJAE9shbIkfj2UZNE3sXvPi
+MK1jMtxTNYH0zIauDuebSMo9MgcnDGYrf7QJVk7R6n8rdtiIXXIdOTHn9x1NRgN8z6XElfJQRwn
zOe/ZbvX1aQP481w0+1GjJ8sSVIX472N8a0PRlR1r8aVSpH/N95v3dn1Y47/3f/xJGidfuoA5NsD
i9XL4HmaDlk7N7DtkgTatjnG7Y0HISCRjIc3+FldSi+XYi0ff+b1jmFsoB6Rrf6bKWUYwElvWjxc
nZqHYI9qhC2qBWxbj/uVNt50v8vZAIbfP33vH1AE6mAQhqjmcGkt8z2vC9rZN98/dnX/7ecPfoDT
FQWGl6I1rOFqLpL6uIlxNSYP1OFjP090apO5w75O8T/niFLcdMoL+/BwyZf+jvpvvWYa5ureqxvZ
Wyb+MUk6gXITGgTASQR8TrkL2tfj8zhAzz8Oj4Ur5GjJyoL1fNvS/ooqJw1xF7uHmL9zZ4JfnO0h
8olTsZ3xkX2CRf+TrvVyNb/jKlJidAf0vu631fjrcPXe+bYsJ9jF6+vYlD3NtE0V+JrYeNHFXd8k
HLDyMD+Udb1a/uzZL16IrkQKeNIMFLxhD7yv6NhbIjBU4J8QCkQv9CY64K2lHPrB97q37W8fkqkx
b04paHmS6/P8fcY82dQRkGW0RLy3zuq3Sj2kvVX/eSbR2j6COJnVx6CVz+taWfpiOYhn7gL+6k62
zR1oYVt7GpINDMgh+yiwAoVecbARh0M0bPKSI6MRCxTlqfK1R+hn8FijoYSOswkFQCWt3UC7l5ej
AT2CXvQI+gvVHvZa6GNziTgPN+xZWanIlGPs387RwYkIUMzZRUiwzJ8XG8eZ0TnHO1HUpRsn3XX7
ZsYvZpn6yWiq2DfcbNYFl+sgUuNWz6hakPiDUI6usKYDBmT/80+IHkFh9gHFSyPhRO2SRBrjwDHg
xZN5hgm0sDXmyOzBHQuccYVILN2R4dxdn79UQRiUDpPTbRyltuEp7z99dSqarUd4Kvyn6sfPAS24
KW6K8a7rtRfOlrGNitIw6LN7OAisI8O3SsdOyUizf7DyeWx2H/cARCXowiItLKTfg/BohEkJvobQ
hu4grfumKc9LyZTbgJ4Dbto+CB9kVzzmetiBULT93cadyFbs7RbUyYmLljd2boy+bu/LZeJvYpZD
AgxhAyE57swhxysXU4NtqBuP7fdIdo2mVnwR1E7YYJB8ifgwk4gHoliXCuHbJGkR7uCr5voDS2CN
kVH4/Z7v8+B6Uc5KU8GljW6jOl69lmDUOCKKk4Tyq3g0ywAl/+dPdEkXeDFzrTA4K+lH6R5UkA9G
km7ExtVfczMpnb+Z4ww8+0EqIkojrMnzpxBak34KDtFMY0R4JwSPwGlrHxuXaGAXkz3/rS7+SInd
iUIp/arkXMXXeTs7KPPoduD/UviFHCb6P6T3nKaASgBf3VKYzuO5ViLeLmhXsQuSHg7fBk4IKVFp
g53D7JNqe49TImedXfbmuR7TK8eR7+Uo+7NwvDCSN5mWP5TWHHvUobfPtCwFCUkkzQyvQcOSW4SD
nxFsoQQBn01OQbzXVtkL1SGE1wj6mvUdwdl/GRTAcPHTAnkGX9lstkRRTrfA4p/piINcD3+GB08U
xIbbf4J+MIj43juPRnzYuq1ch6KnwPwrTeldVtmTSBz+4Y+eiZR/9TkcNQaVD2aUDkJWnDAblhra
00cnpb7XeALyXMBnLlPrgh2N72Ycvf1GgLGRdfba5S01xAmOq0e3mW/2GIOyk4oATTwUKANpvVV+
H7FxZSPMKSm7e0vT2BUrRLh/E3WUJQpAV+kKEQMVVWgGAsV35q6EmT/aFD0+9bo23eGg3tOQNfPB
2Cz7V6fWp6g/tKmIK37Jtw6nEnEfedQpVZhSwkDrjJ3LYc581w90mgNzsHdbjg2YG+PFRVLwuJ0O
for4OFvDvzJS/UGQe6t74z1GGaSvM3A8btQky/bS6/3RSYWutR78SfIyl5WMZIVSfNlNnMQ1HXvn
5QY+NiieSHGg0DZEqmx4aFkEazg9LnASKQGshKAbWcJrThx743sI27JQ5cQu7pe0wVDH4GFlxLcZ
OyEjdiIGqQippsfW2Tmi8RdHOIBOdrKLoDA01w6d1OS8pJnEcgDXvDoBf81oilGg4Wk1NJUspwLi
dxY36Cg4V1bXUymDDrbR9165CqR87NOXUzISDW7CjI9Fowsvkno01bop7cwjQAZk3OLSdohnZ+Nq
Cak9USx/nhKcTY5DYUYI/fYw9yb/aYaupV/sc+9HfgFZ5cVhDnlTs3Y9NXLHSkIUwa/Dio7fEL0C
HCm6USrdDYElWZEzzUahPB/jF+Ynw4ehDjLEsstmuoi/eXdxFdLWNf2jsZzoLIeimZGVh+bnmBh/
X+dtf+a4KGauEFbkrzACSjznmS3JAFQkVVR+fynzdQY01/0V5NDDOoB6z6qYlEQbMwjQ/4nAgDCE
W6QSXcfAaRjk2h1tOgaPA5Wpoqcp1fm5WzDgkRaWvWQ8eoQlui80qahwX849w0NLCgRdvprWRK3x
0g621RYlc76sORyAQygbhh3t/ZB+girrmXaDG2XPTqDXxqyEbMQHiBXjMHzLhPqy14NAYUYhqtDA
UJlQmiYqfig/Mb1j3Cg+eOMduG7/IAk8ISLjg2blQgw0JnrXiOBHEA9woxaKlU7sYrB+2V2ShfYJ
CIqoGPwuf97EF0rONAq9vFAR71Tufo7+GWYZKJAqoeV6QZCeKMwzDIN5mbDZKqdA0wi+mlaLZEfb
62Mzjj0phpKQTyrddY6xYoxKus/YeernJU0/yX4nxbxfEyJR93R5hI+u4w3SD8Zyw5fSqsRkE0iA
haB0kfX8kITYqsOM+gspo7slP7v7r+WJ65bFFYEnPBD66IXiJoRxdd0nwQiElhHkauxNxC3Lgatl
lThRKST/IGLe2JZ+rhPnyVmte2FqQ10xF4ZhsOWeKfwdQY50YQ+oQFXmH2Vr0dVgOQpHaLwHvm1G
FOyc4uv4lzevQRZgAXTzbayqwfNrbNclc4pfb2Wu83fTZyA8Gx7KpTMVKHlGKQBnNtGbZyfxrtSt
wIn5OqUELMgrV5s83IwhuWkRqZxMgJKZ1LADhSEcJtlSFM54rDjfsA1mwXzASKHO5MPMhrh/2pgI
Ey+Kd6PAvqXUDn4xhIotC2Va6V8slX+jz3vuADUA9Fh4ImWv2gQDy+S4gKgwURx981umPN3UJZeW
wh5e4bqNHzSlj22cfvDru0W/bLU2wfbATavI29l4LeDTlS1ANsA1gvS+Fin7OZQZV3XffUGiTyCu
+qYpJmygA27IkdKgqkPMJ6oQR12SChRyvthkzdwTb4MNV82z6PQXO4SZnMYKnnlDyN7TJXtrBoHw
zuOH9+ddwcfnmSkPClSR+DJRtrin0r+jibNxuy8Jfe+90vNeJPQWH3x8Xts/Vx8PzW1x1TxsqoXJ
yfCWb9TdcFNuUEW8DqmGDR32R8i68aGMHuyQankm26mKtSFYHr0BJMNnuQn4hrZnv6hFk0kNJyTJ
Qr/jfZSdjFPaUAJkwXhtI8fh+yAJP2I5s83N5nLygUCU9PMzaUpBWJQLXU7zXqKbik5WVe+Js9PL
f5NThzHaIQMt+cfARNwkUdJ6X4khPfdHHEoKuHztwnHM0FHfgy/6QpYHCuINTRbgwspj59n7fmeD
sEtiDkLB1aPvw4KJB66QfS5FO21PGqcs+C/+pw7gtCsFKhjKtABVb++GWrVnPfMnhx4u+adnsJ0i
Y21Kp+p9yslSFuX4E4+26hrHAUuSM01vKn9fstGywUPxnRW+viHcRCp8jOYSIsx+lZHe2+q9Tv0a
DVdqxlMl2MQQMnbUCxFSgp+L782M2ZhMeEn6mlE4CXoXb7JknftungQ2oGavubTst9u64qHjbUoO
6VMOVno4yMJoHQup/78ZiAXTJDX5jk7wYbLMfOZQcJC26NF1nWss8Z8rkRatWOEy0ExRN2sX4WCR
uMhy5jiPS5nFFp2ICO/qTkypZdjzO8iyE+5EOfszMNAJ9R9AQ65EULk+FfL7Abw7IufIXBm/bBgw
bwKXcwlodbRoTQtn2Igdg1dH3sppbACIPjBOroljnkfskQCTSq4RLqRpGmac9mZC2zdFS8MaaAji
l+CSyjUOWbvQVTWIXeHgWgY+HCSZNypcEswMdoiQipxcYfr7YNKHO7KDybKkdUQSNsxrHTlC5AQN
WLeABVuDWnYA8wTzh1FNtJEFuFzfsAlWH1Xjt2mVpp/F/wT2ydGvPh6jiGfNAZE7Iqe69X011n7i
kCsUg7HHYCF/tRS7PAtn0MTrplcWtAeQo9cauowxusz0ICoveQOB+zN0A7kVtjYT5FggfFZgU1ZO
Y/2VpVraJM/7l6OJ7b/ywfWdOvDz9SrC33DHCNLys2Q++9qlUT2owb+V+K4N1IQ2iHDS+D+lcnBF
yQWay4yh7peRSf5dNhyQcWG6aZt8IA7aLK+xhKcphqVDRzMzvItAYUQHMHIdrzSA6NrVvhq54Q2h
TQdDKJevsFmaV120UuqsWvW0HiTXa871zEVljaVLT2PVlRydqKIq5dSeEQuiqd4+cZdv2bIrS4W2
e9PNp4IIjpDiB0BjHmFlxKoGEW6PRpN5MTtMnwMO06901+erCuycMqbM88D75qpHkzIdKIF+gXth
ijtcndhH7fuBxDEUfl7y9a/HZdmvZIvRXqGwXY3I4LuJ1Io3VcvWP8b8XPm58eutJvbWl766N5qg
jA2MYAtlyc3eN1SWUerf+NwaZx+DM3azjjXUsF16uOpCdFjkGV5OYb4+DgKPHFUWARU3RazhzVbb
kSqtcw84Ck3mej5eZYn2q8TEvDOVqTPh/6hrBO0YHByZFTBW5tgsTDkwFMRmdE4U/3XkNoQkV4pt
ZqV2kKLJTvnmIup6sAIm8OgkVZxPkoXBhUA5gQyxDTJjiqUGObMnPd+uCQosbRxYRrXuuyyz1JtH
H4xQtcdthXwX55/R9G+5AiHFF8Z3vPZhR2rD71Oh6KGIxXD+20a6pB7FiI/pRIUovRgdV3bsGlNi
0fQZeIdrP5o9dofh76aoZq1mosx3vOMEDzY7Q4CEJg/tlQZNRT3k0w9ca/JsZLBV+y46wfW7RHKF
pJvi8hiU0292Uy3LOpaU8PD2+LOOehcczJ0eCCpo5tVlxLISNV4Vc5EtttnnytCOKHZY//UJ9BSP
cv2EOHy4zQttmVdWCeHJNcDNTihFaIh1lR/W4t0UGcIv1j2UGiGccIZ8Cse4CT8/IG2HxUgIVRwe
BU7aM0vWBlHCBd2LG4YWcCKUrl0Po2SjFJ78gtk+MLims8nRvTopFvDetBLhK7tBTqgj0P7p9QwY
LJwPw662yYYlawwU20XAI409c+XLxGdHHuY5HMAspEHVHbQ1EKWEtUsUSVsLl1+hEuQvlnvGGs/n
+WdpoyF3WgqGWMM7RMksjpw8GQgnqVZaEYMOCneBTWONMuG/lxQHDG8t7W/53POe74Doqy1iPQkw
xDpxceXRSwIVL3tJUBKvV2urkspRB8NqPY7Ld3p6FFV8NUYWIfbyfbBKMnXHJYzwfLRWLzPSJnR+
tStgEKn8UK4GxjgmMnkG8+BJbtKfCvogk2oURv1K+pzNRW4NH2S/p/UMtgxC8088nZegJHq+g1Cs
s8h7yZv96EJK6hVl989ZCNeVdumCoWISpvVrIZIfQ3cWgRsEASQ4jt9W4DrDP574nwOkNoZXueTn
SbpW0ztVxPlRY2HKKhrvH2i+8wGiEliCmQe/6aiPzzqWWQ3TCrasU2fmVaoUYP9BQoo3ux18y1UD
eYqgSZCs3PAzi5KH654BsrcMn3gU4YfVcDhnN18Y3XImd3wOgLbklDxsQOzS+FXCTlS1Or9QcKN/
LLBwv6Phd3Jj7ibal55Of4/E/L62yFh2lCWu056uiUDfntqUBsWqEsGid7f59ldOMSZX2sHg8oGm
54MlTXsGiKDl6yR5fAhzNT6MtlpLcw6rQrm6GJooHX4og5sUxZOjQhLmPfsD29greDU8ENne+NBd
v4uPbcyDgBeWNnxLhofpQG8957FjzcPlkzMcmhKL5Eky4UOAQSb1owh5M6HI59LppnAlg4SscfeD
v3PBYgj7gr8nS+3JZ/wdpBEXdZoeP61tsK+b/N5vtDL0oOxCul2T8jXNbohtP83XCZFrvHuRVAeM
/UtsxXxh9u4mM3RPgpGbG5SkrdTuIJSMJRPyWRA2IHxFgt+JCpalbdwCAcLbBMZcf52y1XlnnMsm
15QjDgPD8bLCXc9gSztDwofhGNrTCdZuCpxE9Aj12wSjj25SrhNIdXohvPO3dZj7DDdSQ3L2QPqi
xXYle4KlqpoM1rkSAL/XWqGocuZVQGE7q7qAKqZeY4AFNRN2AmIbPhmJqxI3F9YprzIuuxgRTsc0
+6+4uoISLp8/hT8orPMWYkoy+5y996gnLL7qR9+3n3cDqnAJ9OnGYiyzij8OJEAyjAoAymv4aApl
h/QJ62fom1zryKIB5IJLDX+7LTXJGiYn/Srn9/HquIqbipb9qe+bu++Wo6cI58WPZjqOrEMovwzx
enDNTSDdB/xXdztWKo80bDoTy5fzgkHPBTu/5II3aqTAYAEzrC2yv35k+sR1hsCwyjaYTZ4s3AdA
AOfNubg90nTUM/RqmmcwsTvn6zcXwd37jbJg9U9aWxUcAeYCFkSFnOPdu+AZMJhuKDJFKYPh+Lgg
bJJnBxUw9OHkBdh0W3Dt5sL/YKthhHccDKEiw9bPE2LRCR1vVxarhkuG+LMAKVxIPMtL9MwOQ4rF
1bUElWKW3GMg6fnLE1hNh9EUUp6WRtw3AXahJcoFJxPXxiW8/MPIUzbmH5SSmIH5pu95++lAlQIn
EbWbS2fz52XIXh2l6Z8vqzDFzo4Keo01ddQovMqmT+y8NsaxVL9gnUTbKqIkxbaZntckNK0Kl7Um
UUvX8m7zGoyV5RKWeVXIr0gUKYTQLtIpZH3fsc8Oh5Q2byuXdjzZDTsm1TnFLVjz9WNEEygj+0LI
phibm8lfHdAEuwBHVM4VVRHR4TfyOdS1E7JlRzlb2c8eWqGOz/5s34jfX+6Gg5/sUAdn133eeOZ9
L4W1putct0Nc6IVTs6LNQA0V9ynD+4Hj6fv/3OLoxrjsNiFEPkd+d9Q9njj9N98DyyHzyr5BW0Db
RvVLjN2ehnK+5/NDqwwloyEo3yD+NiZAo3Ery8ZARbv+2XitcLcWDYCHiJOauWwNNoPY7boGC/GY
wGxRxzkzZfC4QRBZMc+lli+tCkhsDGJ06m7sV0ko522oQDzZ47jyraJUvj7TLZAyOaK0WesplTLL
NwBZysc822LD+rnc1gj8LH8uttotecvsabaZ+pjIB91wGXGwS1A3Ss9ZetCorJybTnXxvtaDwE5F
72tR554XM3T30Tobu739ZfpSjHqlIdvILPu/RrKHv+JhPD9oWUD6MGsWJjpKIOZBmtrnEnBKDgY5
LP5jQxIs56b8q6mORwosrRxReziU0X0R0Y5DT99GYkRMYcvNkUJCcCQjHYJgVDuzoacevK1fIcz/
LYHOdZim98epcqg4xnLnfb9twP9Bz7wh4q+/qp1U6PItDZWP9g2mL4R39qRcODuGo7afzKi1Yevs
86Z1xfyptDkQojueP+wi4HpV8MXAkJ0/vZSJEvO6dreNIW2tLNxvZ2uwtRsU2SpOjUd1Jaj1QKwC
QSLodOhuuLVWUTjmkuBTXR4SsCKkHtKvVMWmYFzEy9t7b553wE9IsSXJ0H0I9ReEc0FrrxBoz8Zm
K72GtOKktv6OZQUvrmngD+ysMCRCh07FU8a34jDnzfvaXpCDTtKvzASxCS0uIVZB97JRDuQChOzg
HG0EouFhc1j2UrYzNONj7T/MfoEGh6sseCOLwpKwC2rD5UVG891Mws/4f1QX6TnqRhxQ/1liA+cZ
KTIaxywqhjvtrzXgXNt5S78myx+5dzv0+LTC2mRYnFij5wElB1cwVf01ODlRoFgdpPV9wy93jYQ3
x3LqKIc1ZQzJFCLQnIQLE/Sv7Xj/xlEKj58tJZ34a3LQJRbgkPg0d562ZLAoY6Us7Ga3ZsCq72ij
9OIvFJpF3/yYZ2IBNxMTKPEl1wDs4KNOMoxRCwFGrkKHlS8ZGWA5LWxSQMsu3TgxvUjO8kmrdQi5
7wzGq/juNfVx1P8Ld/oXNutWaRrA2dNxZgDBJ9KaspIMIJNrajAYA5lHy1DxTJIP8HqRo7NJn5Lx
oy+E3C+FpLwjNSyJV6bB3o+zAf2cdddOGnEf+QUYWlbgsoe9QDp+kp4XE8ZPJTXm7JvAcr+5BkeV
86zz6Nsm1RKVbz09pl1qdmSWNwpEq9ZrGZz2o7n3HqsHVWWHruZBEHNyUG6RYkCkGwDgqThSW7T+
exzhznKl9jxBbX+DDD6IRGYYeXS9MwcIUeQRL3NU1pg5T/kolM4vDHaWN42ryIO7saH2kZ+j8pNx
I1luI/kPulJ9TaCFWi12mRR9JKZA6UqVpa4gGBk1jlRR8whtErxjxrb6X8Z0u3+ePhjgQanNuO9u
3I0wnI81o9uRq9K9CPv4O+8XYr21qHsGfBbBOTdcWALds/Jh+k2wSLjrrEahH9hN5Ep3vDJKHjaM
b9sMA9ZOu/5LLHQDilzdDPK4fWow+tOctmTp8ZMZ+h48oWbtVk5hTsrEtxFeuYdb2YLHRp4eEHp1
RGrmuDX2O8+OOLVXwY6dFVNbc4x4Oc7cfOn0iIkOG1yIq1OtmQQ6AkAL+N1n7RlZ4iRuLOTGkl7d
PkO1AKkKckC82tiX8GT0JSnJn8wHGDgxAN8SjL7OvRabSKR1pzMMGmvpQ81CSzDTeTi+eHIVEjn6
3CmoYB+V250KfOpaMkwztXHSYvPrmY8k98FMU1iC7RAl3up+X/gd8UlC9Sw4GnYimIrsHfQaXHyK
rpU1FXt8mwvOgS6f6hPGNuC5XzNANuLbfqAUq8Ze/Qci5uxczoi0PLuuSbCJDBJcH3YTD9FwhZ/j
taWaNRmdlPR0Fl42hsZHeBgfp3Y/CWDyToPdDdsPpR+mPnWWbh5rq+aXrtrr5gv6A7J/5kM9qI9F
44FwzudDw+V7yyCR/JhVoPbHDMBqY74Jxr0G8gSgnrsEbcZFlyalEDLq/EqTuA20ajuQVu2VfXBf
RFgxBDmBclrSx4rDkeXfQh41tW1hJk9bedDuUbYQqxHQKh9/wKsJUCc6N2IU/+qglYdxAXCN+sdD
GJyb4deiaTUDxmRd6gClCcv2O7kTPsXhAC6t+8bjrZwCIv80MPHbRx3qoFWak4+PXHMxGMfP7BUp
2ufT2aMSmYPaen2NBXfMMErTI9uBekxiXbntNXRlG2m46EDAEPmozqLtSHpQQrRHbctv4G292IYB
kiMadvB1y8ArL57kxMrwTiwQvNL8RwcHNaFQCIddnKQd6jaXnR1xIOsOFyJa2e2e1XkhQzlynvSb
h2qHzm3MXxHaoURTfW2E2oNLbg3bIzEEz2opQxJ4ytl/dGDoZAnv4AHq0zPGlVx2klmeM7926owE
NGRk7lyO7Esuk4J6/UZn02+WqGMS8n499vWEXS+7fsmZFoLO/nIRX/3RIulIUvZl699LRq8nN6em
8AubHNUlIdk7Xyd/sWjJIx0da3oSgFYdoSlPRcdhg6LxlBZhPCY4fINQ2kVfSYE35osUfxUgJULf
SuzVJf4OuUX4BUtCYdciM+rPITI9fcKrwQTrDLFEWkMB7Kfnzog31uXQT+x0xYcZ3T2abl9uk9UD
+kh1BF/hydNicGlozs/4iW0l5XYlIWUrgiWiAIBcqc0r/Uo9ukuluydSrNzWzi64KaOFi3asipGm
+U3I87yXBzxMv4CazZM/4YJfN1aF0w24r4trGAN4Yufk0ScBi0K271aAmub5dni1RKaX7tyf3nyJ
geg6awkQws73tBo3HkYq4BNSYubptqwpPTA4/q4mlPaI123FNyX/O8nNvXMP1DMUG2RP1tJ4LKGj
5RlhWTlEfAzAgqJOMzdsUPRDLWvngSXlUzvz0t37K0ofvxmNeWMAvyj8IHIX7JlN5dfke14ggt3d
Hx0W02DJOVtU0FEmOKsPmcblp6Nxi4TCwVaA/M+vcoRzyz8+aEExD+xLwOQh3bujjMFNapJtwQ+q
r8Z3gleWBKf4VOZVM2SzkMQctK4N3ksPqaq/kQ+HPldDW6GOQxzCjMMUlWNHemaOFkWeCmoyrC4u
UOUG0DBJOXvFP7Q71yFxWMiY8Ue9xSi6DIYwM/QKiyPHyqBHyBAPCv9z6G2nt4UvuE2jGZbubT0l
snpvLfLqEfW+unIjNU6hdTWU5qMsgMPwdexAooHhy5fROmWTSdEwY5K+8xASJ0SyvTSxrRhuW3lG
C+c7FZgJZ76eQQecBcx4Z0bKEb/nyxhsxhwQ1U4pwQyF/eUXCQRRI37NYRqmp+zQfSZwRqyw/WyO
QSy9MTwFLy52FhkACofAQlTDfIxebk2rfsANrPl+B7uCsN/1fHDXKPNsIuo0rW9dHX3QkiuhAAe9
FETs7ZMB3eQLGnaW6pVm/fsxxXJi6M9lsiQxG/y3r3GGkVMFgiBDFzix8gLy793K60UnvwOdPCUl
sDrlwmSTYCEBA7WSfESZQcgZpJtp0P/goGDiupRQ2yvQJAf2vfkJJahmWaOx3hgWxMIai9ZBnxVg
xvDZSJdvhO/40F3Zr/2T71UXfUB4bEn0LizIQ168yuMb5TIpmsSnPVbhIb7ZmMTbFmy8xwyImG2y
3hjGFCsPLuRQ8obSVdvXMR18Tmbu7WflTHWLT/e8n4U43LHa+DKhfB3XRDCOSfECp1cFUVn7qz1n
TBVTu+JqiruLBBsMJXnTahYi4OS+IZkjQTL1Ih651ZC+jjwcDiU4avaqHeO81QXmL+5LaQk7br6j
bj9wiGzW/JRD+D5ybbBRO817Uywqfvuru5d9lg1Rq76p5Jc84St/w4dXqHmfCoW+wyuURoIddKnZ
3Bdp3bshHv2NOxXHDfSvJXRuV79UKY/6kmAQH5DmqeRV1rHDbo35M3AEPRULDoliC0BI2ziomEix
Si8KIgDI4uptUE67sRjuZf2uch+ra44lGk3gqHG0vPznkapkoT9pU4HczFa3llDJ0oNWUXTq3ljZ
/zwMrS9gTRwyThQW4a7juUXAUUeLYQtjIqYAGZxdIfBO/kreXGek4JG3Gcfp5+O7IurCgLvdHVFv
I1vfpAKx+XP8p7U5KzBbDk4MErOYZW8pHL0yzv93RAQ5Wmldll0WVcKZoaRlcv/NEkLv2jujMuSj
Doouo81WsHzcz/Y/tgQSRDGIkLq+YuGeBZKSHv6XhRmpXxfNExFFjZQ5SQIAIS18m4Q+vMOJiaWs
UPz7YVVowUGBgHAm1d3UySdyDUOI5LmMAbabSh/4zSObVz+IE2DJT//nJct1xEdiRdgp4ScjfZNs
sALP+NaRWbjJmqFqiBAPoNLPh9gtW8aPUZgbMhGHG6oc9N1qr5ZuNacsnl1D2yA44ufpzxJT/6Qb
4TT2KG4r2zKt7CFdOsl3VqeDRK0sK98eM7/NwBbriB3sTsYiEetrEErSr2RXGj1V43ZEu4Tnbd31
b+gp2M83qsLFPH4iPQNU+ZZ9CsnnYHL5yDFiv+wjXeQbsZQE0w0N3JDd4VCpYNZiuaFPgZGAaogm
tyDlv69QaW38y5dJznifji1wNtbOVMwT49hPbP1Zld8UU72oZV0MQqrIfnd8sx26YACnkD3AKtmg
v5qXx0LwJuBsXDEutGB4r+vD8Eq1Z6UwOWFmz19Eddl7QL3Ho2xqj+7VRs8OA8u3V7G+WktYMWiy
6FXN7n5zMRch66Ifpnq4SRi+j8ZsnyTJgcu2FbYcKn3MOyucZK5Lwh7z2APxl5j5fmu49K6QUXRU
SpMDEUmd/5E3lfxn56K7dHbUeBqV+IsGokXm2b59DislOFKDB3cjU9PD0rZNbXYHgCn/iS+Nq2Tr
J5ndz/92u/knakjkZDCPK+dMcqcip3BQY+MAn60pXZUq+uMbg5866JL+nNyeYtn/aUjdBQRkufFd
a8I26PSppT5M1Im/7g+XdPgrmJ6A3MdQV0MSQxgzHH6FAkaTpdeDAMHbUidIr6N7xO2I0nHMB+hr
b/ne1W7UhXzjhUJuSi1EyA2ndiMnylry4nWNA3R68Pli/9x3rjsmVFw+8kZPYz+paIC2gtVWoQ2b
Wn6hD6Brf8OG2dmi9Lg3LsD78DBBtyA1b2q4uZ6XuRYeNUaVDLNfdAUMJfloA/ifjn9NZEDKEFiF
8EWm0GIhBb0RRxihioijefGMGtFmYCv3xlh+DrvHTbaSE6SpvIP2ib5D5uRIWICg49zaJRPIAA7s
qFFarRzaK4VmXq69UprUg9SHd1+tPOIvNeYbhkplo29zWJ2esgozDssREzOXeCb18IMcN/Z0HBPf
wQdH6DRf1Sj5NS6T9/Ubz2O23FpODOXHSHcncmhNURLdvhyhOv7U5WBmD/SjEev+GHdwIc+u9b0J
SISVssXwu3adzajqU3VtE3/M7VlHq5taIzLzEfKT6fdydTIawWdu91/LJb9NIOnXxy8BtsM3fFh6
VjBApQrO8T6WAQwJs0nd6xk8vwsAUPlJ0wB5i4yR/TRhyeSE/Ph7nu3F0sRgCB+rZmKWAsSnUx5u
xDtOdIez8ZhoYkdkQDd43DOvbqxpOrjOJMVUVMDrXwZesvF8PniAPaCgHhAK6MxtEVgl5H446hqk
9K5H5BHLOsexbR0sL3m/I11kME0TmU+vz8+TDWMFvUSEzd09mJuA2IIm7c0LDAN65Xy4Fp7xYcrE
3ofJiPA+9ikFUn14IO7vMOqAv1VdHb3KWiVz7H+rdWDWJgDfrOVM8qsuJlAZeXXzqPNYAwMilVnv
+eNOkvHwDIRCuFJHfSmXadequA83nhUe2Zo/rHBl88j1ilEzMy0G+VSpE3tqXu9hKTwPgkYo8HRM
zLTam2L5QVEPN1lut9OtuxnsrSLy8t2ujPpIJ+uJqsdC2H6/Y0RrT5hMRdFkE4VIWoLW4tVU80Fe
6efMPkOjQBfizhgX0WTyW0Bj9Wf7zZk/mad5Ers1ug0uC+pYG7DIVkHoAnISSC7Vxhok8B3R9gL7
s0Vv6EJcJRuBOyjbKEka1fXxnTn0A1fz4tbr70ydYjDF8iiQUHul0buxXxPwDXo3CLfk3Alq0nnJ
yItFM82N5tmci2msYsi6mkXCQIWkTVDiun2Ohj+PWUOAyvERtBwTZ9srOBcQ/NLhWZKHFXJJ3KKv
lcgWDb6aM9rMgCwe5jewQgAxrFZXlrfMMyurvasfEqYfTnw7hqvjClVJuy6q8ufVYfE35HI3mVnH
moZFfg+0iCrEqSsyjwtj2F60YHaIcvtFgdStPz6P5/eMGOZ7J4f9NXaScGyEAhQ6yRFp1AFbqs/7
2bXYMmfE2vAvoDTyy/AsGcI19Lu9o092oRfbwpE3LPKM4lIescWa3pzXhn2Jfhc7r3gZpyvE1knX
TNCQUDWsjQPK4H7qQeCdQCFCmf4MkOGdvmiVydIXXxi7C66e7+fFLfnWQ5a7cb4u8ApPFxeEJ1yR
xQ8UCoeQ9r8puV084/49Po/EbefM6VURxUZA7QWXUWQ6ou3MyLmtx3DBKm00Vw9V0UpjbodrNnNK
YmfaBZW60pFjhKc1E6UMeQprHFVaC1B/o2bLJbdv47yLkzrjCoU70dWutsc25b94JVxoBcLsKpwz
qTwS+dshD7XYYKqC1jl0Q/b6YA+J5uwiqGUPlSUkfDaP8lhOAf3r4pyHaYWY24BvJMdETZnyLD4R
vdtAHKGox9/s6pPyNKQmJMH2+TxYRhyns4PmhciCyA9M3VlCbA3aeUfwPwtP46jACGYjL0mjbEBM
wkF8XDkq4oU3rTdexdxiWcjJz8NfCbAYfWL0uYOtKaMemN41ASEOh/WDBB1X6HFu0WJ7obl/4jDa
GH2hpJ+nqYszjIUXYhc93I6U7qtF/KXqJ30nezOpOeNITinZhQiZj0G/5PbX/V028AvteeK8vdgA
pVsvpDSLFxWu6gKZ5FH6zZXqDZkfvMMoD8b+TkGXjnGS+mbN4II9lY9bK30Wz+ZtBU39B6cfoqOG
HXxlM/ymzmPqQk9O0dwgucN7J9MUEsHqyzsXf4F1pG0ppKdxaVQ79WJysV+QeDq5lZWj+qXWzJcI
ExepRzPNek2PCQ0D+3pmDpjtZE+WXpiqK3wo9iNbiG4MxElHQpK6YVipJykZ3x5AJLogg+0pYW4E
SQT60VdH+B53UdD3takW1U48/XN/xx5xenTVTQKLGZyRz8eWSm2IohonDD+ks2f2OagSeKv8l41B
mZegr8gtEn/IIDpoQ35pkrXjVnSypALREmYj5zg1axargQCOgANhBnEqMjj4/+0VP4gl7ToMoawX
XOcOr3XzkhOKQ+puvP9NlimoLcDCv/wH9VKOWOLNq4MiXzQ4Qn1dGjD+lbP/10jvslesFhsmctvf
L9iLPTqIhpYwQ0fq4ELGULM4o+8S3/ev40RH4KgJi6fjFFqqNjDMVvkepVMjnJ15MLFbAzPTGscy
3N0Q2b1DpQbmo99udGMN7Q766hLd/6CmcCgqshNLuvT/n0/mPiQx0ewJdqq8nnaOWGKN5x5luX2t
Jvnen8lfMpCYMpVMLnlEceAIvqxJveLg+I0+FGZu0DyQOpTPoChmg7sdBfxz0i++3xoHYvu5KDFc
dcmYrRUy+8RXxSA3eIXQKuEVTcwWvKFJ7p1+P3DKNA2AMMUJAZ33F0eSP2RHE9jC6L3s1dK7XftF
BBYbJQdhUoiDlaBCouVe8RTQVmWEULGHcBFT7Z70Z5mwHQZ1+ItImtWvbWF+Py9azlY6MnmYMmnn
xXmNPfPHXAXieMqWtL6+OVrfA7WUZlmQc4yrpYrQ+7tBSNTZOxiYhnsaodadi6sE7Jkn9+sD5L3d
OsJKdghvPsRDEZCM/KoeD0xdVJqoq8wBhxKKsUM3SXTpjiVbutvw7o7qIXlsyLtZZjSm2GCZSaj3
/K6M3xkb+JIuKWC/FmLSX9G/MmS+iDsoCfaZ0/fTyoZlB34IJFBMhlavU1wWb1h1NeNiQEwaY3bK
nz5p/VQPH09up50Qg/KjWBRdwTaj2XQqZMy2AhXihWcDiO80aFSLNkaeSi8aRJ1E8GbyAeGE2W5X
CAg6awbOQPnflLWH9gjmfR9GMqhWxAHrIeXejGut2po+CzFL0XZR12PgRPGIJVCYY4gzPZ9mjKA9
wkJSj4d/HUPukXBmzeEimrZ7y2hqzNu1ToDuChg0ezTTzb6fh+KONk6FimnUr/SGI7GZFVjzmGkH
6ASGuI0r9kWvuE6Zh2KUNcaGSGCPIpPPaCMlRGRbLJKYq82zllpaa7soiVp8JGkMbG64NFrk0M8d
q1O5P/FDCo1x+kBpcHj72q+/YVG7PcjiBD1BOlysbOez4bb2uFOH6D7tl6sym9zRTFctXPFRC7P4
p9KMB+aOF5xuHdQaRU2JYyXRONjEXkcD73e4vXold1H7/ucO21LiCeHZn7ZIhFU3/0YqkdP0H0PQ
jJXmJAhZImwrCffZ+GwTwNQZNSAl/BuLyZIoJrvkOqw8oGYXy77HFEs3sM7QWIoB57AO+ELXky7/
0AbmKQ1MP/wjE+ZKCEpukPIdIMss6O1l/gb8/g//IvSJYw4Bfx2iRH4cumvdyFrPHSsqn3nJ5rEq
AAA6wAmh69M8cOj13wZCJD2CKxlxlJzRgGKGNEoVkqYgUwlF6lRi7CaNUEwuH/R9QQI62T5C/xAc
F6Dcb9beiEhOA/6PbXk0hq7etwiAUhpectmPYBw9Fk4khVdaQX+qElRGGocsDv7WL4LCRBpauia0
PEQJvlm8hNKWEkRsX8UdNmcPaaH5T1HMpO4R5Ng72QP95JTCo6r8khqIoiKJYWGyIBAKnBC9NPS4
Kt6Mpn78mth8PuDiYbBiz+AGRAeyiwSlfm8ondZLtNCjMzkQK0gJ8HQh9ierwSXmOKWX3ORbs07l
zYRjQ6caS7X7Yhw0+YQ0F2WgQLi9UgIUGlhkycFdGqUhRTTCstgwtxQDtnkF9kR7Hr2Pn0hvmLcz
wqFKFlonmadg3p418UqFnoCc6wAW/Og3yp5AdCR7ncWcduN8INydCpWOf2Cl9WWLPHCerWm0cV3a
6Cj9DXTk3dMb7egt7LvxhdC70ldEekOMyp0609FsgVGMn1lHKkl9I9nWksrzypkFAl2B7nlfhzVX
GKnJYByRl2+Y3GcQ1MYPeQStBzVqLVzSXZ1gUFc8wJFNZj1WrvAFvGAAEc6XrvkfQbwVU/hd9+b9
S2xj00H15A1kXUyN/AANDX9dWwEtJOAQ2fbZcpZ15+0HtFgUC1KVzQvfcn0HVUV97D5vvwkCOwDn
sJw+zM2DZq57dhoWkGjHuvuVDH+pknIqyO/ik3Vj/dHGMFUQQxET58C38j845fI+tqKLlsFNmoez
t6nbCmzyE/NhlSlmnVboViU0p0xZsTDvEyP/SjQkv92ygKOtX1bRG2bIy3ZEVgg+Xybs+KYaVEha
M/krtpK3CFVCSlQufDh7moU/DqGk+gCGQJxLUEtcWbribuT2ao8OsI/curbQ4mg9VAGUjgadk7Np
YTLl9uh8TAxGniK/gFj2I4/i7GIcWFOMzue9S8PLq+/yO7rUKEkjj2EVtQ/kN/35pa2x9mDt1ETj
9kvUhvzQFKo37OQnxrUVojDzwBXSrgX0PcZ/UVIISKMMPR3OnoJGt55LCyZoOlvvSG14cL4L1+dO
b7Afp0vtJJ1DJayj1DfIr41zVkaWr+EvS96tzXZvLlr8jpxFVDD/fxmZgleNtHEqXV1GLI+/OgNF
5JJc2xLseyzeALU7YwZFEmPx05ls2d9O53rwYtqkRTC+L0z6mtAGUGfLgRFIkL3GkYeRZtUoxfKn
M3cz24+rfvCXlmMbdVXKS0KbwnaAdGM/JT8jTlw4sVYqbiwtKYMZd2fWUDalhB2hAAjfwd8IulL5
54w4uZ4jzMYlbkUWM73yIxVH4c9pl/cEKu1szWSGwXBkJQB2s53lgm2BtuQQ3PyOjxfpo92UdNqK
7WcY0LD7icRcCIcaxnIXMhLZ5YQ8SmZ6zy1sg4RZzOZKk1aEajvYupuNLX3FRFomNS6XP7dQF3C0
QgYgBOJw3H+TupFZTKKYjuQn71smYxsEtjUeeHDLiPls6Sr3MIvk/vY0pUX1KLsTvFLgNe3PrUFA
hTu0Ds6XspTWxjQg8YbHGZwIztC8tki9CweB9RypKqU55RErph+Ldfvba7PUvGFfFBDmumQ767AF
r2L2Fg5i23NgqsxKRw6JsK4Jgb4jbLMza20SjQGF9BPUbicPMNlhNraLXfhcXrPxvjCMnD5l7BFf
KOqU1SeSLjo7uLCAwITemDpgh+BXQhl0YfQ2xVM9PBtHieZEE83FE9f+XGoxvmtDZITYN9g0V4T9
eKShmu7Fyjh4i7Ja1ngLNk4IL+wXTrDiYfjwQ6DAm4/iC1QXoqcLXYGSz6lTeg2w67W7PsSwS0/M
sLEOjLv+22frVRDeB+eepxSBBMP8THBfQgn8x8GI97gcO/mBD/JchpD0N29XDsUfBMXvNcHQ1khM
v7QEUjrd42Itp0oUDsenjGqCw3GT/UxWEAS/DQNiRrAgzVdBPGZcx7LiUqdvsUsy+PHFMKcBX1D7
6i1H4JTklWmeKMp3DLZ5cIHQkmcRjW9ylVnjRB6F78WsaEsJ4dSCFfmqnvhrzIZ82p2HnrmTOPzw
9OgocViRPcElPl/3ostpoICsIqSYPz5yPSXncd3FH9g2Wflvthg1fPEsjS041C6Y+Oz3OKsdRFHm
AKS/c215+45Q1oKpfpEJCZGzUB4BxU9PDtbDUMcyKyeQk0ey6tBRBU2lFESghY4Uj1967siMQF0H
xt+kICuiifDyqYqT0S9mZFVmW1dazmSl79VNy/qCITVUturwtaIzzxSyHukDj3VV/4WvROPBRFW2
7iNANnM/hTdbAkaiYvCEprxl0i1xz3b0LskhyOGtyZrqTnw1UnF/IgWnb5B7gYGflQeJn+6f0/Bp
Or5CzSbxYHNRMTHTpyIp6z7Wobis19d5pNXBtkI0WOs4AmWiUSsBminlgn5axa+leWk6fKkrXTmR
FmHk/zxq1rAI7mLp9P3TPuz6sW0zJMLIwjMZfavZ1CAEwAnojD/7BY1BRirWIcgyi2evRcYldfKg
32fp8T3U+0yz7jWqSYRqyu2HOad1rTCxl3hNXwyS3m8e94DQ412EXaCbbgC1I0o8ntPN5HmQTUZS
CteuSY3nRjZRH8vY3uoX9KzIgzIgn+/H1Gh9Jn1WBi42osKyt+62O7vGllDCJIe3TSmmJukmTR1a
DhNwpBPtouGUZm+0OJYoSlrHJuvhNHR362bjyoYytjuOkU0DnfJvDk2t7ypcp4fwxj8escg/bTXJ
MQthX6McxkaPWF8KIajKtiKwDw3tvGsrH1ZK6vkw4mYceG+7m+Ecp7qLAXdWStAf0Sn3QDrK+m8T
FTZZBFrWKBFBUH/l4jdr612plq6XxW8CuYFAXGItEQTEpUOAnrB3rrDwakQYEqy6GRga7vpF0jip
jdnFHnZyWjChuItSoF1aOhn0QOgNLGgm/hyl42XACNOkBrOgBUo7e0Ym6Q9WUg6EAdIkuxSBu/61
/ZZ7+MdTSEjGHJ43Y3+mgDk4LR9rXczy8VM8N5pgqaoveiUmAkrmWoxABIf7u/wVqLz+5bMfdQvZ
JfTkjbD+q6SpSVu4vwRq6vHPhFk5ZtAFhuEQbkOy6byhTW2zhyaA8hG1oYlPyeyp+uDe8hAD2De9
0LlcbO7DGePQJ4ZGApIPpwR6D3PL2NHtzYPx9RGy0pf8hwT0AO4JL+jA/p+FBdnwULxiN4RVGOO9
QWyXe0+sEVxnSfFgxENjkAuqUH757VwwAOIHq52n/tOemtvaKpetDjHNe7EkVg3Bw+jhqfgoADN7
3zNSGtdWPVqdULy15nPIvaybhhMQCt92A6RQa/+1CSzxa+dqLCiSCHDRXteyfRQNbMAuIAEMmHJn
EMJ6gVa6idAUA6r6dppfa5FrqfhVClk2/LbPP+oUYCAIHtCBnNKnMpB0SYHGJhFXVkUDGM1/yNlS
0fTufskyLtnVQAfUceYkazgYNlNMxrbES0HMc64CU23Oa46RJKitaPeZd2O5TCfVMAvcnFAJA4Gj
qUnO9pZKpeMuYjjXaNQiwgSrC50kUEWw2Egj3LyN/K5nvNJfXB6rA4UJbvKUWs1Hs7MrebLp3gym
kd4DaDg4g66s9X0HfXS7z0CLd2DmPnfEzxWU6zZ+UcYmDEqhrQwfB66jbDECU9RBonKNpUNOcvzX
05/9mLGV9SN8t9bOWnjM+Ewr9FdZ8LKi4AzABMoiYRhHGABGvG+e/jAk1+6bIsBLd2U0hUddf34h
J4bkRlH18IirhYUN9uIgziF6QDWtrNIIRJbS+MtRdps5RhSb9/IdlnPEgRtECxq4n8qzMOi8WnsU
WCJgKKuAx6xSCksUU3kLjqnnmMxG5Iwoy4gGWmyiDbnu+x0/Qx2exMzk2qgMmvHx0otDeURat84u
uoMbj6r0Gt08U2SdiE50/GvgJpMnYLqnBdrubjzfm8ScdgNmeSf/Jq725U8sw2gpPh5P/4akIxmf
RhLZZoaQjKeV+hOCQSYKT3yqK6vtWWfhtJEpYD6bFvXxv92yMTKHPHwjEY4Khyokn9xulE/hVd+7
nuVWprqrj56wf4KV6Ud1MKckJFFzY6VLxx+Neaq6fa5z6ce1GxXCwkyNIEuN+LnXeVyNTlxQkOoH
C2fXGUQjyrqv0nZeLsf2Siy4f6yAbSPpw52j9L0i1+AdviDT7B4AYebVDzWUA8Ua7pFBCA6Sp0Fn
p5vPUiyof+kxJWX23OFOMCd6Q04rIjs/6Lqk+36NG1XNnaF23BxktigqxPyJM7sgNAv4+40eyDIG
lB9J7Ie0kVcqoe1yT6GGoiuVE4onyKgtK6H8Gm+YtckXdHufYLN+1FaIsM+pM9XHnWjWku7mEg4T
8XMcZQd+8gcbSUV38q2OiUQnzUNH3po+oi3ylcGQBt6hMPknrpFpaslxhzJ3hiKTqc9Y6M2jRKiV
22lqOzBxI0HSd7kajem63WL6jsfwKyRKDHRGoOjFEs8oW/jmzKrV4JXaYzCUf6EOBn0GjKGAPdzK
lmWjg2X9zQR9Tp0KTdeUerRpER9cSV+xmegGUUTv5RdupxCpEBnZGNrOh36xD9YMFxmj0I7ZnXfr
IgyuNANWX9TLyeio80Qxkrmy//luXVm1h1ChMjZsx+a7vkrvviBMmNmXmGLH+DFvnKUaWGmrlzno
u0jBgGZgegv1aLsFYGzi6QEXet9veB0XPZKJC7dsUYaOmEaKLgTXlebUl4JF5bgJZ2oyFbPjcoFn
t0LpjT06UCcL2W2VyY99Ogg/OMrL5E3UaUwbxdbH7eq1NtMM+IQowBbO4kAaAo2Oittn6O/DTu9E
3gS/4wSWo61UnZCQjMDtuc6W7MT68cyoRnjcVl5AjeiCFl3/id1d1i64zM9FTp1xQ0ieBQWheF3k
jLpypngVPLphIsp10MMk2YTJA6ALz93IpJjKzjwW5IzP/zbC73xZhOJNfWZoupfQkkbBKtMHLgiD
hNlVYrSrTi4+kl01ITj/TCRCZ6tNcQAdHj6ia5O9t4MjDsraoKCnmSNiKPNhwCOyXxlOqNEn9z6I
FqAhCRLRpAEhVT6/k+MONomb09NrQHlcRomUwNbRIsM3V8vVEHSbxHRrXv5La6U1xgZJ9C0jxcID
JregGo1MypzHWfLXSHpP4UkccJ4Vs5rGCV3yhH6tUEcCWX9mObntsZQUiT2XCj669ecCmTB2Rc2M
WIKZX1Sb6IgQEapijd3/U2+v0SzvKLsNZrYgaVDxUVYSOne3fvZPiQujLj0aUJqa/uQbu0pFLYIi
Za5fIBaM0bcpakA4fdzO1Hpity05Tx8+qreTt48t9cVSVs1rloyMKrlqdFNVTHx568SQgrVcsJLz
qMXbRY+yUKfFewaqIPwkAVMKxOaIGLwuXnsk4YgxngcDiTLgnJD47ItQKpibn4oDEJyvMrDWeP3W
DMzazlqsnuzIIF1HhBYkyoa1mn7Nwa9U8+8dVBanUnGAbDJGLYbdn3FzdsL8vOBGaIZfQ0PeNQv1
WdME5Zxu9CfvzElCPJqg2xCDwIleZMbNulIYKuUVkKxGAGeL0PMAfkfocFy0tz3cWdIlMti8i04P
anhzDpgudABSEybrhyhTttlBzz69Kd4XC28lSifZhiCB9viSY47HAe/EsoaoAW8or+YhJVHl5Zy4
g6ylimj3sAeKwssWeejMB7GHveb1bQ6zfF1Vg5Od3SdhoOWI1j4woj06OQMrKV+RYWcgneV/tYJr
xIqyL0zkb2UPf97+8kN3qWuAWzQMopz2rwo+fwnKkNOyGrYgdBMVGZyhkUQOWW/SE+8tbkkw+3J7
rnZ9K0DKeM6DLV51SDqc1whj1yJMNoSbaHCO2jy3hTLbyZD/UwHy4hjzRIFICyi2Lf3WvRX6nVPq
F73LqpZ+0K2ZrYvb+5L7QoGro/7c2IUKs4prJcBId218Gnws2loVIkoxXjskzk2PTXj39qnyPSuL
/9LsahhRxkNY2lRWC2vOBcBnfWsCqgYMNnWkvuB9XHoLISbPXWMpOaFeuZlmU/u9YuICKnYXjH7M
qZQb9Nrxx0XKnD7yRouvD11/2U8HmFB6Y8RqfiDRfslnx0BT2NH3TWhZeh7VS43/aaDFTYTQ9ioi
fzUsveNtROb2Aj0inab4GhLB/Qzm/i7TDJmNZ+9OWZ/RuaPba72ZiX4We41cyo3kvAPAea7gJM8I
WpeExoBApo7gS53aAeHywtHScJVc9tR1N2/jWn0O8Kn+Rz7QRS0r7Deu2YsOu4Q5TD/7T5/jRpHc
antVMsSO3TuCnO1kjZfg4+4WgIdWm5GmQs7P+LQG99BlnJfL+GFG1Jr5kaPogf+3gZLAyFJgfmwL
Of6yIYqC7ZykmoVzxyj0Ef58URpZMMNXb+Tt53qn/g3DiOtAG6PVXhqw72TlebC0ctcVsHunX8Zb
1iEPrGaYMMnzeg6gZ9UQvgJriE7dvT2xUDOnwy2j2b5JYoOCxkX5faGWGFYxOljKtsamXo5lELa1
Am0axsKkO+m5KqJCMPGSFiN8nhA+t4SbfZdQpJYnMqlrM+LdP1hKyVzASvZFixiOKwacyn/0ab2k
ibXX14bn66f3s4Xmru3I/bJAjOCOdyt9KXA8urDdVNPlLm5ZgypmSi6KtD5i8DgovSyVuqGX8w3I
t4c1cjvYoYm0bwlTJGC9VTMF9Zldmt6npZeus3bWzSrtVffrqq+LEAlIAyTQU/VAuG0DJxHqaYni
X7EKsdtssveDe/TOC/v3ecu7kNtVCdMdd50FHJOKKQfkXfXySmIQt95Ckrk2k/6hgYCw3+fz9mki
Rm93Qe0URxxgxPoWl8NMIcLiEMeA16ZnwCiLAxJ1WsCEYIZ8kCdgoCA4VnEP9I+NLIvgg8USVFxx
+22sEv5g3qbEqZdxNYAWmzMJkrrMsTOHD9FtxbDz4iUDdsG0oZrv6iB4wtnifQqN6shZNH+z7W/+
Jm3tJRYZuaVx1pFOg/yoOOYJWTUTVChwOo9bxfdN11k3/DRR2QeXFh79nO8O26AhK2Ou2iuSTLVC
GzYwLIb9o96e76W1ot+99EW3EkbMUHU5IHt8TjI6s2W0rPPwp60n3s+p8FXZPtt6LqUhWMPLt+f8
tck15F9gXWwt8QzqAg1khXb/g0XRaEkjhdDZlg+Jhl3/6fn63U9DsU9Vmq8jnsF1Y9g0M3PNt6es
eFNaHI37AWYzzk/PtJYmpbLGher9goL0Cn2X3CcnZDsDRPgRsmA16WSLI9aogKiiDQ6+1wZNJskG
VL/0+S7pyjTAUphYiSkEczIg/XYsFPqrumkWsHRe+L6tGKPCbm2eJtvXdaTUdsSy7LZoH38k2t87
OzZY050g74upQdJ7lBZ5tr9WauN1eFfL7uMvWgKqSRin0/+e3M8EnzHA6l3BsV0jPaxcEz+mJASg
M5PdXkzeW3esj9oqCgWD8bcbaev8dhce+wRBKwWSuxH5SxeaANfak+NykD6zDIMPHRmrMhhof4sd
lYyKOgYXwgiUQ/t+aFkU2j21In3NMga1jUG6UoypZcGfmDS9Y8gy1WGWzJTWJ5Y+elX+MEfv8aQk
VxYU6zwZCWaP7Ce93CLfR34aiA4VmTaJuZ4KjncspR2zQAInttnmS9NKfhTW2BuGY9nJ1r3IA7EE
QUvoKB6FaQZZ7tx1p9UallO7yp74PyxXP4Em/jmzPqKH4MOeOs/bWzJG9xnQmIIu4CknLJWbF9H6
pnS4OFHCg802qpV3rm09QY0iLUll3gvlKuW0ow3mmRxGd57m/0X75oaG9CQWMI1abRzx5lW6HR0b
xyMXuJd/rlvI3rg0QW5/jGKLkhb8+Hhkhug0I90BF4md2RqzCvIzZYXYuFRf/3cQbmSpCwtOHG3o
j42KFyxgZGvjZKGstRbh/1wC4p/VS8xqA8u+8qWbzhc5LYfjv16kIJyxH5PRGAYhIrYZy9Rm1ocd
GMtLbVh875rwSBIOhQrROEPkQ0usUfbkcnF/5G7oUdJkcspmBeM77FbVXKHXduvlLNTctvFzfCic
imdd82pBuiDRp3rKGIFJUaUlRQ5sU3+ZiudZU9I/qBvVrqDYjYe8mTXuXUefXm4z2ej8MwqG9svl
eJDpfmVFm3hvXrM4KGrBP07rQw8k92Ya2WdluZ+OWGQXngYwU2wGTrWJJmM3JJmDK+bai/JKG/OD
5p/T4pRBhs9tduLp942rQivcRqrypt4oHqNvVBdAABOEH0CbuQmmHLPgBLXEaEeDBNQPxEM8m0aP
DDP9T9iceDvFlDGY2yvFTTF7sLGfiCbTH49NgW3Mi92tveyLA7aWd7wYvEkLkalAsnQ4vR+9ETa+
PN5N5+OC2QbnWwE0soceHHxqFBMv6TFPrkPbaCec7VvdAjaYRQ92shaoMzR4HGwctvwvfx4N2wAS
EhaQDmmn5Czm80v4C8AtjB6m2vE9gmSuEKJpSiu81wT2VGwYdYq9UBHq24xhUn2EYX5hjwpENyD3
3042qTdKfhiu8sq3rj4HF8ePn717lAUmns3qcMot6dNewCZRFOLX+YSGIfckbWNOsEtZVNywYg4a
CnZ+DoH7Enj/G7An3kGklsTQADubVTAvXukBvn/tHzPMa6etKFoYRzlrgmGUAtUjrOjO+CQ5r0FZ
EgmM5tG+jui8tX2RR/7JtQbFNt6Xr4CVDpQ1FQ3b/1Aw97VPURRPRU7L4+shAsSD5hXNyA1zCKNb
jPZbIzdWdrXdY/I/RoFzC8s896gJFp3MrOND6N44t9A+yjckTy8SmcylHoLOls/mTSlJSQmjk33V
+Zff13nM4wdIx02OkilRp3GOEpRwrOUecEz8bn77xJqKozjpwtmrAmUYlyiF/oviQLGv4gXhPljr
KI3IYlyVm4vFpn7smluP7X77l/3Jvvd+KrlZnr15BkMD0FLMf6BIIhVhuyHG2xImXz7Yy0HYIH3i
N4gOf4bO/xSVflGzuky5J5nr539aGDgs2ysAOC8GFwZsQDFAp6nGqzmopbyrlbOWFtgK4OB9BolF
QUHQ+Kz742pLRirDti8kBAKP6ouh12+F6swBGG1dvcmCo6xy7JPkXmrpg99Xa9/4Q//xd9YWL98j
rr/cIwBxI2a7o9FRreJNB5F0o0BMW7ws3g23kT95dg+AyvApIk9Ejf/+9F+BEQe29q+fxIKbywl2
GLiSBOzEaeNjhTYBQ0cgbi3WHHHH6GN0EQIY7p1XkEBnobC4936LBEDykcFzpp3rRmo4JqngtaWB
G6DiKzbKaeOXVmHWOPz5GndrUJv7v4hV0+UIFATfUDM+hfoUO4KG3yV+klcq+cI0e89juU12eJr8
BVuh/bUeCKik/sEZtB9DQgtx09xSJ2VpjM6nSFonMGXalpFY1akaso1O6i8AycP6+jT31mR2oS6O
+Ip4H4Hp3JCT7qxzUH+LIh+ITiw43r/GbsIa4h5HBWkAPD3LxYk5Fn+IgPsMXL44XPxb4CoxoIK9
mNvhJgrDmfnjCX3PwLrPWYQ+2yiCcNpe3oB/MztSX1mczbTT4b4TJZwpaMbbJf43TGQv6ARV8FV+
iC2U+zUWH9AEk6ORzhwv0PtHN4xT//F4jPP5pUAKWpo2lzxFhHc8O5Ziqnq8bpLEXO34z3OQ+PyV
aLeseLnQLARzaAzfPnUv+tbD9cclauwqvX75BkFtd3mmyn6Lrk2iSJXCOPS5YucUkRwHY2nI+/OQ
5P62cgWq8Rrd3fyMrXyM9T8S008HVQyY3IzgZ0xzkCv7LbSCDZWCCGsmZR9Np/A97WE5fJX54GSA
kEZyW/GGeh8AhO6qsN8c+2WBRj0Mv0jI+2/6DCVwbwdilmW49lRev1X1EKgo0IqUwMjJJKX5mvy5
RaJalYrggTYdTcd5d+tAUNbBB/HAVEfK3hYrAWIBN0WR2popTqrlIouOqAbzqKbio76ynfALh3+e
KF+TRoaekXXzfIRM4cVTqWAVTEj3nV3uA6CDoMySJ1lNjK6n08JIADOY/R+0A4X+SJcFsCEQZZ75
7tdUmc5GXpi1QvbiBmBEHo2O/evcwlCOsfNgtr8qydF+2CFcCpLS/Cd1Xv4r4zdYdP0eIJTDOPu2
eUKk6bU+yEh4OLSU5Xd5/3QNeBK9qygJcquQCVO6pGFbrzWnAnKh0r5FkbzwKfdNoEYBLTlVn3zD
0gKkWdeO/T7DmUeSsyH2GyfefnwiF6gZgSCHBoUHvesbg7ygUD4Q9wX4LpqpqaZStdQYQHfCRuFy
S7jGRrAYcSiVNhr7t/mRAioL/bMA3WxM8NpE0cm85x7fCblImfAp4mVk3z4Y1DEw3W02I89pOgaN
FEs4/l9mna2HXzv3UzO1+eKGhlpDoM2JDHMAmXx+4s1kh98+9tt6ZSkYh2Clviyjg+PvdpG2LPNq
fGlYXBqH7gb8/9oZen18pecaEq2Yi8H24geNMhDDac7oR5nc2hCjPVyFINNv+lWL3MkSJizk2UeI
kgi7wlCRuoCaa+ueVLyoRzjfXC9qlautprSxwiV7yaiOmvhe2RHDmZpwoKjBgyoCO9mOnC3deLBP
tlTixIGSd1iqxgH8P0vYCK+oq2YTyyXf29C3mLppPEiwfMaiBmlSNkqGUVr6balAdmnIXVXgPxNY
YXTosZeiR7815EAHf1XUbLlwF3apWZDF/YM5Hhps1ZNfkd+62gruyWc9pIK7FTevc551I026n109
RXpMFnnGNhtzN+agjv5D7fPvVs9EkP/iFex7f48c+UT7pfksQlJ8qqTMQlxkgWSqmFixDiyAOYIb
cyaO179f8cK8AOK4+MKUF+VAqiJqZR/xI2O/sybbF+6lj1Z91FOqIcCo9rWYPnUl+NOGIcM8j/ZN
6hjiGCycxLe8Rn8St+fVRHKJHLPSUUSlK10RX1bKrOy/MYJVNIl+BK0YGuBPYluKZ6hBG/IF1Z4f
sA8NPvxZt9Pp5P0GMLxruxkG4zprqd7+PowYI6cTeGn3x0iGbOob34Zl3OCCJa3t5Eriu7467Oeq
pcdB+fYXNqUZ3ZnMmMxlOpGEj9HhDOurLiwArTWnWREc0nrwgsKYwAw388Rwp0GI90WIlYdEcsmy
WkmijuvFcQn+jvRqueos0g5n9dmXQpHn3SHnA4YBF9c0kOBoEJQxcr2TVJkakl6lIDvoL4N04FQP
BLHafD+byXSmMTTPV5rcc88/fhEc75nWxzMh9ibKmhOUMaqKBTVk9NhaazY+zra0T9pLaah7cQlO
3yrlR9tqHnZCGIRKjn0RnN0eexJCGgwVkmfGsT2+xTgRDOPmoGEqcDfs7uuZlXQmWoQaM98pGv9x
Zzg9/cyCe86ltVpqT/XYY5CgnSFay4r/UAq8sHTpgZvOUTMOtcVw5eW+qxVKJg2jIdBd3Aaj+Zfv
kinHEIxDvlIjR67l5AVwx/QN73VjS4u0SihWhAnU9EdX07/Ft7A4zp4Zvk6K4KVGeDNZTruUqkxd
LyQXaxBJOqbJuLSKVGfBXO0dcoymbTohwzkSMpv9XlfkHnXrTqgJReU4k185P9UZcNdsnOizkatz
Weylgynl3bYSSYtba+Ct4WEls3rJnOQi9j1D1tik+C5XD40TAZSHgDPdPUSI32csgWEpwW45xXzP
NWBxShBUwlWlzd7DUJ7HwJo/KR3n8XJb85mW/KwK2SlYzvCHLUWztR5L7LetTu3oztvOXb4U/5uz
BNvWd91NPBI37+068/jC1HQhvNBGxAaPwSbg603HkkR1q2txcRRs9ROe484ixGG01fndBxgwnTdI
MUzxOBelCAQ9vMtGN34vv72wk01mnHYYeJRVZSe5SY1fC549YjUmiljT9vewRHpDz+0uaU1ij0bQ
eAzvYKAv6ouW/qV+DuaclJWXzlasNpDuXvzgB4JGDSEIbBmyBTBRDpExTNlzjPLFexzIaXZ8Hqhd
xfqI/nT4eQrDZIDWxTSgV1fHh3feCJJ01lnQCQFfVGmoXCKiqzB7jnQG+SVaAO4mllVviMBbpiBT
o5drP0NHy6dpn9+IfOUVZILDdwQ1klza+HlsAwEre5eH2wwa5OxuYlxCHGwaJtjWVgmbWqSiafdk
b4n3dGUmru81a3zFAG0Wr36c83Zq6c5k3wBULt7qt/+ACzNrD04Kde4ccbaTlNTboloXh0HgEXYG
ri+EUWEANWs9b/CQZb71CAXwYKtAZp7u7TZS1ipLbIq/CZVWfkCsV0iwuIK8Kpncaf1uMwPGsNYg
x0YDGDNVg6i7dchNFne3ijfBE27uvAeuLaFehuGF7w3DRGylMd39T2Glr+9hV5G3nlq7VRsXp6/5
lkzh7lssfaR2L9ReGCwPOCyUpLqSSGMXXUKpiTj6EcqBjUy9GecsuS8yjzCuTEwY9mBJGIk7PiGW
350hdiHdtWOyKkYXuKZCA5ohKgzT/7pYnwVX06X+RrKjOR+xtJbYL7TKVUGNkO8vv6zgBEEXUsfz
OIFtJ2VgzfG9TmlfxEo4vPLeDsL/5KsdCdlPgjGWYPC6NHuMxCVMQ4VyEwiVSLsoxMMH8oVnZIFf
smtzyqFAODIFhMUm/YChRN0CbvcHmt+lBtLY03F/+C6iUgfYJmAdHane7X6R/Lx1681uIPzTJK0S
C0AuqKipa4E7pR7O0EVuh1FvYPcb5Kqdg0bI9egtp7u25gSJtVQ00h7Jku64bmEKspuVUHDzHbY8
Z7O6+wi8qXejguJtheatF9BwEp6y0Smv9ELi/aCod+PRUY6RuJKjNYD4cqj+A2Lh2U7q9BStjlBr
bJvN7OWbppkITZzG5hfB9ZRa10bj29O30swgc2l5e7KXjj4AppKVTiHNwLacKwg34j88ZnOHi1el
ky1IDHmfL/DfhQoPYaF2/P58cMycPuViIwCsA/in2T7e6+v/poXA4uaRyBFvev0zGz9ok4/qelMb
0L33RKwFrFf+sklAmsUzu91/hoOBZngPQrizTEdNea+oqSF74sbuuL+7coJEk40hT35+z7BD3cQw
PG1Edu3+EXcR9B7RxJ8H9KufLh9hVWC4G9gFe8n8MVCr/z01n6vXzdJLmRKa03p/r3olCGFjVDuU
4rBis+hlY9TZHdDKFLJViOAh0jdKrWr3HFxEq06qr/5B3FYajtkAQtXrLUsKtivtdcZ5Fq6gFFbm
X+lqEiopOO1TD2vjZybPd6LRVw9oeLafAdqSkXvzP3yoyn5Sg8oxIFJv4pkwxU+xLqNpNfU99o2i
9r/U725M4TGxvjDf4utTbnf+tflbIqZbUbDZL8lOCZOxzd5JuL+jZ0vCwu5wh9spOrIZ57h2Xli3
O2jHAMS1W2GKK1wKHbhscBjGn5pfG/nU5Mb6R97LJVJbZ/v6u4IDWywCJevNvwAdie+0l+qXkYci
fVWso3fgJrZr7VM4gVk++lFfjAio5oqbgirgsOWL7YwESP58k3n2RbOWqyhwimmrh2PBuLUpp8a8
Qf5ZQMknnxlQcmybbCeYPA4ENpHhwX4p4NGcoku8s/xrgA+SoDgMV6TBffSDiyR7bHapnFwANZ/x
yDr5gHJ4U1o4kvFgFrjQMOqYe9+ZmnHcV4OJvSOKUaART6nN6BDVOVB/Ij/qCzCGGMz0dDAK/TpE
M6Km+ClJFrajjilQGfSTvoErbzKOpgwhF2xdPpt9p2MQNIFT+pYWya/6ue89jJQ91QWWzmes2tM8
7+UsgrqC0nrF0AMHhEWsRCH7ZAhG29hPpEJFd4c1NM1XTzN/qHUtbbznXr5Hb1pG9//qyMAUCfQL
SGyHhxVD7enfvh/iQRRot3DUvfmrRTeGSd1OJAExQbT1RBJVDtSv+3+16U+nE0oG2ZOiR3Xf29Q7
6Lem2r1sOqLEjFYJs682VOXiEETJ6iHhC48072987i4qC9kGMg+KryvoKBMf4hYaA7OWLWLBuPuR
FNKoy40XN37rvYAweU2bpf2JQCBDh0OlmwKmATWvwZSv+oUa3NUidFmyAIiXZEHQmCcCzFOtnA7W
1Xpmf80Eh6MZA/rGPPXXDEmfyN/hf1xjmE0OcsAb9YKVhSVspoiyolJ9ZRLT3BTkleX+xyXdgq4r
zBBDORKxeguFX/QeOmHO1BR257QTllpEA9KVqDxQyiv9AIMZkxQLfl9Yx5pHh8TIyueaNpx8bs4d
cSpgaN1hMeNiJAdGyGzRRkDuGlS7k7htrQbjwzz34nNdQDcSvHLhQ9HcLcgF20aCRqbddLRctIa5
2Gexpoodap8JE/Rw2hqCIgMyze0cwReKVED3h/aRBQGGRexsL9wxldsh7nM9Ehudqvea9d/aUiqL
jro+zR9GoHmXrQlBj+dWOpDSgY0p3RkuuK3Ox5nKU3ZI/9g5lKdB6GW8FIqKyWExTw/vmx8pgiQI
sj5SDbZW9zRv0iv9YQ7qhDqcwdzRkGCXDc8LE3oQ4Z6q+aMiJF5hZeZMKFK39Aq6xpRPJwRyUyuw
O+yhR4pSzJ4HD9Xc4GtiJ6W9D78SPlPoNpUMCUVPfW5IfinSr2VfJWcXI/Mj7Q6xwgrwj0redB8M
zrtuycu3hYNm30Z+l8f9TForH7ldf3Ov3bpffywvL+1NCZ5FK3VA7DxMzs3nQE1UbnDPdK9fysAY
ZBetD4PbtPnLJz/TkeDxWa016pygxIir418mXGwI8sQAn0KpyFXRIAR/YULbGYP9yyQF+dlQlARe
hKhVzeySFNn15tTjohnJDChT6DkrwpAO7uoky+jIdPV5fZCDXPpi69QPq/lNBC5j2vmRPps7dlGt
emrjnClO2GGrV05aYOaNkekqpnt/ajbDdtVd6jUzOlIewCNCMQNySbQc4lD87gmZH1xgh4YcpQUD
NvgkzYwWSn2+HulyjmRnTslyejmuetTJiyIIFe2tv1XaXkpi8Q0sGm4aLEwNn3s1p0IgmvC3Kvnw
g2HYn1h5NOtLIx0eULm8zVib72jI7UY239+2LElKMBBUfAAootn/RQ0UCJJkLfPDU4T5ejH/Wow5
ltkn7ZO43gGvjV8ReX780gq6NAsoA9M9QP/f5gQEf30D1DppoAyibvtGfFbWK3APj7lHjxnlELcO
KwWEOscx5hYCFX2ws9OEbiZXj/VOWA5itZDuQzq/3irLhqMaIERTTD+/k4oCowym3gxNw4UMX7cN
S2RW8bKnT4qxj/TL3WcV1IAtrQ84nKxgkCLHyiMN6Zy18oz5XeI0ZPJNDlPqkagVt+6ZCVuAXRQx
vV+udWvi6JzEviwYqGiGzcAhbBWQMKPBqKeIHriAWXVjxSQqrjBbnUPw2BgGnYegZmqIlKNX3q6k
cQlYuTzJFx3yW5Hf+OY852FPBhC0nQP+4CijsVoQViBOzf+TqfbNQLcLFxH5kaKkw8OJdpmI3UIP
OcXbD/kowloWGTdElaEPDErRKZgflUT64moLTI0iP9oiRXQVvMQXzFDLryLwSKlDsz1Qau8aBNXL
SD8mnaDn8QbHWGhjhzfvJfsUYrb5QFeWRtC1J+Nn3M2LtgUseLqe0aA0mGabTD6cz0dvhunkZ6pw
mmfsaN64L35qlyy8fN5HNmstrRpwShY4y1qvHtYD7fyJGGsxqgOkbkhjNPwZlMtLGn1XsKMmAa0u
GskHCuBkyhW8sINPsj9xI8hQzGb4J0dtDbQwymGyRoUMDtk/bQJTOrobYEsvHIzWR8GTF9oCrO/M
gAVnHKsRdmrljozkSFUhkmW4TzfeIy5WV2f3k0w1v4tnwhwmTZKOHSDreB3nyuZPEKgULc8dZhFA
pOYT+816EBEuYoAJ6u9zxO3k5yU0vOXhmYgcYr4ZH0ZLonxxwvibjr2AXE6RlWNG0WNXFPq1+CE5
4JUitN6IRY95GR6q9xdJg3ajuZHoPZdYy8YpsUa9rxOXf8AcqtJw4xY3kXMqlU0VH0gBZNX4gxWw
QHQQ31UOEmr5ltWPDHA/Pnqk+eSjkrxzefGQb8gbRz1ckokPc8saEBqnRxwaGJh/eyU2m4a25X1y
KMdiOeBKvIfBRbdpxcV9M0bswS0fP9xtYVtk2hI9AcyVB53XH4LjByR+Z3YKO95POop8uOuIU8jg
naHKBd+8DmQiYGf4mxfwc9ZPWfUbs9o+VWxALeN7jzlGTius0jH58XCgDKw7d1wBigzvy0daDHn+
zx9bEuIa3KhYih6W/PJ9+njYbYPlYLNI05QqI+2g3e5I6Z8gLefFu/JNkCXZLs47bFGVcQ+krEgb
YbDWsek4yJxDkXmDcDJPDXi+CsN43NBxM1UUEv0MkepenRQNJ15zA0YRh7bCQDv2l453RaRbtq9w
4YaE76Q9WvFQiY9gLs/M/ofxewQxJIwCgKUUC8BHXHlZi9hJ1Wm+BxvJlJu08cSj3TG+ABQZoHwV
wUpxFdr8F32gG87SlH37EYzwqa3MgtcOz4fEcMrbn/3k9qTyIIh4TEODv280HUavM7yHwOAdRDR4
SCv2vlNMP1pZ9DiiRFB/YHiWzNaJ105Qv443djMBgYSr7Zn2yQ74nHfNQcEju4k9hetFrLryNcy/
aDRpmYtUaSO6AlrP6xOKG7BmXEs+3h+ROYdwUzNptLAwPFmE8PcUksmffGQOgDHfdc6qfKAO8T5D
OrC029Lk6F/s0IljhiF35brb9eu71SW3P3a1P7n44A25TisSY/vZsGtFpnr1A3pnhwNysWTmMnfw
b37wifpujlblebUJMmxEWK/d2BVHG+l+VNt6c/0+AVgTx7PPBmatnzCKmgjiRkrxbBrzIRy97otP
YrYbH8Y8MEbzaQ4Mq3t5g48IgrJi9Sl9lS77XVlmc0w0sLm18MjBKo7P+T2gH1GxcippwHXrbhoD
sWqC5qShr2aoHM7Q1b3OLVFZqQEcNBRoocEsGu4uCj57NAA+kW3iOR0Bkdfd2t8it6rgFsPvvs+t
Orc9dt352turpHr/KDHjc4mL0kc+OfDGuIeaONb+I1jOCct54l22OqRB9zBg8vyJM/jL1jA6o2Lw
6Gn4JyIHcL1szIIPqV/wpIALmW9UamOubABp40vbULYAkigABZr9MuQKFh4GG0COCSuo/1q4KRYa
f2AGaXfI7PjwajJpPGJ3DOE/Be2AKQdA/YDnhGixox09fV5AjZcWH+D9zC7ix4+2fOy8VGi3H8n6
AUWvevKmk6mQGSfI66wTGIfTbwp7mgww8I4V15KZlKyVNHFZaaP8tKRzcebM0Zt2oqhCA6ZcGgGL
HhLns5+f/LlGubLie07VTrJ6tm9RxhPGjme7fg5pXqOix41aXpxhKmvhTav4ybNuzHhR+IxbLCs8
FnrmJqOUvPOH7HuA+0V/ya4zI15ZapEdXcHmSZlVC/KeEFdgNXEAqA5Mb8h/Yu8h7Nsrbq4w19MM
xKFN0dHi1e5BAaRyi7vMs8ARbyrOv86t+tz3BTJUeMxSusaTl3ggFgZDIweT9IqD7kUz4Im6Tqfr
vzL9GsC7g2QhBhCryMObqr8AcxSpbbx1BmHB/akr1j6wRsaLFRqzqyZTcMxaCtM+m4PwcMcWJj4G
H//Rhk6gM1KOjIPVfTDmxILbmu+Pbjhrzes9MX/3V/o9NSmF2cp1H4Z1XiVDD3Tox8frxYt/kAed
5RBynrrs5ArRIs1nvn4zyusGHRZePPyrTq/qxNzRqtome9VqakpP4ZTBx+UXS6iWjAJ5HI/TI4G2
MOdn9QRRl+FEgROLhTRZFRE4LTuvfGLJDSEYBqdrVQjCHSPDBWDG3jIXMZN/Y4bztitYmzSez7GZ
v7x3ed4a4vYgJMGAz2F/MaCJtEiy8gWRPjcOoiG7bfIkBPxHLJWeDiqLvlIHB1FC3MaUtAwp8QyR
5ksXn12MRAtc77YX+VuPVSOoOqxCDs5RinhK3iERKUTZYSInQTaFh3Our4Hn39v4DjSlCYMHhxEi
CjMmPxofKH2ed7JXENLU1Scn9tb98pCFk3YL522jPl6/IBGIJSip+1uSajlXg1LsLYFhQ0oToBCZ
SHbqgLnourk3uTSPJn4wbYHt14F0jnTqR2bl3Fo+1zEmbvF/17BxyM0poNfxlLef+8cK2NOFBVxZ
FgUj+fEDXiR0VetYxieYC+5fK2P33Qp9WAumP5b4q+STjn7DeoCa+Y+ZFtmuKMrvgFIv3Eb2lIeW
fCPuOG11yT0GKlgXbl8mIwEJAkY7DThgKy0lRFQYG/4YYxBmiuQC5JJXFw+6UhDHgWtRYeNo5C/L
QJ5G5TItXmtZ+HenLrHuMAP1SWmvV6Nyp3jFYAKNgE2I2oh+daPCOUJxndwKF0/4i0AZonyam1Qe
zHjcZ/fZa04uILH5IHpZjFm7yMJJ/ZXKhzmhUQNJINVfQn8LOX2SctOG8a1wQe15yAM4/Mwv6Pd3
0Rk3GtPCKansDmjOhipaHKNZKBUWW+IVYEDvwZTV3stkqpoqCfIJEliQo7bv1UOR+djZAM3ujm+E
Rkqe2NswakISJiyZiKqgWAAegXarMvTvXgGUxuObv4B606Jrz7TlTeb41PVyd9gvh+ZOUGyuM/t2
StnDyZmMy4Ir4lxRcXvFZ6zr+tKjnRjLOFYapSB6LkS7J69dRcKnyFNOCM9dKm66JMh0WnuKXe9Q
w9NJcrfEfH4Zi//rBe8H+AyHaRwiEWEfH4c+Y1x8eNfidxTCesl1Zx0H1LYuhPNJqR2TwsIVTZqS
aM2rPOJIxFQF4RI+qzvuJ3K2YtEoMRKytqmz1G11RHovFqjWMxFxvrOiJ2cNuLv6rHO+j46b5jpg
yrsIkdHhC1u5qevszXXHpoxbw0xjnx2NyOiHLUk/2ZhO4wZZxFJxDN6Qyc7gEhNalZdCXlnAi7aS
q7R8a3Ufz7psdGswaKi6mzZNCJQnSxe47dDbl3/iZ8FPqXkqxwA/i+ItT3t1d8FYecdKY6whOhiO
1mBVR/osloVN4U18DQjDx9c6qa1C0qPsToyaDCBG2KrIm8YAds2PRDiKk0ks9hFH0Ubcaf6zoPTj
oT1qm5LNoAl+bOjCM0XzjsFm82sl65stiXfCLpailSRnP8MrHxe1rJiOHeMRer9tW+bqkyCmZ9Uz
2XtyqWX9SMmRWC0lzqGb355yNcO7g8+ZWWrAffeR+oB+IZxzF9JPviwkV5O9RPm6T5xHUNQaRdTi
EsqokID6Iyexpf1fLhF5caR78FaAUTlpWOfRV6fRgiv6RYo4U5pajRLlcEd2Q5K5D5008yuFa370
hiB4//q2Eq1JJGCHiSHzKfKZAHXtDEB+qhro6xne8o/MRw4PUatjIegVbugRDPyG6p8G5/iayLkN
3QZB6M/iET1JjOSesvZEQLhFUdq1RTHbzeVnCvYR0WQoKVL9OuCI/dp1wmdu4+f6b35Jwn5/WHPc
wt4cco0B3aa8+KCLZ4jy0DvOt/QS4gV9UwFUq2LaPp+MoE3W+4gFst7ZEUW1pQ7mgz7s1+rGukx7
fR3OhIFW8u/sFxc6ZOGzuwxPaBX5KgXA5Y0QRztBeEaOU+BJsJRUa9LVcCw2DEb3zA/U1FpC1QrJ
bd+MsN7ObCQJieCgJG0ek000UXUmyQgZFyvmwJoyk4P0jA151GR/RDjshfjJy6JOPznu/0fLO6ud
WO2A+3QMMdn88/Ys9oQYfQAlgycXSMal1ttqgIE0uGTn6DHdK8zFSsIXq/dWdJKC5f33M745DL3m
amiVH+mZ6gyyJNAOB02OIM/B4x6My+UA0JB31ov80bFhGcCSJlT0lazj5a2JMMTeSH5xlI1meqp4
klgXr6L80JwhS9eEIGHVd4bnbmDbtAJz3a7MItalTqD0zb1u8RjsQWVjWO/mllGxpV86MpNKbNwj
9UN09se7ftTA6q3BmPdtoxiWOu5T9ybaCJ1vWY4BQzy2mEr9S/om7vi/Dc0w0tChLCQa/YH1PRXV
43p8YA78ISTYEV9cCAwgVCe1xXiYRy9lXCSm2o7vR7zZ1Pf4oWKTCj352t4l5Muweziy/pHaNYEX
KCNGorUpf51UfFRX7Q0LMHJeeZtWjZpW/caxXIl29TP35Cj9YkCYDvEEgNCLpIVDNyOvU/WLKXes
GuOgknDIqqD9KKKzMKVNa0n3dtwhgXRsY+vcOZ/SEN3hHjxvzvtOSW55jY1IDSZ9SQMdqmDi3gJZ
bYXvhDU1VJAGzMt1TH6gnkWymTG6KCJjQLYIhatv0seDyYSlUcBjkdZ8ZNvps6YMjfQBWhnLVTZT
AJdFy3gvgPL62Tn89bUiL4ER/iiUIkY47k4Eth5WsCaGiRr4158hBAI6inTTiCi+LG4qdSWoldim
7jLIgBTeKN7TAzyWfDuo1NdvfdzqPTx9M5mh1m5rJCd8MGv1Xo1q3qr7MD18lm3wpuJ6hC2biX5v
lNGAHtsIhdEruSsWsdFSKz9rbog+Y240aLjT9HdG3X+ZN5g3x83SguM1z/FW1QRNKHOEbTac6z3u
IYDX9VvpWqd3V7LRgZDE9zlS6NLQuaCAyzvO/almH1rZT4G7DqBwSSlLSrEefh/RxtXEUTc7So50
tDJR+ihuH7F5qcbjlDjptESy9LPPs6Y+sx5W4vIC0jfo3YuSqdfvilLHRkpOJZI8NjfM0NIqRJBc
rrmeKnlfJEE4TWdLAVy4zllZoNUxg1rcHwss3HcLNZg7dRDchtIOZa1L5+gH4P9/3nQnxbmcMNwa
JzknGHqkr7h2KPSIeKhDBgaeC0PjqjgCUNuBrQCKDGX2E2mKA/pFb38RdN6i0cTHDkGbw5p8oQZl
2IMi6E6mc1RDQFYeT5fiO/2pMR+PCxWR1+sLfqm1ZEt76x3mufC2hH1+66k0aD4iM8FSRy6N9Qmb
ft9WzGwAhCSJ10olbhptkl0PhP23G0Iiex6ouIKuz/d9CkEdHY8ZbAyoVNCaYOJxl2nx837A++hP
7rvac2ZfMx4Kg9e321OkBtjkaZR34kxiKfwMGbRguzXQKPexqhwMuCeRWwdIfr6pMLjo/rM1t7fR
6z6OfDusNwz00+xDf9EjxZBB3T+4px3SpY26A9usTlFJdl1brZESqyDt1NpdZzncRMzm26BSiE+W
/nFHn9lMCnizo4GyjtIufPKRUC0qX7sXxta1/HU8lWmNHPAnwfBMfsAaDhtdsV8SuPB9ABLCvDU2
kio8QhXZIxFB3PX8Yh0oywzN/eIvB4+81PFNIyOfOqOFDGicXIUDq+9B+oWAWPJDk2pCN/Mm9Sgm
xXjD8/xor8gh+MzZ6HT54d8BGnDamyMfkMSaTlwAxm/03p6vZQwSX18Drhqfm4DOWAPbVdNDxClD
dMaebIi+3hJBJI6GuIUf0Vk4+1frZcbFSHH9OG85mslzsfm3XGbs8LViFDuk98+uwlU07N8n9CZR
JgsyNZPGRHtoj4I5MG7tF9RBEZTGHHv88Oopj/SaxKCCbGZSA8qHKw75uMC+TT1YeuOMlLwa5g8Q
U2NtpGQiVxBFMBs4tHgG7N2rHHBjO4G6QzOPVbXXQ8tJsxGlH6tXhG5AO2FX3+wmtvJ99RtuOsD3
ORXThhFbV9ofrr0191Tmw+N82rlXD+N42blBpAz4s0tbIBCiHCrjZQ3Jzrks3LeW+8SQyk70ZmuJ
ROnWpynFHegZiWcL12TyvUnZ6d/6/j3TunE76ExkGcYtfXRnukByS996t/C1jznNhhGy6nBeB8iS
dkPXddTc5rgV/FCpzcbdUuuAX8ZJFvtiVO2dnDai7XTvahJgE16TwWI3erplTFpUant/TWg4jPsh
YGZ8D6mRGN21hq8CU1SHvsV9+02Nfj6aOQ8QrthgbA7Wc5RW6BT/PKuu3ydr+BNXyPwTmNIhNeM4
xkoeCPFR7065+lMk0unjLluvIOXiFhy4008RME1QI0lVj89ZXl5L3tpoeXLh2I8uFlbolceadBlb
TBIaURDmzfUo1ub836uQS6h+0QdjI2S8Si4VF7GBsgoFRNUid9FYj8qqNMrT4JBQz20EufZThMAX
r4Yv+zcZ+UH4kuEZ6OLAmMSkEL1Nh/DE3HWZ+R8B+pUP9xL8EZ3AREJ0hMmi1/kVwanc0gyICjKf
X1eHleF9ta0TtBRKbl4n3wM2q2ibWSf5HX+JmUkXN99zXKpx0mJrK6T1jTXZ9qD8FshDks5OHIQr
Rvixoi+81HbNQaj7R4T5m1GSoFhni+zzydmXOZmpVSuZv2/wFMJ3jFOh1TuVtMfez5waf4YhSRT8
Ct4UvmmZ3MvlrJZfzaYhyjoeVFnORK61DwbXeUwL7v2vgNMeKoUqtvif4990R8X6gQH4CBA9iQLN
ZnUm8UBOVlffMIDTzhrmhXoHNVA7zJ5/8vit9qS7IjRXSSN2Mr/lfwtJkWznBqrcnITqegWQ6Shx
seVPOOmmHIoSga8EBqpFlbqhQNuOXu2exdGUFcm/hZg2NRi/KTmO6ZW7xt3X5XfoSAXHDVOZO8AJ
AYFvPs/y2w1U6aCVEIU1qSaqFWTNTGeOS7E2ZcKPksV11dS/AvOziGcymObiEnoHrIi2DJQYvYen
UNXeHJSkZvp0PPMEz9NTs16VN8DvoPG+w4unLrzM9MiSwjOBWQllykiMYKJHrPcutqEHJDLTE6+K
1kcj3XrIYPf6HljZn7L9IWv8wfeBLwsHFjv3YfoQ01Rg3F4FnU9gFFwWVXd9nVMpCyyGvGC07095
VQqse0wb4EUxGw9RelE9mGTuO7QZ7Zpjxqpypuh6op73QRHcPIKVGTz5dpnae1+0coR/XDsLE0rG
WRILVkGgJxcgqE23/aH9EqLVecVHXDul9WZR/OlVhp4HqRL4PsDi1h/i0xaqz9DYjYxoS3CCIuvQ
akWGVyALGa97ed/uQr2J7a5U1u2RDhIi0qLclQLxL1l5a+gkY1aHhDngL3lCjVao52x+rFt1vx5c
6fVn8LD5npccUu8kF6JFN9MX/QHM5NLa1OPxdNAL1J4OtqLWnvBdXiOgTZshujPPnekfsx30uaMl
zpxc7CVXP4KTCPN0kW5BD4KscvlucvmXefpS17e4DvqlT7W/2LdrRy2m6wi91rEPMTpEBUCwUaTl
FlMh9HQTAycw6Vz3JCViMpcYT9rlqHaUxzEiG+knVfF/LsSFH04MtCjo3Xyt7t43rrPtQEEZb5sl
hO3rexRzKf1r1Sla5QWwAnGaNKW+GZ/d0Fyw3zxQGbOsOxZZjJNi5RbngqrY1oe0Do/bhUrMgOol
M5K82VC8o8AuoZiXfVjhL23MZHofbfLsWnFTKkLpLzBrH9T+adn1L27FiMHDNf9C4Ydyz8raGX3s
mD0AKKXMB1vlWPJbyy22abDprwv8JPD05dtPYnFrPSrgVwRlNLohwm8cPHcdkxyoGM9XjxX+eSGx
D1fVS8gA3keB+akeKMd0J1OBznfPuc+VTccISV9gk+HGON1AC3HzsBr18AYUONRiM5x3bouiWIoH
bI7e0E0i7RBz7h7R1nWMR50m7TbYZRxm+B16TGX2J8QNjn7VXPQSjdCw9L+A40AFlPmh/iQFWaRv
PqNKko4BhtszX1+DwhwO6Wr+vv4P1kbazjvOT9Vl2yQzfe53xMZ5V5ap6sN0cCV1LQAZQ1s6HhoU
eQr73aIDRRzly/Ilo9LpH34Fg4l236++DsTWZet8e1rIFC+r7YbmY5vYFz/4deKBn3rIoMkLZT7y
Yh0CUWLBzU/CG6BYq23wY0Dqk+ntx2xlXkPoex5fmuv1oLiIhzJjhUMxfzvItNHOj15y+feyq0M/
elWhjakNTXNTnv9ke2Fz6Cl+ax8ZYFOOv/xxaACOxbq2Hu4g4fXW0RffpyeRRFS2/puDjpvazSQA
8Rn+pgsToHJGkfVoBR3Iz4372nVzGf1yU1TDXDOeMwp+uTrn8XRE0PacLSoL4nQivXOgX51IGdCT
isLrPSRY3KlgYmxHlX6j/it8/RcPt7kjGhWlM+gjM0Qyy5OM2WlEDP9QePAGmhCvTavVhtEQUZx2
k9th5BLW+wqwGdxVlsP+czdp0OtqYKmFpfEKrpZuquz7WinPtgPjRIZvGepUD0ivlJPhccyxP8YU
koheE4SKbpJFFu6oCtpgSpeI/K2Guyw0LkK+WmLKtC7rGzHjxYo4ssqbPVMO58P28RdaOLPez3st
evZj6tWB6aVZXkTkxRcwUF3JJJqjNpjGnWNtE1n5DfLpDoEJeToSFAAwK9vvRC9lIRJer8++DWBt
qzS1LcB4U3vl1+2HbUysIM14Da2PjZCWKOeZdcNkTJsGwAmSugXtgygVMFhKn7w9kuUOQ9cabTh3
DX1weed4yKFLHXQnUtBoJY4ARZQ8Xq3G5a4/wzbotaGtWa5cU+r6eo/FELoF36rkglmtGNT8NNZl
WlUdrl2AI+iQ4H8HXpZfgyU6o6RgcMMmHlVuV0OqUBistH4+yeqSghMGWNFWWz3uikoEpzkKkPxg
6pe8sZXqtZ2bu4yGRUDrApyL9AeyLsQGw+9WiUeRzny8iKbVkLZlpyarWc/XOl+WO6M4eSBO/Fxk
0F2/He+Fw4HR0yJjsIpnyGs95qDLjDuO+uXBpar7bubqM4jkJ3olpt4d1d7lSJpUhcxoTRz3b5Kv
fCyigsctKK0hOx6chhUAmxIEZAXRmuk3soHN45FOgasFb/HDZ1GP/2cZqNaGIA4dTh1g06XLAAjl
21Bv9fTVNWFdzZf64yMcZn1E4/wFXUDNrGUqz09ZzqAGCXa5IpL9G1S/OZ8+Cy4aYnfKFyEmZWNy
q4zFccU0SUE4zjuUFUbQvAM7+gv7s3VjAOZnKDG7OSKka0PzTjPvFCZAnrU4j6EUGrqXjij/y4QE
slCTsHZEtSeTqjgkw59N2E4zFrdrKOP/4aMD4KRS2P7dkp9p+9ShlylSVruN5GSCasLSLJMKu1Rt
5/oC0XgArCIr9AygcLEAFUMSNCXd39+oy7RblLdJJXNNGfeGYDLZhM+F2cxdyFheVsEDrj6ZPBjI
ll7Uez0DRGeT25dag+Pwm2Hvhh+M0xd3un5+uL5CfEFdNmjJqhyEpWmZgoDiPN/EptbO+azupI2g
AzH0BvniDkC47M4WKoczvMFrPNWhz5pO4eX88bDDAbaMv4koU5AoHoolweO3lm0IHjJ7VB4Nhbo4
yvG4XGWAS7ZW3PNlxiGarjoNVlFcYK5rYrwhHYK7RNt0Fzku1E8YOEcPrCllO8FxIXA01YK0ouub
hfLv4uaS/+lkO33Golii7mJYlXCz3TXRaQn96RCpDqWT6Pru77E9pwmojcxrx0+/cozH2VeCyl9p
E2QRZbDoCcUd42dIz3OL5QHx5QQhR7B1O2NB3a5bYw43zhuSZJv+wqDT2iydzUslTzDqB2oQH0hi
jimgFhJP4wALSMTaFhs1GmDfe3uVRPhgz1vHo4lQYt2FmBTOOa69jPeLPWCD+lS5c1pIKBuRsh9m
lABmVUeWCTt0QOt2MDQAHYL1n/7Fxe4PBibnclh6Xf01YcqIlyEcyJXVlihl/JfqikowNiEk3K50
rz9O/ygfOht5zoE7/yc8WRyot4jP97Tp+HENWQUS88DFEQRRilAjQLVve+JSlnmXCgC4vOtMcNea
KYfJ0aERa6Zkj+KSFNKTb92watsxDoiTRM6nAbf7SNNc/IpFvsAABd8mn5MQe3p0NOFU/vhtttnu
c3R8tm5tiHKyDzqz92dkRhiPDqLnxGcmNjCN6Dqsnnn7G04eMlzLxcQkmJAt0gOArKaqXS0t4/9d
+wUSZhJ+vE4szvRLr2Hj6y3J6vOiC2c3eyqC2r89nqVEtWpTRx9puDCTjQzUdX/gIw039hlDCmQU
L9K0OKZ58D4GkG+GmwyBZC/UKuDYyQ2Vk2XG61ZoogYMi0Pc6xtfnD1Jhn6q5KoiF8xRvQldYKpJ
HplOJSXTd3cIsL7Vy32SYXKthTBmKo6TC7O6Lz2B+wBcCuI83t9MIbHNvD3Z6eYfmVT2AWwOdrUr
DzIHInQ2fq2Lit99kAa/dsq+Hajriq+fxpPLAf9KBbFJpD3KUT6gpIGgxqI6weYwZvDCQAcK8oYQ
vZYj8GWr48SmhKBJzZ3ZDzcGwUF6bsLhZN91esYAvexaid6+4vq8UoV0eEZGIaJS1XVmsQhTY/I4
VDokZgHi5mNblVGZe/dneTQGHrFaa8Vca7ifLQzcRTLhfTPn8dbH2D5seb1vss4fr9oGRhHltjFm
PotbjlpXdPLh5mE8pwCKCJnmX3ux+aJ91yOnEdeTnMqLntzLxXxcfsy9lc22UkNom5rdEcOZa5j1
Dd70uKsaQhy+u5mmMywHF9IaPMAiIxoAK3qbmoS5eWrXS6RDNxoIROClpacLSZszqakeDQoW8hVH
R4ixENjW6u3zu4WztNpbHAghqBMGlF/8ZKQVu9IyZfly/cwliF2zwfjn1WRQDOI/EAg2YLVDdRA8
b0/O80t8fSZoGS1fhMp2/D473HLUW349jn744MssArZ9l2Qk5q+2dlqtXaZ7nuFvn7iqFVAMS7R3
MlSR9HQZtry95wIYsPF2ynmVwLBr77YqKE0jI5DQErMDw61yKL8BCj2uVcWWFD8924l0h1K5DFUv
8o6F31WaF6npGBMHDnMbDTUeGvDCmJ9ARkSGW748rDDkNEw+7YtLTZROJMAmzm3aXCL7dlgSHdL2
nCcdBxCdR1ttBODnY9jbTfT63idmAU/yEZAv/dGPJqA+ojByI1MvyGWY8sNFaqG1UDB+o8i0CnK7
NXoGOb0B6RS10i72OEIgvqYyfMzTgkUjnOr4AH+o+kpYvCDCbXxjsT0aufFQSHpP1D/mU5jKI2pD
vrbnJ4uwiLnXkHDdgZkDpRxlYv71P70k1xmtKoCYgGtcHpFTUYHdu5CasIxDmct33yKVHlcB2A3+
hD1v6CCMXxZpX+qtWtQsuwWmPLJCnoakBUAByjbsKZykHdQ0+EW53js8jJwtb1mjyW0DmE7fh9wI
aybX0l9w9YadARZQOVd64DcAK/lM17/1cY7KhfViSTXdiQCeJx7q7dD7k1EDjVWhhZOazVjqQEgZ
67GvTBqOb9mEx5YdTpvNiDriuwP8qlk+4smK8jytQO/oYfhg242+dlDv7OG0HV8zP5H1S7heWJNp
bQnJtZVcIdrBcLkdjFj75xKOT2dafc2m0Mzaezgek//diIcawnQKAG2omdcTQxmcP5wXo2qfROuU
vxaK/fo2wt/SgYKEECvVJM9fWQAkOxqAJsnbk8iKV+eh2KkpPowi0DJ9K3KTkXLdvCbl/0Z2FwNW
3pSUcG+oL3ukb985ZuV5OyJD/YkDVELkhBimPrXUpMD/HDYN+vvylnYPLSv+aTMQJDDBwyJq+ov4
OVYYrtwRhR3ryvmoOchQ7+IXm0L1lGb0UQ58ONiNdF8saWuir2z5chcy9v6lrWiXCQ+Da/QsNujc
CPHUwKqa2t7XfeFoIWz6UVxfjEqef/a+zLWSDW9u+qXLEvxzr0s9vpCbHh6zR1Lqmlcdz99HQZ7h
Q1PO+zjHbdVrZfur+okBOTJM4AuvI2/An6aj5Pun3egg6+8806WA6xbrkjpYF4zaPK7iz5U95Pza
gS80D/lb06DRj/KC2XKckcEniJeNI8breBy5lelcmU/Z0JeaxzUqwff+ou+U4Yz8Kgo/38IErVyJ
dUvo3Vb8X7ogSk9QXxuXW0nXulht1gkb9HkRQpvis8qLaBFFfhq8TPEFnSmW6HjZeOZEbBfG06Sj
D6f9t+ee8kPQBn+upMIjvUCmt0j3cwG20vpIp72JJNlG6xkZ9V0DWfcUJFBKHnpy8iMQZWSCDotJ
V8f9O6O/6UijHjwvKmsR3ODO2PZUxP6mmh3EtmlJeWBOQWP6V4x4a70mzvdzUztsJ2cNiOBz5h6w
I3zmY9JzGEOAWDx+YdSvyyAyGHSkBqwH7yh2izUz4vLQZmEo9HkEmbaCriP6O9fcSdP1lGY4CIEb
TCcJ5gfBkRtQmHkptUqQP7NYrYEySdRwhSALKa25ie6IIoLq8yroygkkCmYPpN4A4hoNMqpkYJoa
d7Dn7zJ6F/6VogCu9QbvRRnX1DSpBdkCLZ2HDnbN5Jf2aihT56d2Sn2wzbvzTfjkHtkaJq9MLfY+
UX7T9ITM7Ymi8x7whjuXS75Fvc8gIMTc9W/RBY4SDFGOfFlZXPZBxCjWkbpI+dCpLiH9cxSjI6HK
nFeYt1SuOBs/nem1ELca2tpzAMoZnZ7arhym4njrsGCZ910rzVJ6851WF02C+v7gaoK+XHePddch
d66CU1csrhXXckORCcB2mTzeGJZpOOXkmtz8EzU0LZVpd0qCDplPZEGPfy94Iw+8MAp2RwOWTOD0
fzIIBHyJlvlymQ9cLS+dHne3TGmd0QwdsJFAaK7DaSLuyj5Q98r0l5LT523g2p60qNlzlG3S5xSz
x1Mtw7fWGones5LVeiwHMsOcnpZ0pAF3AmT6UoJ6J7y2xdKSz3L12RvwipU/sj6e84aTyJEStQ22
yNF7QeoXh3TeDCAWJQDHp/qvu6vYxIaDU4cofLdp+jQNZNABXtqE4VmegNKt/a1wFcX3LGd2kXFI
thnHdHxIqUt9/oBl7/xg1SDXYAcYOFbedYKLeaWPtx6XhWegkos/0zcgeINquf77+yez3Dt6HSLu
Ej5omLMK1fTNzdVjzIA1Xni8m+iJbzeLwgB0UxHXbQ+gebUYfcQiZL0rCOBGkenwVKAUgIDBgfLn
tb5pbO3f2DGfXM0VmeM6pkecv+ilSGOPcRpiS6Mmg1Aw+dexGl96rfEaVnmccw6nxv0lVOXuLbxK
09XvnMXtV74Eytd3QaQ6es16UHtdWTDTRrxRrsXTVqoFcYpHEgkRCBa1Tv2BKyGCZzUrCJXCaeWW
yR+N7S0IsxgVJvROv6P5Cfy6jTbo4IfvxwKlB4CekjarE4KZLqpqOvQqyqb0tVoNqlgZItJf9xJt
EpryH/7HWWwO4IQJsmOxTXd2gjt0gXPJL15a6Qh0WWQghk5QNgQZXEaEDSN/jnZe2mDuTWBhUfVQ
JPneLCVIGZOEe+6k0G+uKAYNvyFYlVDNKL1jXT3yb5FdBSKMRobAlUOG/OR718tD/OjNiXrh2dwn
2P1i+FJxj5JKy5hDhTyII+9+sVNDFM6I05HBjtLiueWa4uITFJc6txcxXOIPAyGw03poLEgs7pzy
Gg11pRn/Tz+wqgLtvgtqD5IBULRjZ99bWoHNzqCr1QKyPFYAgSNXRcIESEoBuuBCpgOL6el3tHOb
pLeYNKVntgYtwTjHRiPpQA1khrQkn+nNsXELiJCPl6zsvUYGcPT1LMo/aSIzU+1FlYHZa/MSKDfc
g+4owGDeh4yIwipJdctKFgTkNVSqFfjahs+D3DNSfiG/xqt5vgREMgjSIyLFksLA+JkSsh7xgba/
ojPTB6iEt6tEen17PdVzF1PIu4AF5egYTiZxC3xrYqvK8DDyOveOb/TSFFEVbdggaUMQjlJ/ZqCe
sEJMGx+7eFpHjgiqB9vqeNZo92yWycn8FVb3A348+aVJDRWzVMpvq4ithhdL7mcrGbHSgPKXbefL
i6pEiI2lJh/++hUdyCizvdNOlbS7NWSg2Kb+eS+z4qJ4NP0tyNA6lhTZJCyJsXxzUDuIFb7kYYSt
vu3U+yHLMbTiDL13ELjPCmemqcrCcxCZqDI2fD7sCoAYK1znBgQwWrTvtCLJO2zHOseTosKK+Tbz
/vAtU/XHT4Ddsz+4e+AMRs899tQIYVUrnLlHCol2kZru6mMTPCl2ZZaJe9WNojUSpVz70AZ9cujE
QiiL8AqXOQNs7oEjErWNS9TG8sFxkclh/pe+oxx0ztkX4rpxi8ypQ/f/DpfYzTZdQDMCEO0MrFcC
cjfrq8aVX8EmKK2X9zmzHOqLj2IeStEeSRDJpIEiXw8xc7cT2TWX2TD7pjBHKRKddNDhaDK2M8q+
00sRMb4BgoujvNDf9HX8rB5Wes1U4UW+mzS602dnyTbq37i7F0+WzH0QwaSfp61kWlhtEFW8bvve
H7wQApGgzRIww4nGuAkZDxhm5wNxv61AzRZcq+Q3Mj9QQ6JdIiydo7EkfsbFnpDcB5CQbVd/124Q
MTQrX/qBUNQCHSG8Zs0fE5uwXcS7tKHwVafw5QAU2/RCsbwZW+2TA0VDjJvl0w7+akyaNJGT0gYe
0UywuP0tM8fTq5WJ3DUoJXBzIV+mnb9nanF/EOQD5cdWrmiRztnzVhzFp9D9Atckv4fWESYJuv/z
uJYUBbJ3tdb4r1si5rPV22B2zcpVf3KID8h4sDCJnWBDPOdMo5pU76rW9Lm6UkS2qrtvQxKt+1CJ
K/m0AB14zFkX8eTQrMbGwpS4bbT8E9HCh167kVzETH3vIZtsAQKyQtM7rdECIQuWmlRcyQj8YwQC
R54XYPGZiuFb9HiJqwggLtXagYqVKsb8AjVPoY2QG9kQk24wRhPZ14Mw01bI2yRYXQOHbrC0iqSO
EiMJTbZ4EgAdvERmL9L47kCWT34tnPeZ3cCYG5wB/AC4nolaW7d9mHFpHIqfWJPUuh7yPLd5Zw/t
csX2G05uhyhdSHvLkV8FT9ASsOuIQkcPD+lpMD6fh1WylMNZ9/KA4y3Rx3P2EKzCzQHcg+k0nEpv
yaKpPehCTB3syNF9jje5SPRkW8/EqU/nWD/dtEa/+x2ZhhqEGkfc0De9CqITSb7xirWLuogHgvXw
19BV+zWvCdFxfBoyGHAEpkR//52y9GZFOD1zQaxF1FhB9bJ4wxnxUeuxomWYZtREfY2YspJzUuc3
ueel4rRMFLLODc8cm0bPZIK7YwKmnDWi4BUu1fFV7C1XznmmvwDtJ2lBSyMcxsX0sr7FeSqjKWgR
9SY4f20/zwt9g6KdINzS3UgstcjDMjvqzYgUIrbi1V+g5YE5VNpncuwgmPB4YHqp+rV0g5IWPFhq
RZC/yL96sXR/tajINtGHLyJ1yOJNey0m7om50s7Mk7Xy3dKYktlTILiQWwjK2jQEGkD/+g+Ljxn3
25GqkCfHoWz8o0+pm/5J+n0WgPxPeyqCUmmQjjBCjmWck2eUY38cbrvUaBNq2MU+REdQCci1Qtqa
zyCcM+dAOhp96h9tnKnfFsMgwB8z8biVToxmO9w2Q1BnjYPrvqxprYzyBhBwSlbprlRPj86VMK6I
joP+hXmHW+ZIu1FN9NwkQTlFYk+c13GatLNuER0Wvc+AYIVoD9ARgJJo1cnysNgZuRJBrrE5B5F0
BeK7+BG9/+qtuoPf7uCe8thjNdK7zebcO0E5E5ujikY6/1J3I2L7OXULtYYFLgLjkEqn+XGN74Tg
v+ggnx9/yekZLyHjHGWXTL68LeZLHN/5p+7Ogamkqu763+q5hgrYPWIWU2Sc52eq2M08/R/MnRPm
dDtkm/djfxRe37pdBOW5jXzgti95oKNJHq/Lcg1x7uUfQ0mWiVC2j+UoVL3RWsS+HuTR1HBj+EMY
3QxxLycytVcNtIF8CSSTh+ACRoRwlAUJ4X7OJAX0jHzxZGQI7FONeLx48U38oz/PFvGs6OXX+iql
SIOwtL4E2vGZb3Yce9ZScIcOWciApI/N30hDTI/W/0KPv7zC86WwNfNFAlHc3t/fkSzyXQ+LPFgW
79syBF2VcfENTk+IOo7fJsrJmo5l2nDhSm7M7wv5OR3Vp5ZL29Ac3kMR33v4OHRLOElK3ARNcS9H
mX3szIZ+wevw8kM535OSF2OKJzFARj9ZUqitnmR2DJUeZ4YY7fDcl25HhL16uSGWXGm5fogY2mf5
0z30WoroCGUjjaqtiOeabc9a9/OQsSFQVIywkw3W9JTzpngZ0mYKauUQIVxi00/elt4CmYxtJ92J
s1f0Gy1SwA7IuVhGthjl1zKZsjTqsoglqccJ3+hZ1QBffxKXm6NXK8nc8rf9kvGuAtu+63yUFUa8
W14WdX9hf5G98sS/f2pNiNAln3V4Hq21Fz24PQ7uSxjzQ50hewC+JIdSoam4aGnZw2EnNCICyEx9
L//psdKByRGONoD1mcMItGQaTXoo9BDjuVeiKLioS7ZSMOJ5KbwP3YXHVbs9qF7wa+pHBVVFIKYV
Nmc/jmNNFlwD2CCap2MbJFjtR38XgGl0BQILBYq2qEr4GnAnToeBn2yyYkkLzHqED1eyfvutGzct
6bQ1hYJFj+qr7v8t6zikFqUT2zNWTO5jQ6JcQ0WkdUZDDKs8Y/4JlBO8f8lzZfCJ1xmg/hCb2gNu
fXEKd8BsRyC6yaHe2o5OKxKo/auETz7+PpQ9rAr0uyqJV637lSk+etYRoVJXxACVLU6A484F0EkE
um0Tvnc1kxfTlnYXyx/MLMq7C8jeePmw9j2mLQgPcf857oE1sU2Satrc90KVhRwSUwL1J2D9EZ2J
p4dq945TVMOAc562+vAPHkq5EGcqACACJb96523bfzBmthdSC/L+JNUEPForqc7wsa8xlmc3oRsq
+Th2vizBRHG6V5eTAxTL2HKwm+WlS0bLSHVxEj+r30fYfGPSoVZEZpSe2hinGc0gH0ggoQP5Tv3P
J91gbgKeIpVA9iUcia68yVA2bkprtT6D210wppuRypTrjmhA1kArGHy+6dVs6WjKSsnxahsBZR32
e5Rrh4RGae0Ksa9BUre23N2w8QP8MC8g+BiPYRM53QI/l6I91Ga4MhqdUj1BF3jFdITVecwBN1mf
4n9QO63sxfU1eNRMQxXLuetATK4nkN7Jhl9bZPXv7AJuaOmI8X+UItdvhlNX1aX8BqpfT8ScJdOn
eKo3ULgVCjWEtd+bfSZKMsmv2e5qXM16vp/h1A72+ph8jEzj2xb6OXUAJ5uVfQGp3MnQK1AzjBIl
WzWmO/h9hLnmOjejw+nDX1JEbXOaZUiBoNMczDTwsmOWl+D+boHpOr9DOmPKh88m3A5NJTV9W+1a
6HXZcqTRwCHjHRL6tUYhg3BCCNBkyd6FBpxC1D+/3kx6VHv9uj+qPTGmBdZmOi8ZDw0i0BaKVgQk
pnJ94Xz2kBBWoaHXKk9Y0sb1NjdRvKCVoIsqL08PtIb47BsG6Hca4unY6MkpuDyTTr+jUWfE2b7f
qER5Q0Nt6Xy4L6HJu3NKgTYm4s3xNMlFP4vWIPsdv4gS1kacDm1EmutArt+SCOCw/uzB15UwZVO0
AohKvO3YMPm7lQ+QeCLBmrOVIHYzjYCEiNUmmgDEMxCvpgOWI/asB8YCcP+LAV6GYtkqgEVTqcC0
jsF6U4kxbObG6uDRZHUXiR3S3U6BZSl7ceDbNF8sAp/9TzeOb5/gufSkCd/KFH9d9G/fhC4sMY6F
hUctYizyP5nd9CyueEAKF/M+/3R1ZqY91rY8NV+rLrKwne+9E9EOVfj7SUi1kcPVF8Io/40FjdmM
j1UeUwDY/GWHBVVIpJ5jQDBcxZ5VPAAB+CvNHJB1VKZH+VpOL8TPxiCmXk6yyVsRkvXSjxxTqURo
XX2kDlLeQr8ujnkokIf7evq6JmsybXBv0fvJvYodZLjU+YrggXSCj6OIszxw8JHqNmQ7tAeLXO5G
lDemVAhVRugOZbprU4ou5KjU3HgeKkN6hNXvblqJ33RbmacS36V4in/scvgld/8m+17PT3K/HlRI
VfU7DM7FYIpWsoOrD6PxvYGW7OGjXleTeLJMy5K7TiNiVeuS3u6Z7LL6+fySetQT64naVzVfVA91
EN7fN8qKceTeKHaIj4/Bya9ZYM1+NoE499urIRxlnSW4Nqk41lr8/xqZHvxCw064MiNeUBi6iGDw
inOOvdNF31I7XsPVojbUtMGo9dM7RabFz5kE2+rdrCCh/COOKoyChuJ6mK7a4lGNJ0gDnS13K4uC
4xL4CwndMBz1i2dbm84mAwD0AbLbVmcWkwfybytsodDog70vDIXEm4g6GEAXGVkDpmvbIgvIiBIG
OWUdARUhY6COzTf02itmWnXCC1vHvR0tqNN1oJPm/ys8pDsu9s5dEGiQKU70t72Te6oNRSH9TvoW
Hu9zIGAhra6Z+FPf7ChFgaSTal9XH0ecFbUFHI8x7x5kX8KlCdu5ACdowFMVtJSux+Wb9UCS0dzu
Mp6INUy3K5pidn0MulI5ckJVGrJ2/X2zJ/iQxs5Vy90lddMxyzFITx2YZdbQcJLVX3KPFTq41YhT
rM+g4OM/YC45xEbqCjGwWbwxoCXIGVNd7E9NWc9FZVkuIkwQkznb3rw6qTOJyGpdifcC/QYqNQV4
NG5S6XtETn4M5f8KYySHt1kmwR7FN/BMb1foG7a9DPnYOPJAGDflVMVJxsxmnI9c4f5klmDWeZsa
F+N3O7kh7tNCajN9V0WAgoCNKp45q8FsfVrqrPtfrlWZJM42YjBQFFMgwy7oTyxYUfx9RXnVDy2O
bmSXbVMcNfGlLKXeYrtyg/J1idszCdLCwyiFlaoKQJTPvr7TULzX3uRRauIgG2HbX0mgcSMs6PNN
U1Xd+LqV/Mq80LnYCj+mqc3nu6olgbaukOyKCUVNmwHtE/DDjKzydSXcu5yg7ZJNhiP1M80GyTB4
cnMZ37pPMotvWfZjx7X9RU7fUFCtn3LJqcnKjgKwFmsco9OXAGw+LTrU1UZfatpTnZc/YQ1mASSW
yzlEKE7+HH1QmH4axzseLqJ2JdjmnAD+SVY/FPjwProZjQTOFA98mrVF80BysMno9Og6p38mrJmY
a5RjqirDiHMlghX4YJMufGdcmh7fG1nMVvPbAQTXKJTBUGfoPAynSoihUfx0YaDFfv4CPwOrycNL
keiAxP/vUbcCahagKYRKibK92d5GBK45WylerZQLW9p2eGTJT1Imn4uM64ggglffLdnnLFumJ1YE
sqF2V+2sTVcw60hdE2DGo34vPYuPp2dC3xzfn7C4Dg5RGBLogJgfT5FgQZEPSzQr5Y5OUQzYoT1C
odwWec3qkz3iJPwCc0+uLU0a9OENaV4KUj+urF1X+65FHu7ihUF//8KTtd4dwUqCSA/RSqKTLD8V
/OBISpXeKUe9+s7i0HSY/VN8yHn0Wb3aNv9wD8HHBvU6dv/J7aMuTNWOH5IJ68/vnffBmlC7+geR
tP8LPJSQuiswn/bd/GqTLp+A0C+DMHILC8oF+Gw8I70HxEaS1W5IIUqghgtO9ELgNbBogy/9Ko7+
XeHDO6q0lE1Y/jI5tNDYgTPgBV1bDK7If+BfHDl5b+sjpsXV26DK/HS40lYWt2EF9M91mesxgJTE
WPetgfbyrnAm0uADSbZTsW5+wQOpEQe0GhjVbqnUAWXQp9HBJNKnKGUzoWxJ6+apeRS2QAuY5cOz
Vh8ChsVs9Pldx6gaJIPivd5uVcDzGk6+9iHVJRQe/DWXkQ9S/qchNCIQJcFOS9e6x1R/WpWieg1F
4RZMsDodtiqcRgdKrggdp/yLG1sMWinm9U8eWOjjkgCk0vOHvx7o3buNvMShZiYNSnSWHnWtB7NS
N7DLTiPL9/ukC+L+2cCqqLX8jCsUw6tNIJwzpGPMWMyGcVlF9JxN7iuine65KlQ9f88Ld4hfzbCU
jcQVW6ktAgR1UY7XjcOzurgCiTPjLWYWZUkDEmYNRXVwo0SGH6FfQEPovi9hGmcRyKEVauTU9nBr
0rbnYNlqZZpnphNPMJGz40Ko1OC1NYF7fczBfU1HRSoUiCeexM4lZdm202nMomzoDAfV2rIHooda
hWkIRIw4CZrVG89MDYDA6p85Ymgmj5TiPXhvdidteliI+qwwTO+jpSQ5ODVTP6P73txHRba6xvkt
3aTHKf7Tsizk/pNXNyxp8foxIxKN7sXV0PqInUB9t8cMvbClj+n+b4qb5x36RvgwQqitU/azoZ7y
C1GwMG6fyCOfomvp75IjyzzDReckZz9Tt+iPknW+PwwHQCf4m+07yU0/mDFWISY74aL/TM4MxE50
xlc+4FbcB0DC+QIhJMNqbRuZZR1ZyQ06BzR249+bTYP0fGcvWpyjSRVNuM4ca+aBUi50JHWYu63y
XCORWHdIZCjPeXA9OgJF0vQ1dkHJwH+B845Jveg+4N14DxlVke0qfROSn9id5Ul9fpj4Pl4qqgkm
/YAdSHLg0ctPiOJT2ydexKGL01zeOG8vuw27/cMN3axPdYObuDhOnCLmxiprQmYJkF2vdRPWJbEk
c54n/YKvfv6VbjSjquUwO87axQ/CwArBgzRthX/qzfi3m10F5lL0z8irZ0+SMjOqX4x/JGJOruhh
oY4SiyowMp8GAERv9NJTSAJc5fvuJRQLuESf/TOyMHVFx0o8SR8GQNWp0fb1sgqVtk0RZqpOX/8B
jF2thBrt8Ys1dg+n4gPL91iBUoW/YoPHVHka+Tdpc+uIrXgMpolzZp5OBokz3E9X0Tk/HgzudNf8
4jXVNab+ksRy4fhRrZviWK6RZTX5WfaopbiSEz1nGzjf/IOVpBGPokJpzNQa+VM8A1E0M1MTAEfK
++JdV9oyspvAP2vEGVW7GlSlGvLn0hA4HfDv5uwPgyNnFNM0EklJV3DH1KIlZKITzGYo7ByDvpY7
5e0Pj7w7erot0hiT9uKEsKAErDIQUMgVDr083kzPpRG+X1blf78iB0/Ey0smb9khcCN7/4UuWi47
9anF6pg/yKvwH+dqEYf3W4/ECZGp7FUsbAxiycjolOBxZ89MtxQrAXV1a5rGO5ROaw7LUDk+xIbw
rPMWO0JPhPpdUJ1ocVvbDnDM2f62H/MihmczQ9AcmPFzOjPkmV/vAOfkIzmg19sX2hD4NzWojmZ4
7qeKOICXZdvymCqPHgNHkTXR22eyJPhVgAowTs6tnujXCfVxo0CoZO8GtEQsT8hhlQY6RDEsZ9ev
W8HenjiCZyq3j0IU6zT+Ag6lSxH87S+sRUDaQxUr2t4V5fND8rT7878EhkUyMoqVYhLJeFyiWDgg
nvppJCrTbRiH6drPHpI6Lc3wHK1ztG6mCA3A46K5daW0TDpF/3qZefo42CwUwXTypbBQCob9fwO3
/2WGF5ubYF+9TBLf+vQdojK33ctJoJSJklCzvua635YRuziv8PA1EksXU5KSHFkiruTcs4iKKvSs
mHzB+1TvkMKXpBn1iPN87IZLXpzWgrR0HOOtIx+bM44leGqtcXPaZeYdEQ0rWQmvksjLwSxNRjLA
2hfwVepUOvzMoEY5nT5vrqxCdWzNOpaI5MSO3OXzKP1bwdWqrKhTTeX0nxBJ4LGPK7TfGFwe2xCn
qeUJdW5F6zkRC8PsBVS5WRa8YXuykgaTCejCwYCorsJfD3/rfes8WHd1F+hrmC7zhAtkJkqKnxhP
8XPKdj5it8p/V1y3LCvnyvDBR6XEyHvGz9VcZVXgXVxUbjwh5jMJ2HMo2/I1+cbH8grF7FIpQs0p
eZIb9ptwbj993IyYCTivegu9UiwR3kBaabwIePuzkMnVWfRKHaPoCmuFVUzk9Qptn4Om2GQe0DtI
uTfCHKKRuQnSCA3K2fD85/KGwyRNYaE+HnnwvUKfNhlezCAW6nhEaUH5zWlvKc3kKu096zOr9262
PE6cijarjesTrm/Q32224qQ12SoOREH2IT6ql/SNKsfEAwxtNfrLWx9F4l0TkZUr1RQx8ZnSd+mG
f9qfDoUtwqxwv74bLOx45K0Lgql3ULatbgnwZROCfVwIZhTOuJGUfARuSGjg/vuMfiWoHXQpzOCW
cQ9rf2zG/4fa3Cx/YEk95yxgwegvzNQVyvi7/eQlSIrs/QR5ox/ggW4fkIOZqu+6Hyp5Rnryf/EM
zaIa48VJD9FxnleDuVXu9GtQV/MRpYKbW7as+h0mI/uV60XxpyREhQUrgD7cLgHG/s+/unFgm/03
KXsyDPfw/kfOEWMQFE0U3wu7yDaunSIrB/k6Imc/UuRB+84LjOPkGD8FwFuX+MwABGpKQgxBnM2v
vsOdFQYkotvn/+zHNYpv5RDq37WIWjx/zewStt6IoMq0M5mwpGipmvnA2MsKDb3K9hIih7HIo3Cb
+8QAy99Y8y2O2777FpTwv8IFdbeqegA0ppD11QBm+T0KJk2Q6i221UHv14PS4W8ErJqLnz2k99sv
zlwrk9XbxwoMKrqTexFmS7Kn14mcizMJsnBS3Nng7gM01TXu6ofGommZv7wAkg6SBSCb3ePSpLIv
neEBkhpv8xclXD08dIFHkOHJ0nz0BtTWIr/hCJspLfp3cynJLaKeVfDgC1sHYjqCl5Pg3cWG3rOh
LVmahjWI0KbUSXDkDSy3cvM3Qm2XTO2Pt6XfTHoIXe15CuBGkwwbCyXCOfcnaw4Nx9xFapUUWaeY
4xvUNxHeky9QLsRlkcIiVJ06EqV8ZFrUvn/JOqHY9orRLYf596PmVyaulpo6zPlHmNm/W4I8tjUa
t6+vyoP9pA7dX4RxksGNGUWsfJOxddB4Nnv9eGQD5qQQlGMKeuq+leJhNsKofLf/JvTw49f+qu68
GJQbOy2XaXJnC9bCvnzNhalI5Iv8AHhJvrm5A/S0MC/42YHxnL7j1E46X4gJbnfQVMX6L9c2Vom9
x7gRiPe1GBkqMx90uYxnkkkp5kUp2hOBlrkvYp8by4yScfFi9zTujvCe7TOcFm/XId/2W24QAOL/
TA3W9xnbYrX0OU0TUwn+mulTfOy11KnC1j7g/Vejx9t9p6ZKqB+0F2OeqYEzDk0A8j/s5Ooju+NV
YiH98DOtZse5xNq3dAIgnPYNZw2i18YtIzEzU5PHB8BoFe2ZtoV4maXkGJQmidBmN4NmPw+t+M3i
3kOTNlQMskJ3e7ChxVHUJ/DoswzRzaOUX+4PRLjs9Ft1wrDthpbXCoOsV53LaPg482FV400P1sOT
VJNOsGPmk6OR1/IGkMHBIC/KMkPGuTGENyVFCytS5VuQfDH9M+NRSi3ILCqZWhdElK4fVVIQHm6f
ymf9BA4F9hDsk10ZRVYUhHy4GZ6OuO7/M3bnzmUCX1lake6d58TVI7Mcg3avw6yHmSOoBzbjetKV
kARb7yRqj1NvG3xAqHdyAapfLhgPOKAEtUj6uws+cdoFCeqUyir5rQyBDrVmhj1aOvXkRD3i4CGY
nTaH9TMZA5s4FQMGuvAPNm5iyFp4QLSQim5H72F/Pt6XB5wJsEtOP9wG7QSvCP3FwIfsKX/AiciR
QkBGhDjXCyF7L8tOI+j1GATebKibvX3ybTnoXug+GEYl1TUTZanXP3Aysgmaen/zoo4oWn83e9/A
Bv8gbWzNyAf19nCrq0jOGyLiRcVaTB2ety9CGrV0rnOjp9Lw32D5vjoS9E5L/GjRhNF4o0axwPRx
nHzZudXK0nhmTSZeJTt0OzQU88dF+Y8C/QH9Zc6e6Y3+Myb2aNvbKP6yfJlato18218QXbPmxv/P
Fp7Uoa7McjlRiBTgZ/TfhJq+FvCg3y58PGzZuLqZq//haHwFjbLvAHBmUEGl9aAqgUCRMi+tSruh
bILAKDJcxwxtHLvtOQcbWOcscHv7mJfIlKz3HGd14aeKXWAEnQEQMPsQz33BoXXjC3Rn8UtgGfyS
jmbVhpXrlKMI8t+PIfd5ww1I0/+RqqJhWJbsAWgwE0WEKm8h8T3VtPRCQfJXMtjOGmVqz6FqRKnS
GUfhQtissCra/HT5dzC40cg9vjCZLU4J5nKTiwwAiRjA4JHH9oRrxCzbpfLQXKwQFyF4TJYvy2VO
w0UHlDp1RwDi9rOlxfefhfbJbGTdf7Cp1dyB2gjPVXWcAFkkQSIvuaxC/f/aJUDVrZSe5gKoxedz
UJj1CKg4GyPG9h7NQC4Y8w3IfSqNvR9AilVG8xTyPqpr76ncV0FjgcXQKGjZF1r26avPQUDUnANW
ZgEoQVcu6AowJ7yZkZaNt33jOCmT8zRedXDYWQYVuzNYU1J7Pmy1Uo212wA4PDJ8NUrWT+6W8yX1
ihNYhhH7jCz4WpNlXzFVvNG4UoGjHCTl8zNuSfau3UThde8NlDLAFMEsJOZTD/jGwpa0Rn2eJZx0
d1vfeBsVuJy1/1KxkgAxJ+d3FsxtNGHgPiXMg7eQduzjO00DKgRo4YaKIw7O5uEVDhWEd4l6J8ZC
cY+P1FFJJl2NsoVlAFdRmqWOqJWUsInKVExp69NrBkjr+jFJY8kG9ypO3zsq5hKcu8GE3KZG8oGO
ZJCuL5bqkqa3oUrRGpksr0iQHGWXU6aAKeIvThD5ULAtXGlK4J9kv/C0HCDuh2vxEBjPzNjoKdJE
QmwlujW/was8ElPkINBS7fLykYfvvp9c2sxMYFCLfiloLXREsSLOi+PUDNkHmS7K31EBtTk1wXQ8
wEqIoPcORsnwN1T3nSA6Nk+Fqei31diPip6xdztksqBmZ8gycq/4GhmSYuKoj+HqRbAUI7e8ptpp
cfaIJlFNmHP38OeZNOwMCDKeLPgM1kzEwnZehDAT9iZ9BRB0q2XbrWYBmDDNSgvRCMbkKbA8EE+K
HSTTyHlVA7Ganw2DeNuHTaQ8O5Q2bCS/pukFQLEsJ7MEr3sqHV8lIOUlqAD0MGa9vYZtPQtQIfwK
bAeqSlOLROWb4I8TiWmHQkOKGV9jkO7Y9pdUYn/slUoGOMDc8cP4LzpHmdTahU+llimjHqKqSs5S
5+S8jRDEtGOmzgsgl9TzERKrAXa/luW2/f2UvAVux5SO+mZDtKA7SkTTwzDPdbF0VzzIilvS8EkT
uFf0CeMv7knsjmtxyalNvBmrXqb3O4dyuYT+L9cSnZobAGSb7oC4VH8k4/Xel35HYjDADzhrGm7F
l/StdrSDjUgmhSY/AG5YNG3/OoeZfjs8N/g65/liJzVWZyAks36p3287eyn/TckTe1NKaCfl2fLH
I4DnVnhVuG+dnviYjS6svstgQN5mvLJ6Rbl8ZNS+rriyMCsdapUF1VqsLeq3pMFrSFGNTwvkimPy
SL3UdHQeeHceikFOUIez16EfojMu7G/6tZbuuDCIUEgj8oTlhQKnSE6B5dSnaBNEJygHpV3QAJuc
yUMsHwS5ZeMEnsbN9BH/BBnzO2mlzMyhI3jEXGh+fGrXVzb9sA/1o66foKPf8TpvLfIp/Tfc0N1z
y20ntNTACppkxtILPYX4SoOjTE0soNwGa+PB/s4mDCF6ODfJPldmzhTe+W/xSpzt9Y4zJU1rz+mj
qLO+lcjWTGE89r/ou5E3RkEndaJSI/W5kV63NlBSpn/7Dqa3UMd9VSJ5E2KrcKNFhX7n7otx9qI6
pDGiUSdyoaj8Ytpy3IYaL3AHsrVRDt83+rgKx/c7mmTIH2E1MGP342UC4Qc99U+AnLqe79onteuC
XcfHqSuwtCmgEt2CC6Mzw5EOysuddObyJojcjCs8wzOjFuT86rg7X+QdF9qk67MThRNCfvpbHjdb
oPwB8wmTTrCpkFpx41u8GGKZZb9cRIURNlZPLByy9fuSvO1R7slUGiQg5pK37jgm30z+i2OThA1Q
broRm9RZtHCo3EIhY+pvduIMHP8ccLuFKCnfsBqPf2aKdreFiki8mw0H+3lx/0Zj5hNsOeXR6uXt
Nff29vuA/JHUWxyTCHrWJncT9gmAhE6Frdmv6iz7Jo6JB5qXyc8gbapRm978EcTY/1zeRJtvJZY7
pbQ/Vgrwa++/YSXSshZLveW49sTf+nljiMbx3PB4vEk420B2LRru4BKGRxH+X5X6tEl60TCZTfi9
JKpik4xvbhsqz4BFTkzE8hjcZfawd9emGLFlqOdcA98AezC+mTcwQriqDOFeWxYe0AusIBugo61F
qdk9FwVyS7ignETmmo70zO/3Bdjkmc4waD8sBaglJER6FIxa3BS1+DjzGktHTJaHFulFP98DKNi9
MQ38QPmYKu04o+5Jeby2FuGUlnvx24JjqefF2ZGRUb3jYgHS9p4FVxmXwtssftgPQRKjojN2JKwi
IjUL3Pj4J9qxfBVNF5k94q7c9JmwozFdsS7cdE1560jIe6zqGr5ChhEyiW/FklBLaEmmCf72BKUy
/Nb0b8QS/7V+8Qkf3ClTtrFeqDRKp5Yr53+MKOB/2Kp0YIbRuciqeugKN3O3G1OGXiP/ZWetylqh
0qFYQNXayAdrNqUH9TUMoKUMdIzUWkWuA/WXSnv5JgbrSR/84P9aBNCTH3aTnWA4fAkGGWISy/hV
PkMI78EZ4ySwM5vrl8v+C2wOz9ksZo7iPP/MfOWsvmVUjXI9y/5gP5jg3t7XAZzdr1Q76KZayCXk
AnbesEouYZwPyfdC/hL6K/jNOdABr4CzdVLYYlQ2kJr7Bqyw7D/T5y6d/0v9Qgk53pqPo5OkCNwC
ZM57L553TsYtgCo/gXlInLVT+PThtZx/SMfbckLUjhj1NmYtox7TFuNiS17qKrCgHVxlMG2rH5pA
HQsdpP4UeZmUlqQRfGsXMzxOdehz97pd80AIzOHYcg2ZHGVirg7ehR9IAyKEOvmRQD1ug8rFScU1
i170JbH7iz9EqzRKa2U17ZPyA1BjX+pehWnOrCEQCUvNs8JdjQ0+bMEhyM4jfct39/TfFl2vhq2g
7g/Qn+eepzLXKOQqSx0q0DDkn0+lJmdAJRUTy4bQ51zAIYrD7BLcgqUUuqXZbED42krd7ZK3a7ks
Y90ZjT9hKFjPBburKm+VX0YLEQd1PQQVAD0WEnpclzdmxpV4J2WFChvkXWBn9+qNDCA9++RWbOW4
ZTSqxZpE1SmO5TJZiqb4X2ba9Yq8FRPNHvlafgd4kiwposx37PK57jTGv2ucjRJ2TdEMJsMZnVz5
DQseSUACfvJ8TCelEwV6aavHBOGfYMXdLIUnMZLF+hb/4cZLcczlr3QWuvCGfS3Ez1W+dbEzjY/V
COXg0NDD8ESqnC1X5PLRB/Iru9OIrXGattQjxFlPplSmYzFSdxKFkPLRjKhpyCZ9kGLL4vv8GwME
4sRki97MXggFskbWbKL1jYh4/Jvv9eNGRbRx5BKK9WmMT4bwiKipEDYBmgYCAOsE5a82GzZBzeA6
DFflOxqPbIPwB2J26oaCOcCesKc4RY09EUmnh5fcEhqfBiydF1th23uTWPwZgF45HnYPDd9tORaF
kEFdAWDgtwpwEfpY9jLOj327ECYW8Ih6orqSOtTl8fD5WgrSx5RKpUjOebsGJRyS5SYm1DJ2ynQ+
VJdIiw9Ljf3/QKmif03BohzqhaJRqt66BxMyWQvToApym6qAr0avfvOpl0P7Z2Zkee1vP5i+x9GE
0eXXntMp0LH7+H0BY6c930kokr11hkWLsXc5b4x6t916hujysN0YRWDayGKhnZX0UwhOWeuvnMuQ
csLzRrpwaiQEB+54y7ERnuJJkbCF5MSIQi0fmopG3fLpx+RUWQqHvc9G5erH/lI/ZMPan7Tmm9a3
6DXxD6UbwyeSO3qVid3rEmGvjG9auDdCVt7739DE8dFPGtODYgCYzb3D32skHNH6euM/XWYXBkGE
J6tv9BL2igkh+/xK/Rb7bfma+TLA+60VgGjzotz0OtgR6TVw+e8UJonlIlBUw68zgqYyNx4k4CAX
OgXg7iOGKbkaJ53GDO8vzr0Ku/nlVHBjci0/e3kQgQe5xiKHpn1gDoRv6JcpvRfKOGFH3NvD+KIU
dVIblFM0ALPa4hCOTzD5kYjAZvkYG6HkGQLqDIlDTJZ9VYHWhUR1rFH0axtuYzk9HgrdoPO7OoON
tOM/0UceFzxUKwOJoMajuy9KAOpuXnq0H3tM1NwDO2/2VHif5KiwCT0qskFh/IcJ1uepID2Y9+s8
150JLQ0GGAqxPNtv2I152MX2kXpQGfRaCJnLNc4TobGhcrLUYd2LEHp6129x7w/zbst8mBzBBJkh
WB0ZB6CHigoxHGGhG9FxtUbSTGSRYdY3WPOQgw3ZI8O0qANQSBft7/fTIOBgr8HIsXLI/P8Pra3F
EJmqdP4evfAz781Gz86Y08NtiWuBp/xwpfZlhR6i3IOgRFylf/OYqU14dxUoBXgWyD6TgK1ZMiPe
t5S6ackXEfLMNERtNcoolZC4xHf9D2VpSdiNx65G8UdbYczWogjKouc7VJWxBiX8tCBCMgbOyeTh
sivQRTHaU9hl54oiGXCgyxd6m2cAQde+xSwHWH5Ln1/wXJo2qeABnPlJNthqebvPusxsQ2m16q9R
Ji9Lljc6W4ujn36q87QoDeAImjqtXW4t+O0oGcLBBuNr55tYIPKsVh36Fz1mhAi9flHXFiwGLNB/
3UT6U5KF1FPOhJ1SDjOByEJt+QQLfvH2AaSB/9GA1Z+ZEtlO1lSGFJvWab5pKtdwqptJx5tysObf
nFb9qLNFlfTI3u17HTXerdVT1O9rLi4taSgxrggg8ZklGIes2YpCVeTc4Y7zdR53EFbcU3ctBa66
86kNjEnDCx4rQufEp0kPMahn+FW71C/SZ5oMqQWSRniz86fA+P2Nndwe9iXIH56IiG6v3leHDZ5Q
I61tvMOieMZs/Fym7QLWpmJVuXzuuSTLEIYFiKmitG5+OfA50/ajzpXWPSo/aRvTqtrhoBgaY2jH
P1jGG0rS11m6j3w19dlJ7clcZRWjH9TwghoIMg71CI20VIMwLkMzLo8hx4MWIRW+CcOYn9LlgfU6
7LnrP/r8fi+hs7EDlhfvT0FKgC47xnoQ4WNVsJ6kA65qbbz1EFgPZ8dHaBLnE75DE3VbiSEh6K+y
o4aPP0JkfOACoMC5U54jaMOhpUghzvYHHIswHeDZQoqsjhDAtQQApjWv5y+DQamMddYvbNew0vAl
iIR1uPm8KsBn3VyNkDBWL13IxnksrkhyzG7n9OVXP7pQOu/ENMVSiAB0TR3DxwwpOEpWjQy513li
3TCZSEzyL3Y2285avrlziMatkvjmv9+2lZmpdEdAO5uJ2UVR6fxMD/7nSpgCrvCZ8GI9gChmI2u0
XYjrPhAibUxUNqir5h18GEPhM/FP4UgmXElGw2Wyg2S6aJ/HgfJOejCKQaFFJMpe4FLSRkx4lRY6
0UDMo4zp7tuSaSBUqwszB8xUOqY5WdK5h1vE92VTmGAldc/RnzrBXLL5CJrqSQwiWk2KXjVKcMpX
vvPyFLOKoOV7O4eftw0PY3fC/0xvBIqf6PqYVpfYZixG5+j3F5NEN62VZ1LKpsFajLJ1wKPjqs9u
HtxWcS1sbvUySOpW2c45yZwtMDfrdpPq31ZRkk2uCmENRlMh5ZMu8pSQVFxUa1x6Upe8AlUUIcCq
kj5BY3XjXyKmCks1lCtoycIVWp2wXt8XfftaMIkegc9rZC8k3Ki7OUvTOMUQEawR+ws9BqDtHUKJ
0T1TvS+CTYYqZTW7z7v+2v/hvOAaSPRCINi1P3P1bDhjUxe8gG+Zt9BtdIYGbmRe71OATGZY9B2a
40Z56Y5svv8fzuv8kA8H2KvMoa/fnq1E88KcmEM+Cwi6FxOx1QrtLnwbrXJoUQnFlikTUf4BedRg
F+IretMrCAMkrPsRPvqErl6EbKh6qhQ0hWNiNl7qETJ8R8sDjg4oE39a+QfzcmThI2nsZ6zMOorm
R6PVVJEVDwYibIoZA+Dw9eSbUCwzljvAPqFO1NCsEkcj1iex+KgCO3xfczBSWeKPD2z9GNLHpxkQ
pe9idttZ+JZ7iz3IHEv3kwGHvPWek8990HM67cUWDmC9SYaPdY6RC2bfgOnNcGLuJcyggtE+7Vcz
q6TSOhSHXFQ3/FjN5T6S7p09QPEwiTn1V3rru8ZEpo/b7vX3drigXE7BQeMSgGqvPoPcaiVx0Do1
ms4laLfQruA54bLkf5ldewJ87RFVx8eIJvuIehjnaBn4CCODqrNhBPvR9m69wJ2lRPH0obn8xGQS
yRffujh2CCQ5bsqDVgjICroc4OpqXpamfwG3lxwdLk2ohMa+8M9aJ/NsDJZTaSl/OxGGpMHZEsqD
52dZa4yzD8s8oTbvFyuh514SEdPAAiHc11Zmy0CkK4TJ2NSzj8ucvotsGMX/hE6za2z7vVwBglSH
dfKpLvQy0i5CFVckaMxqUyX8Ub4TkUUlyj81pkfxa+ZarLbm0ANccFM9KIu85dh3A/hlIuom9J4G
EOTPHi3haqvGooXsltmjWREDPXxKPPOlJxcfn2Bd8MDKahMginguP2H9VBqD3/RHhsR42XysADlN
mwj11B7BHKRyihGWiR7KvDjla497yFLJ9fonC9Jon34KHfpTI1Weqm0NtUBK/HswuetNl0p3JV6T
OdXh2zL9OLOcX1F+2JzXA+uxRvuhKue5wla+n8N8Wzk4OIwfW4voCr6w8j59FApgT5reeavqTOyX
0zQPYyvZKBh7aML3wsJYrxI9oIVuk1VqGzdVxe1zHJNT4yYtI7LXgedMZIhhCvI+dJv2TagCk/g1
v3K41XeC1oeK4wR4Jvkta+imdbxeuCCwimFxhTnk9boBlD2qTrpZl2CwKu28fVxLrwwrKxxd52RA
SOsYFMdLb6m/ZdhfQtsyzJxTI9k10nAJu+IgKNNLjYbwDp2vBQ3kupA5ZAqpJSwO/Y0HZEUe48Lg
u5obkohk1kEMzfQ7WxcmhhwXf/xB89sh9ONZ3wQJ8JAYhasIgRySa10ZKTeNsMMwsd5vQ/YikziF
deSOrwL5l3CciaAgJSarruq6i9x+YC923wk+PwoK7xNIqzHmbBFferkxAg36b8Hr+h3eCXy4nAcm
tebsQIoz9HRO1AS35nwAw9xAqZSkBBoOA8hIEQcWNersYquTCKw03AOr0Nfw6UIKkA/RSZc+GWHa
sC4TVea9Xt7+ca9bJeNPSfH6QmJoGPZA6VPFsT5ziN9IzxuofUrXQG/y6t3w4baCeqcrbtwFNeF4
7bmRC5PpHzMQi6/uQ9K+wU6E11TiwhCoun/LZvcb+ymIKIbCaT9FYugWfAV+Wbcg5xQ97+UVjObk
5kFBjNnVbm+18BXURz/79vpWTuh+v+KzFB+2STXPiYf+4nNA0nDvlpCYJoRH9xsmaxY2+HX5rAFr
YNt8uINkf2So0Wl/y55p3rLdhayLcTjRYwa41VVOQDKQdAiw14dKNk2iUpaPLuVzbGNcgtZE0o6p
aXvp/VOW3nZ0fl5XFZRKPBAAVC19dLnqpYdf7lEOuI8EM9n56xWnxn6Cpw9uejsNXrcHUq13JTJZ
yk9MoO2LGKtXrhfPf/9gr5oschQGckRhsU3iol7nIkCDxxDGv4/OC3J2zTtn4DqnlHr4jyL3Nky1
gkvZJ6A4s2nV73VxsIn+Fok8x15nHBXQ1qzkrgoeIu3jbgz0MhRF01ngTK01YsfK19k2p1+yRyEZ
4/4W9r5edBxY6foqaRHkj53P0ia4p2HhPXLxNL5r3BuXvJTK1D0fSkfHenh4sGKTHFKzJGxblpif
Moop8mJrUxDgaDyhcV3SaqIunvlKihy2TfVZbiNDvSl4LXJO+7M4iVaMUXFllHS8hPCiB8CLlVhk
G/HrBluTw4Sn8edQdalJqCaiC1VMOjjhGQ+0W0QzyHwv+PY3nhdIZtWX5gmNnzxCxAAMOEo69fc9
4R6qJ+N7q7drTnj3aNU/JK2JRLTQ4pyBGv1g07fZeJ2N0aGfrdlhzzfdEN98Nw94Ltt7acjpdhNj
PNv+rd9dPXX2Jxqbzxe3A9C1aGnlQBTXKlmXedoyYG4S5p2ZVt+NIscnuxy4pImGH0vJCJHbGeGX
Gd5PMxmzpYV4gy/5r3RLm2+9RPcQ/1lVNA2Nf6Kply08xLcCJ8RWdsPtQHgh26m3+xipC6QDbTd9
xzpFPmhXMGbsTUY3ZvMIKYOnroOvjy/2tpd9NikJOk0jK/CSKXNXePs9IUHJ9dR/961MCj292ViU
unatLuono0VDN2iW2n3rS/nNdmS5H4XVbUFRK9Fi6I0BgiQxyO5sAOMs1F/7g3RJsJWpKw0qsFhD
6U4AbrLbWJTGtU8R0C7Z4LLPpEb4aNn1uiQ61Y9XduoVgoV5vWGq8ivdk31z48esd6WsBpWqFdXi
s+aDSZeZdx4UEM/99hlaYXd1AX02m9tteZIjwudoKTpvdutXibSxALXs1xiw/oMQRxUFWHUcD4gm
LIY0vtQzkvLEzsZFChYQ5MSAENPQ4ihgDJcGWjPQrDb2Y3vZfLAvDeDu0viLpTXDKm0v84JpQbyv
j7do9sRKlPTEVdW8vTgbYLsQk5n92ljGu3yzZ9XBFT39y50VKnlUEhIgRGN7S+hv3bqbH+50Q0Rc
xK8jVc9Q+r63uRGhr/neO6qKreeKMi+7IHJQwJpxTHMHkT17TIWXzmLp2dz7L2ifiN+ehjSTmEI5
hwi+RXQU1SnNWVuw7lenHEMwEg6lxFqviwx/yBAlvpenQL0/K0MElGJGU8wM/IZILfh5iAA7TzmX
BwzLbUFPnmeL+ABYalfrEEEhLWOKyS6iY4i99433VSkRg6K1F5nam3U1xBDr5sRVm2MGcji/dqO2
KdsNqsAhGmSM8EB9GZ+tuMXcy9rG7c85g7qlPuWPTQ7o1fybLqZz7icVdTyebuQzi+SulOMbWm7C
rnom3/ZzhREQ+1I3aKZfBFFNd6Oi9tGELnWVepH8eLY3Cgsh18Pw4idAJHnKWqwz/bO3Lt8MkJCA
tzaWHKqMonBGGJHibeM0OMLhwnTRf+MZ7EMoCKuFj44dNZzPMvU3eRHTtfIIDMZWASPtLMP9ycLO
M83ueRIF6B5omQ4YbEqX3rFt/gp9fzcDUdwb0dElUmTDwGLSS98pxoy1grpy8wesfpMKRPa7m0Lj
o3NbVJR9T79gg48/EbUkX3M3CCKTWkGP7clEyNYWp2fBGXQinM58RoszPLCA+W2FlA/qeIcrAJRY
CyP0VaY3FPKyJMJdGNls1kLj0LjjUgt7zc0wbp41xytW4RE+GtGsS8E/2CE1lk1CUcS62T32tcvE
ulmwoWmOII8UXBFI+HkTy+8Jj8A0sYUPpS4tssWpqp0Bm2aU9Jef1836aTqvVC66aEkyJh6DyckH
UJigw/YKy2W26E2+fUhI7zzlMLSFK3aJ/CV6hAGPsj0ujYFA2DIf6snj5clO6Nk8ufdpAQvTR8H2
lwqmC7Dq+WckRkrkAPyaOO6h+52wutAPPkRaM19huaBr4DeZwDbb8mxJT2KOJSNxXhzz/hPZE5g8
+8f8UKiK7F/5AqVDfpVUlZcvvZeRNOk8/bzmO/lONBMkHgWVKzBgz0bZeMxC1WgQPn0wqug1XrOB
Bj4RmhuJZAi19zo11WoeWh0UzyQaFRK3GxWVCdDBlySeHHV42rAytmm9qM5Th8Vy9d/J1Xom91qf
FuI40VM4LdkhobYIzrGGxPCUeSkJU1jPQ8dAiOK88cF9yIjgkFkxzc6/mmsb2lSBQoxqTV7X8mZJ
/d1tzkWHtLx6uZj4mQJHZONCpPSrndf9QGSp/CrdKr+xwn1qBVP0/WB4vUqBkKQ4NoYEkXIBqFxs
detPVcs1x6W7W5+1VtkDQQYUPZLTa5o44GZwKFqWBPu4AdGKTq/ySfewCjYXWD4+G0QtL25G9jHT
UNXrql4m2qe0MZ0ebYxNwvcTH7KZ2QRdj7MuL6w8rKHQVEzu6dxEjFneutIw3ACI1YqAYnCq1FWx
v1vYN3bJLpR5biFftBIZ8OuvtwzXgCrU7tzU7pqBmxyoLgPVcbCrlpPebjuCUODzHAoM5YxXukLX
944IukVVQlDt6Cn1eRsivK5y08y1KK4uru5Q/Nfu0Rg61OfFsQVBlsIFcCd+tWUSWy+RlZP8O15W
Mg8c0URKvcVK7/dC09Iy5K35uNZZAPsg4tK9GpoDih+VOVd3vXvh5cEjtWVRGBg5O/PFvbRSUhvR
zZdx3Sejzh/rGMCAzx+mBKNf/6jWD4CZgTC52o0NW6K/OECtA2Kk7cQdIKHf0o0ZCuNF8wb2ZJ+i
eNJizn6jNxZM2/+vcPhmmqwut5ndWg6z+ksnch6ruEw/ydv925VZr89Oh7wo9JAxMnGj6A5b0Km/
ZJxSxvZ/dwxgFVxYlnZELRCYa0E/byC1sUrbleHoi4kNLP1DzjPGM71O7xySFKVz7o4RO77eQGHA
+QczSriNfeNNYEd71Ud1G4nnPFf7B85ohdf7rbpJy+/w2D1HEI5p4XxeHi80SmGny6ec8QzJ/m9v
d6TuO+eDeaQWXS7kTNDzrpvGLVMTDG//rrmZl3+YPMcJwllGDJIr9DxfmAhqdriozQOU+GgzDIcY
zr2rDiw30tTvjQslxturmBNyTbaCirzrZvhgKl1Og8J8+NWmH+JnBRzF9yB36tJgiIEY1NGYBmO8
R1rH8dH1C8ZB9Rsza3BLe2gcgUJyhnpHh7W0SyALncPnDtGkvdVmazpGDcv1jfS01TFWh9ifBTE/
5mbDe+EcX+tBUROBZRVdB1Rgwr2lj8lMMRvzrnrUKOEat4BM81wZJFzDZuAsengy/Gi1trSLCSuW
47PwQ1mC5+PISmDBIvRXZex18lk0huzxYQjUtgKiDW5hifxIsDZ9ElwTQzF/3J3LEnNmYJ9VjKq2
r6+AG8gAw0dzUhhN6mjhu8Brww5mmK4Y+RwIlMhQIr8mLrWoWgdTXdZdkNfwisRDQZV0+rIuiRrd
n8C2Be6uBR8pPjc2XnUn+TfL0f5v1m7fPbeqEIqJNjTlQM9uONS7ouxqiGKMJsB3PqHt1vT/Iqgf
+kMJ80UFSw9IoUrpuZzKEnZO1n/CSRY3UFrKAYllqMfxiX6NoO6hqvGcDSaqstNykE1U6ZUMrnQk
g6l2RC0VqlGWpSvK6xt5eh7UW+Oh1ZqZ0HNSWrrFK1gEhNAgu99UQ8rO5dBy5lYeNYdBiQ9W19lc
rOspymZu+5z8ik0o7t37m/ZVhqVniQyMcPWiDTwYc+cwh6qiXqkumtPNyP6z5MyJYfbysAIJWVxt
dYT3RyEDqC/urKbfpvuzFYIhVeJWF/QYL7Y9Zzbq86oWoPfSFqznpSNClK13I4WbU22QbTHOH+ou
GdMbGwmsKnv3bODW3BrHyT6TPzwLgJlOaLeF8p2yUSGP0AoPSak+JrjflKTL1/gt7z2YRa7SlkOE
O1pBPNWgUPxh2e6tw91D1Hz8zlH5TGSs+vNs5vKKN33IQBwm7nJ/M+fW+4i6BrWx3sjH55Mzu/Lz
QsxhV4uzV+wsFdkoV/5W+ZfI7LWL7fQu8Uo8yB/ckIQyyj0tJrIidx6VG65MUQTIxVWAU63exJj8
OFqYatdgE98MmlegSQXitZ873gMPC7ZyfPFt+5Oaw5bHXIr2xGYEkd6KXUWn7ZSt2RwZJnDlrP2+
cymIV7SQcS08zJLjMkQ0J3uGWGj5EPGTXcShcyJmhYp7refdsQ6KtJ3gc1fu0urOsW6OhhtpeSxA
8XE6XlKvKqZab0GdJSFVxnOYhd7wy4kMOZUzrXBqUA7NIKwKxiNHWzsaOdT8Yx8tsjx0UzAva8tV
/BnchRh8lKF3jgOslWlO5oIRJeQQgsnR6jwlXWAYFhSqgFf+gi1mXDWUV0REe/yVCj/H2+qv9klt
UysFW/n1R9Bs4aClGEx1019m8nSs5m0DvVv+SngUqyMj6td9k6UX+n/mLqAa/DgVMJpw6bagKWJt
R9/w85M7aZGVg26O8NL8l6rlu+9VOOVRlo8y3F9Q6u8tGZj2S16xYYcnLurpnme65JLviPWx3skk
aleEwioe3P+P42LMt58MHtvH0cGT4CbXfEeGsDet5Nb2xPKSddJzDNSiSg4S4D+NJiP1gXw1uFwJ
WU1qH1GrhqQ52/OcTcoWRMKxT/Wzi1jW5+liu77RqL6+t4cHigAbaP/oDS9bxseCalExt0X5wvPB
FmVWN6NO4Mslr9DCTLndYN1XqGinobve2RZCChwvN5lE5bs/TdeIOSzOemu1VT1wgyllpIERLY98
85RtxqSNvrZv8+qRJnQmb/y1oGcw19jTA9uaZdW+m83iZ9kAy+i1mLn0fghilA1UECKwazEGo4gq
61HbvDSUdbJuXs1zr6F6zNmDEQwX4Mwnb1xfW1byginIwwkxMtXNdocHtq8FPf0rMsRyOHIdD8KZ
hk+Jrt5JOZ6R91hNDRvkpE/RZvfV4OmgjoycgfdjFi+zArByYsXX3AVUgwu+/dPDZMdfFiSMWD0I
BfLiLPMYCO3FGJY7i8iYi7NC9oy4BU9wM5kXmAGcBPls4+pZFnb84UoLZmvLb3etzLWbA5dzE1Ap
vSw1GxPYkJi7KS7IooDT0dAB/CEGDdWTEF4dP9pfUVwTimfOChT6d1inu2tElIKfOzcL2EonKaY4
P9DZfP/xSHf2WN1Ah5pmfCIr6MrZdjQ5znl8JrjzI9l2htNUH/IIsaBTomb8ie3ZBwcQ5tL826Dj
rHsfe82Kn8IUC0GskJYVtKMZ/SiRAbdP7JjotXvSjOpBzixmQGo5iC0HemrMwsSBokqbYknkBKoQ
Ss9RRsR11O+MtO/luA5h10Wp2biOG82rNRWUyLs+af48y/XtmODr4YWPcpiLd2qtJ9Ts9Gv0RtYs
oAFf6qWEDj3lO3Ji+2ccnAAkt9l/PRf5T0CRywF/qMFc+B6eSSt5qG4h5WEQDXlR5SJTZzMYoQgB
mVTNEWx8AY624/uSdEC9LlL5szVeD0gb6YZT7Nnhg1bfyy7hFa84DqwA061c2E63WQ1iPpQOLorB
2tX4F29k14t13w984ICAhkTiu3alIabHUz4CTYayOvKc41vdqvFozaR9GBzaTPRFIuLkDe9AcR+v
AnW4c+uQXmbHoBPPzHoRzBQ5ik0Imx0FVfGSg5e9hmZUJ9SyfTgZKKbqUsggyKdTFBRa9POPpM4a
g4+8X+YgdRvmvc3WkcYHGlrIyPBE//HntL9UTMuiCKlK4JW0WPpIELCiNZVVzEqD/B0mMKOEvN4q
2R3YT2unbYOkK36evGY9U8mugmSJ/+xXyQEaC9ozyXtZVgPIugf3Qqi+lh8kWbxMQ6nueMLTXYgN
JBpU1lYckSp1lrehjjZ8sPcE7DR4PlpD7gPRfR6TENw1BxmWOVn9udDZggCVNLxKzensrLrFbRMA
9PYXzN2R8dJi/vRQY90XaINKdxMN4NXNJj7CoZAOL9JAD5lwpRv0xZU26L19/TBMn400UdRUlKB6
4fB10Ns/jbVi37x6nWvpv1CfJrfryenBd+3MRljYg4KpxPwCTSJ0Q3rftUlc2eOOVIeQicFn/mNC
XyHLevfYOublXJiQFgj4yNbtjy2HgTWTtoej7IYf2JmOT4fHNBdZqVsoNjvXk3eE7SblZ4TSbuzD
WFI31GtS1HLiiHyI+7y8ROWhr+EfGfpav7IRLulpfTcRkfkkOx3pUpwJT0zpYOgVTgPtJkQ/8HEu
jX6kw2aJJ+6gYnL+5f7G+BoDWySx16oZ7yeoeAyRcPsxu+/nubPR2qK6gFjtlOkXDQLBk4lvJcI2
wiznLBCqf3qhV/v6LQYlMqE8JFlTDMsncsJONUiJ11WAJ50rUVhUjk4Rw7oB9cndXm7GQ8+maeZM
F8zBY8pXLwV4qgJl+OxAkumN1MFH+XB5F+Wi288rZ5bxtacr3aYbm1QVLiTI52iAUFb46/fgUguI
zDw8NblKc/af2IpEdW3h1dxThc/JnhWvniArmwTqH5HJ0mQufyWHvV7yvDX0nYjHlaRXyYvlfuQ1
JO0Ul2rqFsjR8cqdx7ln7+Am4vwKZTaEDdpbhqqP+c9pR+q2N3bm4GTXffQTmwGobO5IMJfIfvPL
zLatK7nkH+/DX63UO3qbP3/tYoRg4eM4aot3Do0oIRC5/LzsFjUw8tlISH7sQj1HO7jL1c9zzblp
wx38/JFtXSJXYF1SKubMILiO0kjHHatcwe/+Z9eq46o3gCau0+v2hmHiEWXMReJy48x/UJJba0O3
muzXN/yhFuXjbuBCvS2GqkJmHXXpLM/b//I5Kze7QDEKpoF466pUejawYqaAMZ/LhhGJPmPYEwX2
athbRrZwmwF3ijuegrwch1/ORu/k4JSA7Q87+/vYSDslp4/NE+OZ7ESxuLFFpnlXemQZEJixUye0
8tF4yGCgbQJ733pqQyGvrDYDZGZBOOnrTKM9y4d4vqn6smx+KVseeJ7bKEYrZ9sVYztkOztcxnok
uO2MV/kHw9uviVKuv9+wJkfjryCdP3IcWjwpyNL8Ukr22B9rLZY/2ZQ97+6uhd8Oxi8l5DjAGHZt
hfPa4CwLTsnQkj6aNTOMG0eC4NmhjpsuEDc+mopQLcFr61NZfMYVOsRIUl8cJEtmeNfdmAICqAA5
Cl4nze21nOAKGkWazpUanb0uXwL0aJH2ZeqPWhzhCPp3qpe8WLGOZJUOvbDIj+oGV71AcU9Ur8+Y
qHW7rNw8I3faWVAM/EBrMiM6N2sPzgx5+YdyjvDskEmuXiYGQ7qwnloTMVtkqDw1u5RMLQeR2Oyt
ASlFEhOqmN3Yh85VjafPHr6wu0ks9aIsUCUsitJ0D0oSDSA7+VjPKzi1PVkZSFBeou+zzoeAkBio
kcXFw3TEl1AaUNc2najEsH+sccHgEg0JXs9UkHO7KwVwWxKR0RhfNaBZZkKXfg5jGfbFBr3pDfDt
XAOwvhYAN3JEM18gsophe7nVr1BmAB0+fxPR9qlqTWFC2nB956dv00nqk4ZXsKKQRYBoQ85hagPu
9It41/wLn01ay4wilxR43IWot+zUxL1HzgxEtPDs23gCl5/nzP9q2JM2Gr3/0TOvSmBDMcNyIPox
YDd2kqCb4bQ8Ard6VauVN3T/t90jYSw21+DITP6nsJygfgpOc+OVOGR04hTmyh9nF3CpOuJAR9jb
BxNIeAogA2NMPShEx+7Rx6qAT4yFvZo2fXy1+IM2Jr0fWl9Pf/6rESLfI7VKJii2nWqOe0t/t51z
y+F0ipBVhamRmegBYxWFyxGHzapi2Tly53+J9qm4qoygiOWYSybzuO2wVha0H2cWakGLaC1TEToX
RA68uZYfkXCQz+oESgEV1Jqn8VuMMBBCuyiGkOOrbE89i64jqzJiUID6l+5rIj+JjMgPJdjooriF
QC4Kd5c+KDy210Qe6JRv1nEwfJLxfYS62+NsFL1aRxQ5iuad/fxGgyAgkqot1mjBUQNpWUE4BSFz
9755QC6XN5zQdt1KNCgjQeyOxSgGhKVbCUdeLSpzciiWr9f7RVS7BKqsSe9CTtXNwNgmQF0POo2C
HumlEBmaUUBrnsj/gVIlzkRPv3xYTysoMEH7LBhAzQ36Ix30Wf5XOHvLaX0uymLLQYhyH4b8zyOj
A/LrMs2UNlfcwb5C/J5JlFqw37EqsMTwQ+RLlkZbW4rS8SEPGGttfFxz106Z+9XxNQ5YAVgE5DAp
ViB1mgvwHTJ2cejEK7VHVOOrAJr6FHJ6CHAeXm1Ni4FQbtTq0AfDN86SB+nTPL7wjsftzeFO593I
Vlo8UpuQuJzBP7suDgfpUI1BcNPBlNb8f0gF4NX84BfYxbzpjLqIergPilz+cbPzlvMpZkWdP0UW
F7ASDIP/t+H5vxAqEhDjTY85oUlvY/pdFlbNk50W1HXdwGzhTDzo+9//PtJTEEtnrJ0br/YN05Fe
B9UJ9Bmf8ubKGo/oIWGenHJcRvLgscBjcNZfoBegAXzG1jYdixK9jivZlUSUphiGQx4c4Y/9/23I
YZqYsDqTVG7iDK0L3okZj/oS+ENp1pH4YH77YQiZj3FInkOA81xyrty7DGoqdOEOjKKbyJlmNRyX
yE2OhbK5mPD2RWQBAljtbYexuqijymC5x+ngnz1VOobJTr3lssrhltXnyrZ97QJs3Z1uUw1JvCUM
n295SKvc/T86dKFJmaPu2xXr3kJE635H5dXKmV4ic95ByvUB2r9LeUQK8pQWrUvYTBolKlmxtBAY
P3tBIduzxRHy2Lfzn8ItcHW8yunu1t0sGhp4gsf6DOuEsnA44nMn0xdCegyvMDtQcAGBD1FjJaEN
7nz/H/hmri01Qa2ru+OkpvoKgrFGzS5L6xRAtaZHdKyZGDELb8kPyyFu47hrpqb8MNcarJ3IUc3C
2if7399wTAfA5PMPlPjUMdKeg5GlG3WC/uaiD1tH8spkvxOt8zoetfNWbvK1avl1oz1QkYczHXiH
LLAF/vkKJBQkQ/PfoYYsYJ3CFWY1Vtd5EJ3TMC/qkRnj29QPtDVi7VGuv4ZAmoctBeA98ll+xjbm
p8TDmnbV6SABGCZ0D75JO/8Nk9kygB+YSkkOJMwMEY6Z0/Zw8jUNJZ/wyAfOHNDcQHcL9zP7w6YV
ALNH4CFXPDSv6gvVV/seZyCWkH06Y7MqRK172t9epiMVXBuq95ei0MiCK+tTtOzjU5BTYyjiOLLq
A7iAmwhkcscUe+MP5eAajlk5tzPGN6P8tgTEeA2brMZo5WBovFzngvokbT4KesBuI8AFOAgGabmQ
S1rxvaVqaX0ZsI9pFYVq1WOCGfFXAFnKWU1G27tRxVNbWZMHKcx9JUvaByNwWw8k+hS7wPKkFy9T
+PWsQIFNGLuWaqxqlqQUgSBUWbtNSGm0z44kt+2QwayFRAiAhC6DdBurqcJFk5prMTpeaSCGAITE
7ILqTzN1tmHn+2198PYZlLS14KFtTcVRBHnI7jgmePLZfZQXgCVuSmIUuxn53Ect03TscvUAs5c3
yEMO6jtrldGmciwQNYoNbosYDh3dQ1EfOfXwMgpcLOL6o87VLemL8KTh+GiYnA8EJDSEnxS1wORS
shd5mYMf8sggh6IO9Vlo8Nvx6JNheW42RmVSigan+AdptCE5OQqAY6IDQzcS8ys6hECmCkHGzgua
YOgeEEm5SIrJWtKbci4gJ1dT956TZFKaykSv52oNRkOc/zIfZzjAu9WQ0/qkG7aiZ8wPUkDt1ouk
ElfImGqs7jRc5BgGo7GRLoiQA1arsZeKeJ7zJsrBYuRwCuBcBJaAlm3Rgk2EePF6QwmhnwkrDV/V
Lec5rjIZyVwdEvXVfd9hBG79KWQ4KpkQEDBehPA0cB/Qqq1w74dr21fwUWd5ux4fIUQ+BmgBkxB7
hN9erHstj3y0b5LqKljRuB3ULKQKisZC+vVMu0RyiroDQdJMjkstxLd4Rc644Uh0+H9Ma0lU3U2l
Tmsu4muaBSTPUFDn14UZ2Wuc8+wobef3vsFrzRck1K71MNKg1D0LFZBlwfWwBDh8/IlX5p01UjkF
JLugjp2z2paAuC4KK8uDVx5LpXbOcdzUdT8g7SQib9yYLzMzMRFnBi/5Wh+zkxIQ209FKh48yK7T
GkKxb80pQ8Zi5tT3QmqoTcX49f7qdfd5YiAFV/+CfqDcyVzeCRcjldVQVmwZYRTFTv8wIhzJ48Mi
VQwXl3nvouDXVHShDlcZv7rbYUZmenoyQ8vm3FFEmbwKj6NRgbF4yrP+17wLK1ljIQhZpy7jrsl9
u5anH1Y+pp+WQMVDyPnFO7AZynhliDKI4OhpJabU1weept2bWivTPmXYhdR8r5s2FD/lLlF2kBUR
te2CDqCQnSspo2lPCZxCVtvPyupANnnWFeSlhe177Gf4yckrXEwl7K/9Z6aF6esQkLGONSNAKpSE
1kXXhxr6wRPekX8OKo5JY5nU4Ng2Ye9YEacvFhIGSNVjt1ZeEmPdTYdylPSCwkSu4Ko5Hv9nWSAs
OL+RfDDtcYB57atlD8HFXbdYl1fINUOKirvcxERresAA6WrHW9GhNOWpXvck2c00VT1RNtQjGToR
52ZGA7f9CJ7UFNVMAMHdhxiS5zXs+TJvhzTl3gP9TBY4pQZvW5uYJ4/riHXjCOYZ2G8cO/B8BJou
HLpfNCBdVYFMYd7FbiktZIWHSWUX//SVKDVt9eafdx6xlSa8CMrFgC9g2qDFxj/jYlcrZlGM1gaz
pYSEtqyZ0H1qVCLz/edOPnhVkNu9s8PDXax2DztG5lcR44DmUtzGjjlliy04GJzhr4D/eukyVjxm
NVAo5cVZXniwS+58aZSx2eZW45XhyKRWaJrmDP7yofcZ85FiFXnTN7/Z8SJj/CBone2pTkHSBdOq
VndebJ+A6bWLDFJsivKmklGPwlCCLS05NWA0tc2rVgjQFNKkhHF5T738+ttpOQEOAvX+/7qV+Tx/
DlTNmy8LxJhhQ6z6dNytHmoeSAiTXOcUhD9Mza3A8rskvNdfXTaXWh329h1hklxC+M1C0GsAf8ep
RBdOttHA8qsFvUDBDbiYkuDS7qMnUoY4gxGvoqcKbv6SUQsQcwmsc0shIpZhZQxf8TazDs0d4aof
ML8Cup2Yxwue+I5Icf/vBIjUixdf0tIwv5t/XQyWG+s6tLV90XLZ5w5DknUrQNVqp0Di+VHL2yLx
cIf49/eYrGtN6zo3ra/gHiMFCBB0XalAcGWJCJMrMs6tCUg9oYsxit4mGgyDKiPFR4AEiaZV4m69
dXFO11t94kN/P+PYkT5KkKde9BHQZ3dXrhEcNRjuXN9mH9j2cSY7D+ybSMkqGhRtGEACvffFnUNx
WgCgdxEERdMe503/wqdG1ndal3RMvjLrq2lKa8ELtdjut6+M6UVOKkKyHMg7vYjmFy6iFx5CMewN
HY62f9okymjs/RgfHZqDdedjBlsV5ivhwb7mgeJGWjLbTYIUJa6djUexzy2x4rDoHjkr20DKiPAw
ram21AnXS4tKDttntkW83AruU0+H7i3kNr0NSQucB2ajKmm6O8UOz3cLjxwgKa51o3LJoeO6lrig
3/qfJu3/KGWOzJFmqtE++bnZnZfrMQ/grFxaZPT7mupwyfO8FQfN8bmL5qCUrBO3jpGGazQq8bX7
9RbTu+FvzJANVGedVsn2K9i3GCxUfWNxqHfL3x8y03xR8E/c3J1flTYheVdfdE42PL6VebCV5fVT
WGaMxfUE0RZrI+rW+NJdr+9xpWTm3oRMpInIVur7Te3pUYOtOTY5L/XGwFdo7ircMah+XY5iIMr+
+nxVKC0RuKgR2EPv7Wl5c1j1zg4+0EXUViFcLaChyLdy4U0/UY9uXo4vRkMNNay+cTJQP5PFWluC
mthsTK3fhQXyNUVPbV7iWrgbClr69Dhx3xTjT/C39vVkaQ4fZKlz+vR4Kzn/QzxvgoTrc07Sx6y0
djEpSDos4ueGR3/E7Jd4jv7iXMDuOjoS4Y4SBnT0+3Bm6AITWleia4ctJIePvb/xTO2b0JUooMhK
sgxeYH/TvgOOFly1N2T73RKYaFVfvay1o2mj6HUfih8c0AbBdtpvPS6au2xtZo4rk+sLULsnFXFi
CCgamNHVAw0fJQeKK/45C/eaXkX9FyFRyCZHYr0B9FSDSoAEUQu7nE8wmAa1ZbD4RnvEn+bwu0Eq
ABLSO5acXaxO8xrpavMWpEIFtqnZZUOUp2vzvthKjbIPayco1uAL4CHHT+SnWx9N9f5ZHuODc1L7
xiSt96oZ2ty3Ndbalug66y49uFkPk9N4n0H5g6Gemtl9cVx2tr0aMh/fDKxrE0Kj4S27Vf9haWxE
Vos7aevqqYg78MZLHk7qUD7E8qPVDVJxOkF6W6nnDdKNrgmeqIdLk22cBWXlAirRB26R4b5YvUcw
zfwcmAKOg96THrZqIZpRlKI5ipcKl0ABig2xtaAAGNG8PTWodzhZ0N2uUDpzP4cSbUCe2l2xr7qa
aM9nZJqz8aQd6gsLl8biSxfsKvUSVh8q55y0qAnt61Gjr8ndjRARl+dZ8UncoIlmDq5CvbudSm3Z
oSk2e75KvgIS1oko9TSecaGaJT0nJSLPvGE87mF9uU4p4Xp6XqPT5x4ZSYwummSgXQDlILKL7cd2
slyWZSUFRvcdOoCDJ6+XVQfhTorc+2lvux5qtR1ewx5aiFZGopwGNf9N1xXwN98N/AegWHwkN0uI
lNjz1loa9v2Ge2tKZArvZZMtDN40r2ZK8KtI/sxszHAxZ7z0DMNfz/YHZSa5Hgxi/TppilMIi7+M
S9t+hgqkL0C1VCNXNqG1ZCA3RIgglaXmHobgNawebucI16m5SsaNhRC15luzyeMDZURl7Fu42ZTj
EdiSDQ8PWiY9NXOsLjeRN/dJEEWjRnFBvBrwYzJGX9us03TtnNCi7RW/Z+TjOT6ywqf4QQmkxwBz
1GOtf8rS2f1Us1OsXMn2ENLUmwJb2+W+EXJjHeReBrz++kuE/GQpylm1eAD7dUALxgecSKeI0atv
nKpXUv5+994EHWk5cQ5z6zddqKsqinBDvGangJCHe4b+LDByl5l5vH6qf7NOBXG3WsI31ffA6ybN
vqKt2EUXrigA8OvuORTzc1w2HItPQmB+sqxaUlAA/keI0PAxc8Xu7ztvtJyJT4XLCQICOYjRwJ1l
6u3nw91jTGUe10oximCDP+kUn+rjqll5Tm2ajjdV4NN564f/H+CQPQf+wVgkSgA2WjC1wVU1R6Xy
59OQlMgeGFw2k+unC/2NNbRqEQCCpkOEiPBFh5/Wu1WcoFDjqnKZNZflWAoLVV+RYZ2vQ8jP3abs
cj/v/se5IHgerfuYU5+o6Pxwgw1gws8syZBNRVExBIUVanu4USP52HDWhhYCbXS/EEb9igAvRNEY
LV99OebkI4/4/4FBk6qvDlrfGzbyDZJHVqDO5vt4cVV61V0e5x7OT2XodUc18yY99r/uhT8Rq+Cx
5afbhQqzvcDtI/PYUME7nZTLAEj3p9Elllmo/6v6PWH+LEtMfj1Ibk7NxT67SBV/Mr0xZZQeSA6N
t4Nvoo8E9/VOE4CU5KubOOY5Dns+CplYw4wSGYPaJv+qPweL0hxzpqt1thEK/FmJvrjf94OEvVTL
owdFs/sweHZo8kDgUzw3P26JOXcGJyO8R3qFZuo/CbKgIjKZMJSKumSGQW9IbydqtM5/ozqTbE85
yqJfM3DoyCM0ZMAKCKQSccNnWKApG8OD3tXqzy3bpxLRmsaNS7tMNxZDGM0m5d1USBzGXb/Lyg6f
ygJtHScW8jNzyG0hCDo6B9xyf4IgjGqCVpVDAAax8aM3AxVCSJfXOplZin13H4lkz560iZBGOWmL
xN0+krTbHqmz88/Ckl9kKyPaqOQqe0L4e2SXxSx/sulxxz3xLRkHOfCqgxpDg+QOZByXeLx+t1mi
ubsYTtuZ9LCzTXKcWkhhQVI4PhYyo12uwk5jI9kXogUgXxvqLFOZk4rutiFdDudQmxG/Xzg+scGi
ZuJJh1MEN5znQip86FSmHYfS66/tMWMomFTNU56UIZ5LUYb6o5lFnAybmp/2J2D/qrhwkf8Duo2R
aIu5tca5WcJVoCocYm9ATH/SEBwlhfImMCTJDEMnOS8Xk7h8dIE9MmyVBZgBuWfUjAYSTRJs1w3M
ieXn7oDASoom4LG262W4PH1C03HCQICLsBoBXc4deJ6LH1BG6bW6pkvB2gnc8VQ/03p6UrqpM156
REwjb5u7XMF1D36oEqqJ4J8adLHHI74ku9eRsjeqcbjU0VzpogS+OOBGhhkikZdBRFyrDqlvZMAP
mf5C4tQ/yc8q5QgH3NK41dcizcQ7sbYhBUvLpVwhHFnUFC1AnXbZ7CpSb9nQduIQRn9FnqDHqUmA
QidLFzQ+oepnsy38ogrZRkoTHbqy0U/hdc1saPQ0v1BRCfP6/7i8f0INRjXy4r/9n80UKsuHP9/Z
VLAhD1Fg+LaX2JLTqH1JuluZE1nht9OMU4NEnZMKtkGDNZ0vBR6IQsgb4dgF9sTj6ypYB1C/TOq1
99Ezew71dtZ8E8xKB9DX2MzFsIm0V7eSGbM27DC7UxW9K2q9rkICX+uscN794g5/mlO5zKzWDQEp
V/dlK0qcXuRA4aIUWgbmp4lgVGRgnjgi2oyB5BDL3ttB96I6XIiWvQcU8SdsdrGqjRAgczgLc1Ey
KAlRAzF0DD+CVVoGd4gdLWqzlpdUZU/maoMHDuQEE2KNx6rreQYc/fnwTBH4gret/FtZpnCxO6ps
50TssFgJd66yyUI0TJkrqkmgzaxP0/yfrm4KStNUy10XhivyjrcKUQMhE9SgPPKe6x8ct/NF2zg/
96zELibZLkddcuILdSpmUnpToi/q7mOOGrPkWeHFr+/qvC4VHNzBVkd/6j3dm0GjOi634H4OfASy
BYIGhlS4xtqZ7bwYbr6xVKVxWP6JD4kfe2UCwPAfgp0k9e8pUxjyXR25N7yASHUlD9J09B8W3cBh
OAJKhf6T1WW5sbHaiQQ8dbHk5Tem0F80/OoRRI7/9aSD/RLMb8aPBZKkxVhvOultwUfaQCGapkAW
YoaoO3/Tic9TWh+UYp1ndXbpEvEy7vZO9R6rGgMrg8rmroFiqnLIB35Ow5xeEU9SxSqE4h99fsA7
xLkEIrsVbR6+weK4Zwr7gc63x/HiXW4SkkEJhhXwGAG/fwh80NaR/s1c75UiAQEZc53bUy+j5/LU
PtALbJaW6WsMtn/4vL+lYzCEZ5QCqteVTx937MVPVipcr7JDevQyyb1j8DHc5tmYTAHpfdeqpiKq
yFYSunjQqrs2lQz1RfcoX6t3aVUlXS8+i8GUHY8r44uMh1nneERY7nuLNkbDfzxShRZwjjZ3t1oy
4BRQakUsSYqOhdkz1C9QyW0dJdo4DUVvBJuq8OnqUGIZQZK6pRaVG124zz5rSRze3h8VQVcFR4BH
sNS+ZsF7jgXRVjO5P7OzbY21HinkiDVh+u+IgPxWeL1eqEGTlLl1n1Xrq0Qk+nODP8s3ETEhXKH4
FZMOrW571SV6qjXb730MKYzAxkESXXMp7gyxtTKsk0lmaMw/3TxTBDUJyvAUOw4HwbQMUzemAZD+
paTqIPUFawRbuwE3xufeS3jg20PyzADsCx4+dHEHdOZGWfIqQzwr7w4qQSbJTymjedihhLB3p7zL
Zv5s4rZieHvwGOe6si97/nX7MA7LCutkhiauKb2gP2ahxAMg4VyGmnJMPo9Vxyzx3EtvO+qDjvex
0WQG+/090VGPLx/1Iv4Yhr6eh1TzY8K0KWWb/+Os3NOFAgC4YBAHC8NWspqsSkBSBWGbfFQcf0wn
sMoyIfHevVE+7WHXIclmZtmvkYRq4/001q6bZwYgXhny4Pf+74lqhDA0OoqCx60vQ5sL7GXlSn0p
hqWqt72NxdrFjCpqCgaWUKK7TNxx7hFlKcq/R6j9Al0Z8tW+Blba6lnERxgriAVhcS6jVtmh0vS4
xcQxElFr3LN38st1mJ59xCpbotQl/DgRZBtFo7AHpXFXNWuiaEvAvPWEIUL8/BT/ypL6dJg+R61j
dD1IW13DpobRFaOJtBQEtcyCWaif1ii+dO2fO6sFh+UbTa3Trsqu/lD0aKlGenujqgkcI4KRf8h5
Ky6zOEY5Rj4ikmxvRpVooUOyYWMoG8Wtg1cMyywbloDqxMpc+me58H6uPAb3NrcO9My2ykzqZPIg
O3fYtI/rXjMN1YlJjtCdnaHeMZaYFbW/tK1E/w0tZNnlQLer8uDQlyBsuvClyzzLE3FlqeVz+m3z
+uQpfO4oTLgc/LiIMpF0UNq4UGaWif6h9hT63zT+54VAaMlzIm+86LPZz1ez+DvGP8swaYZ815xj
g8lixi3MOBzvtcTeR8JZwjTDdd03+2NERK2TgnuUxNeqrdWhlVHJtCt9uEfDnMa0TCX70d8nneih
6oDVx6JOGkYhUrJLvK8dZlzbnf65WqQBoasHq7YKaehT5VNzu+vx14mJpS/p8haWfeQngC1SI8nr
LEhcbd58HjCgc10wDs63/FEQF5n2ud2hdiAcs8rK+stSO4MabTmCZam4vTgHd2sGWydD4a9Oiqj6
UMpft2C48OB0cJyJBw9MiNqZ+eYljuMVPKkswqHLcjOB/MdvrDP2ckdqPInzH9ntvSrzImAg4H0O
l1oAQKfUzVxwQKlFxCI/ktp0MSDl+uIYY4iF73wpniDlG4M9W0vmgnhHmoLG2V3WKXgJiAZakK6j
SgNGvKPU1pe7HiFJTnmp/x7gdGEhjR1LN1TUKHTNakJbvplQEfEzPmLR9cczp7rtGKxNGinIAGYQ
NcTbhnh2MHoDFdyeAEWKrQttGqgo9f7viuMOpTVFsC/2QhSV9UG9ttqAJpSDoyjtqOt8z/MXkthJ
fVAc5JQ8mkH9f3a5ocFzmfnddMViL/z51z6w9MJqlcopDAbFmSKQXAF1Rop8VSg88+T+Cyaclp9o
Am69YD1EMAlmZi5lbYpt1PZC0662l6zLGP8sHZ3/qtrh7IjJXbRuoiDkVML7xPoKmvywynQPa34D
CqoyAukIEus2AKARaJLnuZi4usBPtbTrK1JsUfJYLit27CO0IZuYvA4p1l78+dd54KkPff4s8tWu
eqeTeK1ObioH+sl25uY6+uPb2FLifpB5awQbwuY0AxBGLasMVGheyC465xZhBJJYtvZMWko1WLth
b7Zoq2oJsJCH4ikuqkhn74NUUF5XqQjlCjcDicmx+ZcvH1rIG23UWvcfaCQ+T6PW9WGV4BXTSYiz
xAc1Q/Ji15X9dthnuyo8cFBvllT7ozuQXh6z39koBR/oTWbZ92GlkS9EmBPlqRkzt8u9kJWhWupI
NDNbky0THfh9LOrpTmiGetYL3HQnuuJQ9jv6gpAneirA8s2ei0zWV3aHYdzMUJdJG0cBYnIr1M4o
QZ9WEW6oRLAHNLLALqA2dC5jEcArhu6HvjXWdHykejS8zX8J1au6DYE2o8IIwvaUjFwdhh95pP6r
uJ0EuMoVS0z+RwqKlGkUikdfYue00O3ll82xfor7DMfCojQCBxG0K2mVvFu4U2M4m/vUFer9NW90
gyCSMlSAttiFudGjnL1mc/rwar0TbWTL6dMN0tSEpANV5GVmy3hZGYZsLhKmqeQwH8ntxjHyj1nB
k5is+a7LJMaWqzSqBA3fuxsoE84TTkiz88XfYTkvRZ62GKrB8bXPx3xQF+9qdThtAATbAH1YPT6j
wbk9PqII8sRM+RWWhEAPnRcqRlTCJyFz1nxTVUdEY98ISCXowIgLTr7kunPNVLe+droCwMAe2Ut3
1qWXAVFyFGz0n1pzm6uA7u1xnf9LoIfDKRd/aTBHCbpOpFH8eWp9LgFYJD6Sp5phu4c0rPBn/aWV
fOHLVxh8AYkDJzw9o+F7wmYgIerpM+lNVNOcRVglx9x2kvrh6pMUOSBicZeP+/UOelV7cGegbCQe
fjVveh8gdGxRWiHIK+2y+xCXjSAd1pCZ33MA9Md/JuzgcQi60/4vIfkFAda/IsSwSFsExk1TP6G4
k03JNPFetybfgNs0lp5YtL1dmA7GZq++dpcvBGtw34ND86Sf6ssGyKLFpYmaZTIAE3hIv/XD/+uR
aOMcRFASEWy9Gq4L6gMnpF0F8ZFnvkOndQm7qf/eHHKKqzkTI/q7OvJi/Pv1wPD3G7IfEP7pYyKH
8NPLKaSQg3Q7vX/Swxd4mCgZDClZDbKtlj1LGjVqIfnf0tAfsCdsrnegsSIkcfZUV5p32uv5oglI
oxwT952HnuoFql3FtkMDVA9odM2LXG+JIV5PBS1ZFnFBJi9t/SiouVG7mIxjiGqZn76Z/zPUhkav
eoxG3TOpso51pBP/BiK9xFyZHKUof/PynqrYSCLo8Bm7mcNBIK8PQXujsTvgTZCl5DQGIX4G9QYo
+Rk4udHsGv2fPOt+RdLuyVKOIsMsUp9hkkrgOQsTTHiqOVuylag/noWy16Bkow3qnBNH2bpIzv2I
/FIFbZ9RhpHnv1TV1U1bX/gTSgIqxcV6BrHWhHoTUShWPgL4Sy86U9lnZn+nlGMdJTnth39TWw2p
lvk7lvag0pY9voi5cO4Ybs5b4tEsCU0YRxxGE80rHWaGzRaxJsZkqkd/Bc458w0VMqSu/92kEknH
0MewTctqwwQM6qcp6ASlavbmzCNwEjNn+HVSVu9KMFCxi7D6ECu+HVwpYscrGCDsEi6WkXq/2N3Y
mxrPJnfcVEOnBo55PNhBbEomj6THlMgNBXTVYRPfrnkbQbyr76Pr1Fdu3zU2kOjjAOtVbLInXW9n
Hmobg+y08gs7DpujiI03ZNDnAdoCqgfvYyjkVdOtY/fsiLlyCSbCoVJO5IwE6P9xlC0b9r5S3zMa
6se5HORERUTs4hfgjX2qeVxwQoxDnHTCpuvM+xwLKbZ5BXUiIE7Cmvzj2I3ezor7dF7yV8MVr1dt
g7OsPCzKUxLpeOcH5kDp4wl8s1sfllcMqhJM2Hq+Vi6kDbhehcaoDT/EJEdQCv0G7oX4zbQJF+O3
NFbCr4tVOCjIJmZXsZn+XjSlrkO+FXuOwr0SwlYDWCw77e+Rd9PePBewB4Jm3RoaEe+fkZ3d18sW
K3Ojs2qv5UV+/lsTlHbIgHyFaVk2cDkJ/HB+mNXIoN/UbeuePvPcZ7/36vw3q2anLq6PgdSEghqd
7uQH+0reLEwAM82uBKaDvPuBahVlJmWPhBoCSBDrRtj8/SFJgsKc6ovdgLuFWOyx8AmcjGL36bfI
/6DIxAcV2hES8mqN1m2o6DDgIh2MMkQAFy1QM5GQ8rV5KM3iNAmR9LLSgy+0m9PC/qBurlq7gQDc
7h1ZQ+EXq6/VKhiepokLEEdz/im54Z0cPs7WkhsdjCeQzFqpFXwXy/8IdGe5sbPDWGAaphja1tuu
uIIWlvILYAJNeY8w+2lggOjSCwaq2vZQUftqtY4lHLfc8mmkjNf4T64pLp/cVMJN5t6v4uBjUXf0
B07PI8ZbKZo5CZQglCzebT3CIhuGlk2gxMj14eOcsjERzJ0LymNQh+tY9knLCMooGPqKeIN8lgzt
tK9mk+/CcrIaRwTZ+4nhLhla2BoHpxxJfIt1R93RG441GsR78T4fNCNT+6aL0kf4xkV7gO09l9pZ
MwPSesfmI0QzSslkQK7kBReLx5SherQXCEhv0sPsE8yFve57TmREq0TN99UttcXJKfwXWgsIYeod
rQ/mxrupBLetg6BuWhqrNWg2VSKDqPZZpA4mPMFawyuVr3l5ntSedgEtg7otolb+eJtEQL2JxWI4
d7N3FOGJ9cJvt2dLvsv/IZ8s+3KObBsHdfgjgfTJnbMB8Br1HFpNJYH8NjCMI5YXSl9ygN5fRkVK
No8Qew1rdtFHQxMzQhflq0kX+ZlMoqpP8B7Aqtt3CSRSrvyp2fANx+QNzy/0JYu3r0HgYx0R2+UG
qWCbXhzJbkOQlGVc5dQ29KexppXo+4AhoxUz7EB2wSi456v0hqwf36Tm8yM3QX7G42sFgVHqifpx
UrKMjCGkAnKwX7juY/RBz63ySlRkCKVFlL8iPJtShb/BXDYcRuNgUR69BvN0hyOSay0LJggqmA8P
GiMyM2GV8G2QSDC8rTDjeHsCUIxNujCIbgnVaYLB9Gt+9DmwRpXTHHOtkRjvX2k4nGxjSJGUCzDK
TBHW9muyYoWNC5SK0nSmHGb2c97Ej0zYA/4lxqkgFZrzFNec/K1HRjaQ66MVtpyKkw/Q55ara75K
RNdhP5n0y5rUcKePn0C0eaLv3MiHaJeHmjD93aEyKVEhO1f7EGuGIAe3ynJI4lK2dBwzHCkcAlGt
/nAPTBSrzgI0iHZN2wKl/BcfB8sS4NfO0n9m0+Jd5hdAnUp/xBdzxvZmUM2wuVp+3N9m/5SQP9jp
YMKPVF1cJNT8z+WDuxwCJebmQtBp2m7PWshrxkJDrXzMobQdlgxU3R+NT3CdXM9Ejuj7R/fZpJR+
Y5hyNmvM6NXCGKYIvkeRFjR8hIp2RV/GJlTi6vDFi+/Ds6vBgv2U83/T7UytjaYZSU7b+gIbMryl
5PfVT9MnaPqVsJABJ05OGpwVPjKsSpIACmdfGrd/fX166L6bitLG/MH8F5W0fF8ZpqLXOK6b9rs1
a1Vp2t11phhZK8Ib73m8GEy2IxZYJcWD4HnyGuT0xTPlizlns8QOAQI7cCTF5M40lfoiBFj8ErPa
9s0U+TIWUN1mfn4Xj5OMjxIgn1NGTLceBthMdU23Zz+WSGZ0DnQea9O/+E8d0sPOJSUO2m6NImx1
98GmYaOBDMA+9JRUhcYDQQRNdvolXsL0I/Uc7Lr4DrnRidxu86QgmKKKcrsZrI8MVMUStmW3pyM1
rOrGlPFY1QtLb2Rbhtvak2XsKjej5aMqzqukUNX07FNZi0nnIvK8upYFnhqnu6SOZ5S5bxn05Kd+
l0/e09FimE+ivs8JMGsTP09ypMmCaeHcrp0B1rtlnIeX89OJmwd2/+vX+NoAbb0FUsZ6hhIFTK9S
2n2TRhoUzWm6Yklt0ieAevyTMjuxRHmnP9s1fkA8AiN3r6SNyRMCAn2Rrvk5jRew94k0BqpX/WsP
wIFSlnV6XW82rguXSjNiTBmyDWzmG3Gj7HuhtPU/qVjIqM/Yk33k1s2EdigwYuNRNo2U8R1Cts9h
VxRTTVJu7DvokrwbMnfDJ8j+p+ABSPgYdJvBYubh7JIYwyjCnHB3UU88L3PcKjFpFSXLfesple0w
GnFM4A/QkUyMPOYeab+YFoJeKLrBZdzCMFxdV4PMedOOeVoqjB+Ppk43Rj46f2hV1cX8fFYHA056
Is5/cDzEe110MGt5wwj4OZa0e8UIw8uZjKuGZx+9eC+mZMrNpz59BPptEWfbJYBKSRgInkMFUP6J
42UvXLHHVQJLkIPBTo961JFLVlPBXZlZGJbFK4qz2NolxuoHgZkBtC0VrMx3KzRwAKUYzLabVSAs
bQcOtF6563b1F7/5Xe5pHFue++eHk1d15iNS32j3Ad0hKKiKadTom+rjQdXjmE2g+1URz9bLWQec
VbGtZayDenpNjEj21xZ05WFPvNKkIy9b+uITvbFd866+B3xgUDVlxH/Ra8ZxNlL5yVo/FMSfh8ZD
T5xKBqNp5UUvk7z1AnnUNpv7WHXiGTb+jzVgdFn8qJ/zJcXF+6ELjVGqa+rNWFyC0qYcExesgST1
xMoANR0UhjegeRp8HI0vIqjlv49el6R36HgABkHnYBgNSOz1WxqX+fsSD3HeT1o8pB1nV2uhrnDs
BnhFJgcWLqd34j3yIglMqr1Y8y7bv7SRx2x2hdbuqVTDFKyCWh/GO625fbEq5k0lhHP93oqGWn0j
Qt1B46VdQQ2J+ksY1nuakF9SVScm8H5e7GI7f5M1AtxVzj8woPoDfRFpBy6BFZ9VEqtCmIEKxGEw
PTNm6yx81kxzTYwbkhxqc6+vL8yL+cS/hPhWMY9BBQa36oW3TlEcLseqQhsxjEkMFqLFwEqMyw/O
z0+CD08NdNl0rT5sOXCe4Xcn721wIbKcriWnWoyRZbfop921qTy9ri1UiirSr7ixzO+0DXBbks+h
crSvKXDn4QZgVhvn0iRjmbHQxJ9t8yTkJ0iFWMEYDbVY+6eYzLpoeG16lYYk82/1U2GXUhvL7o7k
rurAJocAxyp2z9LuSx6GlKMytkmwSGUKk1iHfDwZFz1igqpq+TFVNbEI3bou3dU9Lw+X6i/FCJkf
C4p8aU7X/pHTP0nXxnPMMsNhUUnJNsMa5ceYZzFi9RPGOaVbGqy9+9fBN3mOy6Svjkf/Um7gTwLt
8B75pMuvixxIplln3hKuIh9GWyExkkx7wqotKIxF9ZBK5VDhweBU5q1wKTCOEtjXx7uv8UtOSn+F
RXdF0ceX4UKHcDV89AuoubFQd/FtpUdRNvD2nObiK4mzPjTBZeVx5tzbhAJdd9aUZkTmf6tJiwNs
tNAIG/2iR1oolUet8JgD9ad1IwWKKd2o6kHRjsgHXqx7wGmwJcDC31k6m+TTlfDEtS2w0AuaZ8sa
L+SjMukiSv/i0Xk7lnQR+yt2CeftymoRBezcdYJNcPIA+66mxMSoVv95sh8QVsDUw3H0yvdzCVVD
QAD2A3lc7q9BOqtR3zNVjJW4oP6IGI35xosuLyNRjWtwAUVh3hDgWlP6iLoiPJeJit9Dtmy20IdG
tAJs9J+qpS8emVOkknaym35tIyhrobEBHiRVqtbth63mzl1SEnQY3tlth2PfQxusdoPuQLbNRNiQ
F72f4Nwav6Z50uh5d7qlQF91GhNKTXjRXRobkiNpxbF0QODFKXDjHBfOqUX+823J29vkhTRkWV6L
YbDkJlrLSt1IwVNMs3rlkm6ZDwy+fVYygeFRRqXu86PRey0ZDv7mOMhXETlQc2eN7TNSPV5/y41Q
j3ljh8D5j9ehSSZyy32tF6Ghzhuu3wzvkzHaxQOBFQrXR6Lt7bZHOcYDepSN0M1EoZ3QP9DzbTq/
/cGEklgOZZ40UojwgC87XYqNne32eJdKt418cOL2mXkbbMiIxOK7Mz4OBdSvtbuSS1u8KOKDVyPb
anDRrrNc2vWXTtmJdNlFIqLRunHeOAU/EDCBoUURqIEDzYaYMR25tE4NCggoUyimPNRir94nCW/O
vN/GRLTZRTxhL1BfJS2fbc9tnKHWPWGVYfi9V0MqgSN5j3BpOQnjwACuiCRGzBRYy27h4I1K7Awc
n5rfBXvEDuKiGYwlsrGLdc+0PhBn2AoCuFHTnCOpM4jvgBwp/tt82ODX65DMsGrp9/k06Z24TvEG
JhO9Ji1KkUFb2NfNAlDJAUMf2W3gPLIGRFP5NjgcWxl9/AOfUH8668mUfWFsdclM4NRBku7CGtkb
5WctJSGPURKYHUfxdEhcFlKfyYyqSpYKRiPXQrytm0u2O1XILcIlJXsYe4b8sEK64OYxn7WAeKu8
Xf1SNqD7gX4GiKP3hL5ZuhPUZOpx1fUZMkZM77UaVZOdnJrCYQdL2jPB2WTFwsCJdH6jALUg1C2+
wJcElOC+1+zsR7ZniOMNlX5wzL3SFP27Otlf9dfWr54ga9NPYrI2AIqerGk/+G0MOlKjgtl1lTqn
MM85VN/qLVSEASQUBQtqY0BFEl33s8ERLiJvnDBhPheNZLObIzlFVWSWe0FEc+St6mmjGdIdAWc/
XxDRAHsqF+boke0HHANDcZTbK3DK5sFM+AXvWbfpuwFxrZuXXlP2yxxOEQ4jfgFE1Y9Z03u3rfc/
PM2rcdueTwcYsB/Coa85YF6arfB5dUUQdxFQm4ia2Sm22wJmaW/UwlTqGhCRZdBwlDEtBj3beVQG
5MKe5jb3ICU6MsQGr0aEMfjc2vEcE4HpndV+SoXJ5fMz/fOzGmt7bbEyzBiSGw2GBTl3kyTmzkw0
8HsihkcfwzJuhxaXWrxWUoeXPTzJmJScKbslevgQqIXbxtmiuoK/yiPn6nHbycK9fTKE/f3UZotz
asF34g6YUjdK7Ux7Yhk2SqjNl+YVTQ8HEGRyD9WObSAW4I1ACqRzkL2n1tFkrIRHTUFdz9/5KC8L
hCIu4UkWzP7nc4bOR1ZU5hqjwzszFt0XMVbZRFuXbhxKYHrEvx8w8vxgquyhuwFoJFpeiK2x+a1b
IK48hDz42vNecQn6CNpe5yesBynlGpW4CzwzycrEitG0sGun0DXIIEsB0x2VvTah79LlTN87F6h8
yWx3lgiGO5AIKer9wAb4kAr9H9JNlqtl2afxdi3rlZF8H6DBP5dylTCQRjOYdhksKi3Hu/xcwmx0
ShVBJ72wqVo6t6ZMgQeYVSTRmaNd3TYqEpTK5MOjpF67UHqi2VZ9D1NNTAdO2Kl5aFLYB1snKwKW
RNP5gZUS2gdzFXLjFevL7YYsyfqs+2YJtLS4gmQD+HZg/bBI1c3+cBpkA6q1EI1YJBGrANNt/huv
lnYMrUeJx0EVz0lPO7/ON6OaiReMrAUyt614XNQtca5/dnRwFcso1g9ci+WtmukeE3kR5lFBnYGK
C4gV0VJqs81rkNaVjN6B/BSjuACSblE89bszI/yBRDlE3aarPkjpeI4e7yLhSKJgGSCSdFpbx8hO
Ks0CjFItQJfkvJ+Zhpwhp/DCk/CzTQmqUG/jr8HUz29Lj+P0UfD9Gn9zyKVsbmK5q+ECJ90/R8hS
bjni80VWSHz2ZByGzXPp+SDpIXD29RRH8qZBjKT2TGcaFEXbpMVYnozFK+FhB2G/MyC7PNB7VncL
7zf0OsCI9e1tT25hUhHUOedegAiaKTTBmQfarlwH2mRJfTUWH8zrB64bGE6v7brzPboYzt/KmodE
f156TvwJ1IFnuEkmZ2zb2Qv48olLicOox+eSkswdsnahJAjeYo+n2gLaKBQpBcR/N7N5SOxU8t4E
6FK2Ywfp6+nrhmSzglBSmcvog3/dE42oNYx2BU4s+lVj+0Jt83gv1LtDLTNOPHgjvELpXUpKnhQ1
C94+rp3ybzyZlYujgDiRBEigmjwmhNrgq+ncPfRTyMh9RtDTfIEVIr+7Ugou9UacWkuZm9zZHUJ2
ifnTtrO/I//AIH4wngdG6IGtpjE6kPBaqVRBzbqxhZqqsWTrfqKRAGsxRtXVsWp61KlD2xgUPk/k
znY6rQOqMcwUol6ujfpPTEz/L5pzzbskZFpsVSkHV6KMfxpZ8biZuTkbKJiW+FzdEAqrZSJ1TiTz
XVjtAXF4Wq92U9P8wusQ9PDmheWe75Gnbzu1wzAcjNUVPD3nxgbPOtFVJi8rVIkau2kXz48uETH0
iVfmiYgXC0Nz5zqpY8lNxOzUv/U/85ZeJHA43XVOyYqvhi9FBYnGuy0yvGLcy5mQYeItnOkhuujD
nU86Wy7HHZBNI7kX+woTfgkjtfzecX4bF4gK2+xfa9NShMMfk+woB03g8boOGscUSEIqILJXF75O
anSJXs4miPBPDFD00JR4gTYxI9Xmb3Aj4v6CzrB2fg6KT7L3RPzzeqLPPk1bSS3CNJfRQsq3hm72
X6bMAQH6xojex2X0atGJUnZrSGJyxfHjTacglsfGVZP1HGNQcBSQ7XXrozG+BukseHTjKrZmixp3
IE6chy0TUJ+3Aa+rHySe7rXg/yvtsCagmjgzdhBn1kv0NNbiXrUiS5BIo4H9HJVh9VyOpK0EqLwd
tj91KpzvYKsVXwuzufyZ83nvmRwE+CP4k6nxKj5v4Zd+niwVD8LeuLbpGMD2czxOG6RAiz4Ng51H
WoOlXzgtxJAyBJ3y9Sm4NZnf49hO9QfgPEdccDLanA7BWg88pAu721xoj41oJw2IKA+nPLSA5YJ3
wYZEWEeWnG5/FOL26peRPG3rCS4zTtRUeJa8MssMXPJx2v+7v2aHPQ85or9eR7NEArqLTlZ7jejn
FkXpJp7xPZpVO7BHaBwMivroYeB1i50Omp8Yn0fNMC3lt1bLZtCDowq1Z30vXAWIF/TQWF1wKybD
zD/x6maolFOC+ZKUROBd9Xl/xGkHf8+h/sBNYkhstLwNrmjI/udbGJFqquuHj+mLRtBub8rKIcGa
atw3gaoCofrx1E/UWpKIucKf4Rvs5hStjEBRu/nLZ2GXEux9V3bYPiHtZeMOCVifhSSZfd/pNONX
yMSIKRwyWvtd/QHrMlfUT6FBQqiFgTM1YWX8tX7hiRc1wJt3HSaJuVx6SDetTuWBfZYlNiGTDoTR
1U5YIMD+nxRXZO4D9l4zahycpCSriYHiZFb4exjRJyKamVyDyhsTH/PpuImesdBaNjcPAeR8iCCf
FjKl6ZaTLUZI0sukPaqAnGI+OLfwCn3UcrGEPKniEPwa4ARuaXyzIB07RcIzvibkD8gNLYiSb6ll
XpyV9RtxQw44pCTOxO7sRlKp/SKYE1nFt7mrExarnOcDQatJg3ImPJhSolwMr5dNFTojjPo1AzRz
kfZpKLJPF8+OefaVYi4Ggduph4HMwS2Ez0G/eiN00A9XJ04Hg5dnw7ugiYYg6gThlUFQDfTgCGkr
FuvQJJp9QyVfObh/h99Dd/BmXAJJp4xR6wVavhCWxW8tGBYWrOQj3P5qYxXLfV9mIZwqdAwoHcw/
ta4iQ/O98Ie+KdNyRetp/rinIlkan+y+cFfsWUDVy+Jl/ifazuULvH6jMd6Rqg8FNNb7quRREoXW
uXQJHC+Vu53suFsDkmBa7328k9O0qWvtW8dE+5nIBvBaTO2D58OuolbSiuw5ybTKv7fO8JgD+ZAc
UIFieavGucGHB8TwETZHMl0L77GOluPaTMyLvAhGUAUkgXjQmUmHekrbB4J3dlS5YtSQEEO4WIrT
2WR/KbBfHggSZT/kUtN1pv2hbkQcaEIR3mE5aPFYvx414At1+bQ7jenBHyceAe1eAQhPYywOQ3jl
GAUCUgR27ezJ7kQxf2LhilJLHV0zbrOps+X5GUF7xhM9V42IrhGNEG9dR7VVUu/FJ6aQwuGQm1ak
uvfot3sJPGFNqB0WcI3u+8o8q+0tJr171XXrBMNAG+XFQ9TASs+1hsSgvwK8dMGXJQbwfSj2LE9d
3wg2yNI/hJH0Z2SpNYP9lTasQKHzg1WchjZxrOOqwdNKsZu+OC2pg4gdhiqcXFpQVx/WlWJNP8t0
AYA/J+RWAWWjNRaPnHTwjGMbxN7+eK4cSxmD8ghmSLSWOOC3mx4VXSMCGxE0kgX8Jf/Pdj2dq7f6
8nJ1whKwy9jpgkfvsW1irso/D6eNxeF3nrnwBfUaveW8ug5/N04m/T81Y/T9/SzCzX42EylhWO8b
0m0ILSSYlNh+7Lh2VB3tU9E2CPIxSGv7OPS6Sj8bgRMHToIOJsccecvgMZT9blrLdgeuViQwpLqD
I4eX5/4KLFuvpo8Zy9WeN6qNcHOch3CEWf3G1vVCzLH/PJ9codJnuNWaHOdANWQ3wu7Ag88StXz9
sbZY2rkchA1wQSjk1tB++P+Jz5wvEnD4XfDU72ax8ZIvaND4MKcFrCcijEBr0/cj5pFvr9WB0yk6
JcrDHtUZ6PORSe9fwSwh4N8Rr5ECv3k5aF9OYLRd94QN8al60g/n0vihaWhxFBKwXCWWcuFBQ+p2
pxGuFyBEPfsV56i+DqKoSki2VvWs0d+F9m2PDKOFs2ANRHllWYKjX1tD1TulH0G7cf67Jb/QeDRa
9OPcyuSrQ3hNalWh34TtL2A2asoK+I7LM/eMuXexR1+eO1+OdpDUhqIGoaD5F21oSRa6Y6+R8sAv
aUGZR5CZ/760ApEkW+th2bNwOqRoFQoKepDyYP0OV/ahcac4QOH+Rzx0tGVpso8542QuNMalhqEP
8NNNkAHInKLAtzmxhU8Kmny8YMzztMKBG0czA5fwAtIaAX1NGwLGaeV/eirqvC41vRN3pppGZyN5
5PlJWvM6iVQvHBcnN175U5gEZhgF4buxvoVQyBqxob8n90eSfiIFfoBJatUhizYFxovSI3s/enxt
TwKrUMfrBxlakBMGqeMcpGTVXEJFg1IsirFm8LoMla/wGUN5BHGKUVKNaZkfrLbXOgePb96pO/Nv
jOKIYq+ThuNf0y4A47hXjeGNlOCGhPmPQjY0q/UCiaRzzFLEYPvV1vKi+7bkut4/ztw4c1UhWrCt
Po1XpTHnngnnEtK/yRYOKAa4QulSyASGL9laVN8pI43J8aqzMLvFOqRTaxWZLW2GiSm4Ec9Ku8T/
GgeQMDuJ/4419dbBNu412OtHghPU5vHwigEaU519DcOwHnR+SVYeWdrMqIXFmLvQVDQW62ZjqciU
NYMyC6Q457shHIP2oLYmpaLlFsJbanrWkwy+kDVtZ/Tprb8r/5Tl83m8Xmn+kSLvgrEHCfurc96W
hMyJT+UTPcXrd+P3R3O7mo+qT+aQ9aN3Ct7d6T4muKi+pRkDPNNLK+M3vGndA5lfgic1ApXjdoql
hby7lO6uoQllqpW7bhGHAdIsw5BqsVLIqa6dB9LxvsKtNYaOe2Abt8wj6ZbNWlWzODSOC2khVnE7
pmhrQp9RTA4Hu/9ahw9H5sguZG8Mp5DwzWtqIQK9A5eHQWmf7pDMvEl9LQfWYjJxKP88d089TcTd
eCFDtP3XfCzeFozRUUjJm0rajncdBGRqWhQlT8Vl0AeoUWajI1Fxdt0DyYXgpiBxKn3LEuI+I09k
AMSxA8Yas1oIBKDb3RtFQUqriLSIUiDttRFjua2FFRp0eSOUP8f/+oZ5W9gwvnJdi2d0fVmWq4Qd
ljxpjwop4zynJniaARs0uVrwSs6jngvgnPp5IRYAcCuKV7QAhmaF3fHScOUWsLSIUy7/PFCg9u5+
/Zus9xudqIeJV4HsxuBDsq1qNgK2rSA4xGrYE2TfR+F7NpIfWMr8FMqluL1UZTTz9c9aThpyqgFq
Y+9ECdeTvtbzelAksdk/s9clVpNcK8pa9D6Pu4pMUzLIn0xO93bkhegA+u0uHtOVkws+qe5wIclf
XSCZS/NbBqCps4kXj/kusM/6e6aau0+TaBkIyEdVCUyLaMgkal/a1nVWgN5+SzXVfqbLF0pfTPt6
Pe+Ur7vNQWACxqP9Vjlbf08JWxnjGU1zjJdQbeLJ8/Gb0eYrG+KdwQzYMOcmx8PzIGinVVa79j0+
Ocu/X7OV47hP0OC8kzOQ03M/+sLhdgGM9xLnjgzkjNBqGEdqB1UXZ8KAnIPOi24NSsh4bYDgBQ3e
rkHzn8HwSm8eRoAOT2gqKBPBq4LU8Ho9wqE+5zCLSQGPL8qoX/7+hS791pu0/IDbP/Auy9UkO7Ij
Vku7Eur6dDopFlRVAjzHgAB7yacBxrJBO3EwjDHLI5Yb5FA2xe9POCdAtl/41Q+PBLC5atj0VW5C
g8CGhIKt4WH40Zz1oL/3FLi9fwiQJrSlWmLF/iN0XqXXR5dJtfySF3tLcC1qTexo5QP4LI1NckiZ
4KISZL46tEwpm/17opsEspjiFaxT5E1258ckwe3qLEaOXQ7O8rY9yKMCx8043QppBG1SDdFTVoFi
n+KUgIs3If1cSk4LreBK47vx43eId89jsiWK9D8CnBEoNeIOeH6WE3p+LBr1LGd/BkfNNeVOxdr1
/gM8qFn7dMXhWJNIKH09n+rIe3xm6CDKEilHBxZxwuSQXitzTn8vbOyATp4kAuywP5V+34SM9R+D
4Hlaxio+RiB1ceeo1CR336Ii5YQh33xJULX1L9HTabzH3Xc5GtfJ7EfJcvZpFvU6u91suuIi0Qb2
txrSjMnVzS83GuOxm/3dNmvfxiq2QV9FbTxeQ71ThKwmxa6psxrOkHAOQ5XOfOR4f997IYR2cmAW
b9zUJlnrVjbzlNi6gyGqBWqGtvTlU6BWwHmjAIrqIi+Va9Zc2Lnu3WW2FyGsqCBWPA1MwuFZcS9/
Y96uXapefwd+1dJz+cLjWFVBSS6lY1p1k/l3Q828eImTK1yAIJCARfJjKTkbjNy20BqpqVORhv3/
PM+WOsMLKyoXOAYZoZ5hPdpO/pSCduU1yfe5FQlxTi1AP5CVcBxhCc5ZLnvZnuga3OysBhApCBOg
B/BCf60v/XaX/1Q0LsW/jJRfSttx9vEx/bUXciLQFQanf2TRjihS/AFXRkkrRCtV6KCgnWEe9qEJ
OImZYNSFWlcfAH3OcD+NYUx2q6nsA8C1VOMpJ3IWvkyNlB1zPOAw+szQwSCVrvZ/TZSFih2ufIYG
ES3nKgTS/wogH77r9saaZVag/jWOCBZqHov4EDO/9xLKsr2MckLeNwSFHOADjaOc0KvN3F2ueCe0
Nzn1Zn6cEQXsZJbl3CFeOHOttQ3Y2A2hdl+wRb2mKd+PGvejWIxlln9XknlYMW/jpjDxV3x6PqeH
eaaXY38A0W4awCLRISQv+z+evISwV0sr004cNS7LN9kzZPXgFUXaqe/XDkvKZyc6oHC/AGnt10Qc
1NRhdx9augKolFcaRe0egN+ZiilFFAxlABszHsGIVzI3fh1XDHiRF5fKjBU72W+XADUVNsIv0elx
D8mX9LPq4KtHPoH660/gsdzNryZJo23OFtmVp5+qP2n1bOiWC8JovUNc30e+5T1KDjC3851tf/bC
MQay/qSpB7cRi+IKcXP1SQKWDXQ9liKkR0hAfWerneORGGFMp0CaLpqUxI7R80ATYlcx3wjaZD+M
GtGDReXr+QLjP5hm7bfgqk2Mym3DOapV+wdcDXxR8rtAEa6+nqhV9CIdWWyTnO87+CeAGPeamEL9
cvqtlXJU1GeajJyHDnGyK+HW7zO0OfcdnLwXQwktTja57kBXrl0W6f296Gx2R/RZFlNUXHdSqV3A
luAUSD9Kiu8UIKLOgCuRyTupawyMLsdKKgdf7cSnteLGvQ4so/sL5moKMs3HQ8sTxlDxWiXWFixd
FBZ6zYBWlqpE36i+m7uz7E7KD8oxAyqWoWY/JYeKf97pI/cGcT4IB5lNlDb9l+pY0q3tGJ1tpNxT
E6tpOijhutQ3Z4kzfAFb4LLhCphqdjl+2IwGzuvrvqT8n7dw9J6NOQjp54xFl+SRVw83FUnjjqQm
xdPiItop3FQ4c2SaeXk88+TrfsdbFdmAgWqId4VFuPnJ1374RCDX6akhfhYiJpiwNc7EM/XeWvHy
EaxdVgbjluMNNzvaFEa0mGTLm5xWBELUKfnG7+0S1PrmojrI03+FgI5EWtFBLsTyfRP8Em5aK/61
ASRueybMT+JKO0Ux5rohNeFZHq2sjLVPqRouzdnn79mUix1WGjeBrwQ3g7HvaZTcci88MFzJPvpz
ezKAVEgMbGLddMCeZrMZUQqFlOxJ5396jJ4yB5QyXAruIze7Rd8iYwPQvVmQ7v2tSOWvDsKToF5J
6MVmPjOt1c3I/fa/3PeRVaWD8uIK3V2duFQuS5au51hVEON2iLUONI5R43K9nWB+4BXs4UOz3WMf
abjUL/v3QmbhLAV9SIaxP2uFY8vxanJgKzhqxpolarc1mO2dDvJqrSRYqlidksqgmpbuH2MnV8rH
hbsFAvdMO/vRltIT+70ufUIQzV65/zNFv3pFWiJ/SqIWfkXfcPseD8ZQ09r+qaXaHUQxO0C7m21p
Yo4R5xkRv5XNvOXWyZ8OMujpvJ4BEC0bzQvVNiFpdExvU7klF0tV9JgacJvmBDUtVuFR+bb/enmq
iaykfbyxwNB/HP25Df/wi3gNpO8HzWBtKd2u4nm8KjR5/J2kT+atcmX/KXLMnG722qusTW29iIey
0Vvtc+ImVGXuCyddCnpH1gAF6AoUaNjaelYZ+aKKvgSePCrvmZG+06XbX9yqW9EL+E3PEuRnIcEV
wdqmyC0m8rRwlgNo2hCDe4Y+pXO4W5GsyxFiUEOYV9FKHq0GtD+YeP0mibBWOTbeB6b/3/bzs2ns
ajjCVlIw0LMes2VPlz4SoqSL+MOudNJBzMp2iWZWmjosv9tH0bra4XJ3s9e2Y8J4aTt2ndou5YDW
/myOy7OvO51noC6+e0CrH6DxQINjWkQetCx3EbNjTgyMEJZHc8Wisd7CFV1GUU8fKuTtjJpVryCc
RiLkCVhvxMjzCs78CkhIOAh2QPwpcnEhhMBiTVNGcWtZQ8WqyTb7+mymA3eQuUw23lkrBchhU2s3
0VyXMBfLtrhU0Pj8E+2tj0wCPSriKkjbhJLYxt2pYAj5b5YwZlqUo+8owTQoFqUeyU4uTxH7VkOl
pOZT0A5hJPnXGDIaEPmnqSxgQ+vtgzgmzxvoqkhQEEnMfp77qfppFFEzXp077OVOJ4I1EZr2pY+t
vUOrqSk6Cd/kSQOPmhlq4kOJWfSVL20cnHLdWJYjzRTQmBhbdjzmDJygr7jeD6HPkvp7NT6ZU6VF
kVqS2OgFh+GimcPLlIjM4P1wnSGgPqKgL2yraODcUvxBEzlnHJwgzZNt8gPg6K1Tv0h/SKowlBkk
FmkqFwPrwOTkJu8+lIJcI55Z9RunJ7YS3QVmXq7jwR1Llc0tGS3qFmN4Gxb5kmZkEu95qDzW991z
EE3PSTZ1muIg2Dbb7zuyTyu3EVKg8/alpaZlkbdkP8e54SWENnLaG3y0vkTzThu44Iqx+0LJz3m7
EUAt4ef4oYGpcIECXE6GXlbmL0HWKNpIWiLTdlTBWxybMRc9vXNYqtkWkoaWZtB2AUxiHu5jQzrd
LGmPj8DRuKDrYtriGNQz+KfRpWpB2HCojfEC2MkjonK4br1TNqAjzzHLaaK1yyeNQAaz71XHR17/
E6zZInHkF6e7tytYcvGliLX7DIlQ/SHS3NKHzyA5UzIUAtTdhXt7YvBz0sSMWW4A0rb7KH1/oQW2
b4RWpA15+EcZbo/rGjuweDuKg63pSEGTrLD1ZGM0SXpyU/scIS1kdU3VJwt/O6Y+QG2FA008rO3J
NhUMcU2JXzV3735E5144nwswX7SlS/8rLFOy94lwaPR010mlJtGkxzpXWpm32v1BxTAIUq5+xx2X
a0IS6FPSrBexUsU7PC6TKgRfeWUgTxSOs2Wx/Z/dZlDZ5v84HI+kfTvBFlcmyg5uBv8ilk4j89Yp
dRLpuwFEy7UiquhXcdgsgt4rMqFTkO5snCLlned5CoBLSbEWzojqAA87HNjLLZBwdZYQ6YSB/yW2
VG2kBEzcWmpDnxSt55LtOz2OzW78311sfIxkgmdbdaLMzZIziTb3ts1P0C3b/YU73ej2zOvayj1X
N8GNr5IdRGH5HcsmClTl0UbDLQ3YESo5HQE2VcPsoNe6XDbZuQO/Rx6zv5CFNqCn7VYAV3xJpLcN
Sop4fw+JLhYF0mjEkAeejjpZPiuXAjaIE908LTzwh1KECNX6Wyt+3QHLL9f0CtaK9l+Tp+HQm2fu
i6i7EieLI3QH4lhAbkdSlZS6IYZpVFeA2psyyRvzcvSYPLS6V3nWgfoPkCOZJFl8BWNun70sOjQS
XA2+45iYqGlkEdPVyiW5TwPrdpR1nzOW2/hRO5Shbj6GSoUuBwqgGorLPwSKUW/w8+XIyocE/RCU
7A5u34WH5ahD/S0j5rckFQfYXChL+7DJNtF905bZf40vgqFyq2k5SgHosoGZwnWyecZ4ZW/g72BQ
XDvgeTehq2djPPAxqeOV0ojK7okkZl2n4PjYUVHO+D+CouqEZd3vh4EzQrlaz5RK4C84a9roeZvx
X+Co14EEZaOa24093/1ibsH5yXIavKAHC9oa29X+Tbk2fFoMulQtFmx71zVbq4hE4C25KEB6H5ZC
ewElSfcSjfR6qZKScfgouh++AVcRi7Rx5QSvydHkNmoL7yuxhsLQEamRQ1x4m/l2hp8DNP/vadf/
8TbVYctVoz6EKwOo/PknF3vMTFrW8lu0xqDMY2wzzfSsqMO19GFBQ3Ogxu2vZZXB4eDiNNX3DIXz
HEd3i/tH/NczovgXOHA1Kh+NcBuQKHmZFp3fuT1OwkxGrFOIQ26/J96mnVkTR9bVWU+T2lRK0YhZ
xvght4FyJCs69Xtxt1Lc9AMEAPGcgefhWiayXnh3p5+fPCGSV0LDtXykXWzq5GFYclnDIinE76fy
5YSxjISAHubQOr5V6h6cCMgZ633ylUqvv2vRJUINriv3mtZq1h2tF9RRIXYSQhohEfyZejZyjs23
cp8DNN8A7Qc8Hx/OOrs2doc3Ad1hF2FAMp0uej5nUmjYfxscyKveBr2M88uG/rQeci901Kj1QuXL
AKu69UPzcQVwVjUGr4Uab/yeRxePksjuL3vnh6jUnm9Dmb4rDZL4FOSPbuIwQvcffMCTVa5ypUBv
U9oW0liZdoob3zlm69MFIf5l1qKA7BMbgdLU/dMcPYFHk4nEizqipkCzPciVFWf/3pA3tsfO6pkC
1sKKJZ8MEPDVCgxvwOAXmD5j1qTvDNCd5dJ755hZo4tnc6chIUMpZ5AP9Uwu3vebsjtDs+zFQt9J
nGmlQJQikNArW5m2MejdxErY6aI4a02LVbRSk/IsSAoU/RCqPOEDcC4agrJ3dVB2EDqruR5WsF/O
1XSLGI3pXHdzJIon+abeP+wrWVuzd7ZbdU8WFAKEZYZs7brx0qSnTvLApx+B5pHDc1uS6FJqFLJ9
6vZj9WaCWk0tn7B4k5VM7WemtbyXiKp/GVziIOT6rIMX78Ra9U0aJR8o6iU/FjoSTysPl9StJFDb
PobD7Qa6ucvf8FjeCY/4JfFJqGRnB1CcqLak+TTTInIJMYfBkFVhTpUTRXsLL3bG4jPlvqSdnsbe
6dg4Ajyvyuaa9n0Ol/llv5lfjlq94SvvzT4RIzG+sRWhV/UlsvAyNliIl95vsdM+GA+oX5Y5X31+
u2Z3HzQJazy61dZ6WnRnk3HkNanjjbUIUXASwPWcM8MANfky8DhxIZGgwibnkDTiuU9KC1Fyq5Fc
fMnsl0cheIaIrRewwXpZnGebnrlOJPwHdAXi5dPejUt5QD0ewRDY3J7bj53RlAgnLBT4ngj11+a8
der6JGYFBRY08m+RtmYF3T+wjNX+ldrm9ooL6H09e0X1s31VNYu8cG5myiX8qcGJoCQAfCFzu2Ru
UejhVBvtZHYl6rl2TrbFJ2CxFbMapK8fJtVCSNV/OMLDJwk1R3uIa6bZrNbUd3FtjWXOlrqQmPDs
ry81SQhUYGeKtaJ198Us98JOGWwASgwr4KuQ5qUuaTelKZgJy2gs2ITUutbYQRzM/qISFtbt7Ak5
LADCnJBFgtI4D7W6Mkc3SM0vf9oKahBprIlari73uovis01c1pPuCAUlXylQl/NNemJHuUkAG1mG
kM5U8ua/OGGNcrVVn/213D0qnKoUX+xFMkISqDzg3HPMfRfFEDDMNYgNARpnUOKuIqK9Il4q10T3
VGv/vXUeL7WyL/bPrr6peKYwIt2VKxP2KyiAzykFzZ/8uZrE6TIk6ZGRxmMU7roryVD4V2In2yKk
n2wKFY5mrOdr1giI0LNgrHntEH15zBjxL1owmH8tEfKu8nVhQ5iZyWhyAWAlkeFr5QnJ4gHra7Ck
SlDq85NHCL2m8yuCeVOB6CDsA4IUw78HkYKzzUjF6l6U7ybYOY9gLRGLvpH9jRQXO0BaulV8SWuz
dvvsACvgZXfp3hjakkAjd1RdwHxMxE0rKejH4dR6J3UtnUIcdwkYiI9P0+zZi+55/hyv4YTFlOBo
0ChBwX8wi3ONLal7MW0EdR2D9GMv1qwLoszADeSBXQ+LjMjST+xy1Q+hbuIFw7VrlMUUG1l6R075
z9ye4HAyJgUfAwzCUJVMr1njXhJ7HIC5WPriXEVHxdhTWpdd3JahSN86KZUB7OdT6I8yMuNU3qJ8
CTBA0SwIJ7/ATYzEfmHCKBFFuwZlzIJWMgWWBbGLhMqqoglhEFuBdyLSVrs1ECoTrjzqL9H6g9C4
y7C9vR0UzJZw8/RA+UWM9zyg0qResN8y8cqzPZe/13CtnEmIDhOSO0Yo2TtNQwutjbLSiHyL59mj
d/z3H1CoNyDXD5xDohr/3qlgqfUjLG71vTkhjdQjJR7Z82brkUOSGg1ANnsz/5MWuz722fzZLw8w
RdHn6/kFglyVkxlOe0nx1p2qM4owWHLA9ZL9cMeWiBc0UQIS4EkQP/uNOEf0m2Ms1hNhdrML/Btb
KqjzMZcDk4tjsExHwh186u5b9UQn+lplOYV1osEPaoXiaoA66KOd+K8x1AdI4qTL4J6r9lNI3gpG
OXzBaPevdgdmeCgz4dSm6YMiLR+eRHl9PoJ7HSF6lBTJZDHOA2k2RLGZlPkh9hghLqi0dHjGnZKq
pkO4tXBcHqI5trETyr5rFG4QET6dmJLAAvXUET/tO1FPguVSxb45slVlXFTcEDtUZhPPOawdJbTE
OZcNqxtoY4S7nWHymQF5TFMDj3IB54Yjr7JSobU3vYmSamSz72ewOefGfrwM1UErXVkC4z8Bw5wt
0wlc2zsFSwu610L0LEthLrirNeoMX/oogv+myCxHQcFyf/GuBY3O7iPOE5Ktzhl0iFe+Wp7NlTT2
m28BAt83qFuP6jWN06H6/MUFRokzh8QkGVVkE7M3lCOB523hFboWlNFa0Nj0a7U1rvV5yB6WG5Vk
eOFj3MKi5GQBETDlf2ZbRqV8UZvLGU5T6IUgehXkOWiXtNgsJe+hcG9l6NNt1R8hfaI9ZyV1iZt0
THKrU8WDXNOe21bpAr3TK2ZefE+GxPywM+1TNzNIG4Esvh6W4x+/Vs2bohM5vjVJt03IDoOZol8m
VxxFJVsPNyzs7PM6fV/OfK6x9w3ZL9vIRqIW1KggIEjYlhLeXt2T5w4XLJ2r9NiW7SDUZoNcMqgq
iIvoJkwbaaWpGfeaJ3eiooXV6wAgzyKQDaUcIF/8OUROm4e09Y1Oe7ggZAeJmQos5nZM56H114tj
e0Sia//hkB6NkBEeyOyxDum26TKN/XH0Otq6SxDLcpwfhbL5qnj+pORXY+dMXJLdEmDBq3LxrFif
03bJlPo7DLvG0GseB2YXiUOBz7WYl+PfGj58IOSa4HCvGcKSldMsjav+lazqjKrOwxZbOEEKEUm8
oXismEvc4cmGJQZ+Nt1sudNlkhdOkvTNJjbzLHSHc7bAUwViFCumD5Tb2tkZjaPZVJSuOCH1JuDj
fp087xpt6NfkVI3D/8byzmyH0b90SagVbfJ8Jw7Jt8kP6MAY4cgqQlQnQ6/btAGU8OefoHjfbqfl
H2a8tMO1YYld0M/+UE5upbL4pSYEnKGJu6mIZo+HrN8KnjUru3KEaeD6XA4tTnHwVrL+VLoCZ0z8
QydabL9/ktMDPAHfMe5hbdvxUDCqH0TAgQYfF8OoVR0+cmbqDGq60j2Tuc1tdDuRtkaseU0xjrch
X2j6dAS58PwcJCngrPhn9gcjyVRaPA1vblBTEL01KaPHqJtYDyP05m4YWHsj63nhdO/SVWOJivQL
AO2kdHbBwV9mbTZpALAEE7Xta+NGiOXBQt4u08rGNzyQZQdXFd+xmmrtOxFIUe7JMHuef9gcQnNF
U/bQ1pfnwbgkdVuASyx2IYvs12quo+qbtB6WM/gDNis+Ie6Fh5SeL9Yrf5AKw/25aNPtNIwCcHS4
k5On4RfPS2exqAs68XKX7q+NlIWewB0uh8zO445iJ6Ogfj43gS4+lkCa15NWGn40DjJFlWJ17u2O
7SqtmP7lrzvbxp8iTvmid+86TzkkK8cf7ijavUAQunS1kAeN38Mq50Tow1+CjMtcfyhYyqtLu0kC
mEhY9RNDVhKWov/mk7bRVxmA2L13I9szfMp1w34CsAao72DHQwL0s92bJiHDNoOYBuZozI915re5
ErhQ+7lovKvKR6gscYseSfRyD0N63JBMz1/9L7gG1Jh/54/ISzZWvHoMMuF5Ykq2r9kEhZIJ7sLi
NMIu0r3jHm+dpuSZxrp5czbChTRqtSsAkUkak1KSqoPTWoQVb4pPTbt6mgswmuQHHp7+MRt3yrfF
8Oy0m4xnLaeo1SR0/uVIaBdAR6QBQ0Ta/RMc+eYPF94hpdIF/4UXSApy4BNZb9FVBB0YWgnhe/rV
ez1jo/aLahSnzHBr+3xovd5bMe5o7hs5Ww4F+nmTjaX1kF8HW/HzpQYucqZogLGVBIqju4daAP9b
Is1746Go/KG5Cmu4hdGE054W7yME55DgHRNsBaPGRSt7eZJDR1y7x+KPN8RyH+qnsCSHRiEA7C2J
PuzogW49Bv8vyraQrPWBS2lnIhkWHkOltwlGgnRDUPemaROk3kngitDcKEybo7lY68cLpIssjAwH
HVVXA+6SzCQ4jm+HZfsHQxpJgINfSXeEoHbqXS6GTHBE5gKz/F0AxL/ESf6YUVboJY0Ib2oVFisp
bP3MwGyhAOM3xel2adbzVy7oRyoQ0JhkKxK88+Nn1NoKWXyihNquc4+1v5JptN7wr7xAvw+DxxuC
/1ebNTdXtQaw4cR3xdAkIILlVI9i2+5QSL+nTUDKhuTWw5/UZugS788MJ5moaDQ1LUUwHqwjeLlj
51+bxqomSNrmjm2eT3lcNmo1sZkTXxvM4XfrP3kVhEg50JZdKRxbOeEIB+SUAZ6MzXGAqHnuAJgP
l2N9sx4hHm8fXBBAjKQ2Q+4N6wuCvOpkxNAoN+fchLPwblsZ/6Lg9rBxaSAR7X9JDKKGBlUSjBB4
8epDx129hs+prc+ZZyNEFRGIOKISySNlLOFgZ9AmDbvA8KPkSdF/wl/rjxYizjzGAh6UBSblZUdQ
goHPSgE4WAFCNm2Pzwumc2D71u7g5CB9O+ASsfjirKtF8PUEUPz2m9+TNnjQfwe8Fh8f4U9WyMi1
hsz0OW6eI7gE3XX3S4QacKeOQguPJTPSKc6YBG3cHAdOvUP8w8iroY/SRQnyNM+E05yB3a72M9IY
fdsmQlzKfMfRUQ8JNoZ24f7jHrcspFKQ8/dPk59O30+KJrCR/mGmwv78vGHw5yBYDrwsjDiah2ns
ZHdFuzesdYnwmb6wH1iEwwZFWge2yPy1jW7EgrkkqsdrFj6F2MsVc3jiDczBeNhjKMYTxJAfhQhN
bmMUbMZFwFVYpu3Kqb+xQq1lARvXXJT1z8luBKPUMUBD6ABRil7QWLX+GyzbBKUoLLzmy+o2iqS/
bA9BlaQGJlsYR+u1LFYR3AAb6AaxU5RroJqcLo/Oo7ZLjGgQiO4vwZqRIj/AWZZI3mXGeNPyS6RB
gdPQP737wlZuFvPdRejCkqwFw89x3xp8TOLdFiAw4xJhJtZm6otAKAch25r758hPFW5+BgMdp9zr
rLKCPezN38tKuRILvokiEOayCVezGh5YL9g+xOrUh9IBARwA3oYJWTJ7qHbHV/PFWYYL+xpvm6rf
0B0eiLzG2fMFa31NzBRONQqWNTdoiB8XNfT0gAJXAjRRP0c7U49fYHL6VShGc/SjAzExV1DBEWb/
lL8jKdDRmWRiOSA8VpZCPqTJhFlJ+DWt27j6RO+yH/fLHOMnpr9rskDCHZHXqXlZ01xDaKXMW7eZ
fzxuioSihrNq8SroSkJlhVC2+nbPtdMSPSSJ4mioaNzmycvlwerXoHN90uDiTfExSLZ2koUev7wK
A78ZRr+R9oe4926ZnexwtchEBFaoTi9vlJJ7AZQ1SaH+ovuJaE793GefOm5l86HPJ8Pv4FKFTtsO
rWvhwVPq5zAEs/BCQQXWE1p2/EqpGYpe3Zzx+O93Hk9JdDY0d6U/WkXUXVGy+nzReqrQMSUzBNWm
H2+37rorzmst4UYt2gTNQ8OtPC5/7ajHAhLqZkcj6Mn5EHBvlKgbpT/kJdqycQhM/WqtYr+iAb8K
JCfBI0sr1648KPCYmKJQdSpFZI4yGEiDWqXDd+CiH08AYGgIhD6nKWbKZlvmpaQuGqkRh51U0gyF
k2h39CZVckCJ0ihxZLwCcwzZtLbaPIiIsUYADqM6b6wcFxpFQWvRBpaZHgxROqL5ME54vJhPiQ05
1a2K3VYnI1bdKTxr0e6yCWrRw1xQjrogKxqz5BjjxgcMLEpP0DfVXjc7UaeUFZ2Q2aTRpH/0oAtx
M+gYpK7aN5ee01eOAIQyrC3RppL11HaaWPVyCbjfKIF1dWaqLa0phf38cS83NdQIi7zenqVJZFNO
2ftch6S8kL/A46043y0hU84ZIT2IwDlXiQK6RBje+93qTUy3nyMDLXR4IZCZ1+8Oo+Fhx6eJ9znZ
uveC41FIUgUwc6Wv8Hp2iU4MDJSbGc3Y01jXXrqXdgGu5zva2QOsbGwpMTmSpsrenzljVzOWDF8O
W/OFYbHo9MjuZPRv/TSSGEGtoZ7lQOl1TyHsIu/A1SDXQxdjfEu8LHniONhsR8nTjy1yx8QfBnuz
ugvlbw/uEHxR4C59SkK1mGSjZqWwBJOHZTPxFl0oyLFNh9x23tqO550316jWND+yXpjK4iMNEVSO
/Oo/0yfnZSV5eAou6vZHaUCP/kyoXIU+n85Py2qVTYNzTgm9ohElk2kZqP79McAabF1DRMuabjRQ
rQzAtlokwbS4dxmyu4cXMPH9nxXqFWynXW1pqG2wFFVi09FH+rpTUraPV773WRkdRHHVDsxveX1i
LLUKP8C+zFHkgBDls0kifa71E3ExYRdqv8+u+pIqHgaUbbwvSI8XQXNWSDtEGxAcSyIgQ8RrvYJU
e8hF/izmEvGYcqtlCEFXv2tOP7ZDA9qDQoAPGdwVomg4QLSLAe1PbFrvNBDaoJ1WHixMax4Wdm/W
bgJ/CEMtWAWtqD0970Q3uOWjrZmt86znIDLWnUBl034WLycXN9M/5AcFwWA+2HxT67SgAWZg17hj
1Y93ITL1z71edNJmZ0PUrM4OU2wF11eUzLe9aOUEXCEhKelbd4cNqDJSUuRrdGkFcZe1z/yiTPwT
zqp8TthGdPf0G91OUto6hg4/9fgK4vO+Y1RlVBYXc6pq4JkVLVSMGj2Y//sHYfzHN9pHXIHqIZ/e
QYJq4kCUNXoWYWchMdrnaHJKP+ampyushFTpZNrk1me+4k7Ms6awL0O6yUHFKiNE7K0g17Jdz+qQ
clBcx60bhkP1RII0mKs6Y/jy8a+JR2hjlMtwtQJbK2HXZCNPXuFNrG40akLGKqUZXCCpEEKfWHPb
Z4wPWY95KCuHkfnVSKurUKFtjKPnSuVeYExE/10nKIPSmNZ2f3KNZ5xwOjYb/5cc3XA0FY5eudYG
6KDjb0NsWZzRTma2dtR/vWFU8Rrx6qfxCW71p79lAeIJv087OVF9dWQ4wfPqcMAfEUeq6fpQFoUn
HQadKWUQ/zLWfoJ/hFnW1SJjaxCYKbmPz8RYXV3DzEpuj7UY5ufFeJ8J71hIkmfJK+SxhUhJXCRq
AUmeSONx/mi0PDxyMrZIi30vOpV5pxEwWi5+367GGJrkJOlho8aKSQjMOX/WAOIpcHs0CowDtVb/
B9WA0snSYSSj/rOd/4NG41rzSXNkT5JyeYrgkCChF4V8HnIDWy+Lt9KA/WS5CdmfKBKiexTkLvJ5
z+Ch+LpdjPOr6htro5vQU0GAKaDe/o2KVWvBRqYw7DJE/Xn7lDdLkD6h50896+Slov3CNddGMk1H
OA6Cy5nEOLlqML1Q/EMns0dHGnGCUJX8WKcEJBE/4dChetCHDd+pNJl6E3dAo+Syy5JI235woeVs
EeFY9TqGVSpWoi57oke9ofJZgo+XtcWNWQfHa3sACQXxox5g2pgkwG6Q38MbqswzVZkZH3LfSrkz
ymR3p+Jd9VMvTh1F1Yn2SkZyATrgC69EiZ6z12z8evj28zz4yakyew0IxiwAh3aUUkekSRRjHVbc
yDHRSjleWbLU7TCWRm4miTtevvOpz2pMi56YWCjETOmnnV4TUrAMAsL6vThMmMrCUuhr2BV4EOkz
BxWblacVI8D+7z/0wWO1uJMKP3mqX06QU2kdab+QKjL4xlVO3L/i6YI3XhRSYbycKJQJ6NQNdjFi
O10FmW7YxcRDEcZ6kOoxnW9OJtpP8QM79bAe+OCEUV1U4H82G6KACwSQZxnUzDdcgmlgjau22ADm
YQkAKsfo3tLG9FDx+4Hvv5JKLqmqQA/7ayv+7t5raRtCNEMtcqXrAFj+lrPyB4E1zD0KsVmb3Hn8
/EeBEFeOVTAaS7moKuXchYfhgw2nngxUdKGas7zqAFLZRnOl5vec0XSV1IKgxx27V/ZOkIjiNmvD
yq9y5njG2uIhKP5fQ7F0bCDrLe5E45+t6DiVcTzshr7m6CvQmOTLAjNKshpk1F+s0M6wy4EPga7E
nxpf39X0yWCqAnoq0h3nPBB7P5WDcWTyyK11uUfaw39QBGCrHdwK+jYreULRWHf6uDVjtCOxutuu
HT4iOKA3d8mBhUULyiMZjB34HeS5efrK0qkyhtQUjuj9JjnfzLqfUe0n8occHLm+t8mBNuFSab7C
56nVNX0MyMaIKcoySpJiCYsDwaDJWLlzd69PNXB4ZdnG67XvfNuXZAAvjP8BkWveORDBq6VCwJe9
yRtstR8Lo7UUd1hEqpisp0GonSzaSvDKTqDNOgG2pEwuD5qIrSxO2t0bbxB4yrwNZt2XqMoNL9Gr
BI9vvDquscaknhIRuVOB51AWuDhse+TUvPfYjMDbAguGRer+VxgjT4oBJzuRWCZx2u1GsHZAHHmI
Ij3+aXYarGDKsIVPqvk94sGhE6Uhtd22vaZHZIr8h1oAKFBTMc4ERmpMff8Li03zKzmLXo8rM3FW
iw5GZjhFn8K7SZKEj6kcNxqDlk6/CBPn1nr40V6uz489kvDFzlFgqJDTcV8D+pr5JfRNYsQd3lio
BLRY6cux/YonVkcjniJiTBaCM7pw+Lmys7WuiKJnAOScWvNypHjyAUDwwFkkpq7u7bfEKx5G9Hrd
1qRzgKN33iFYXUPO8dOgXj1b085+9YOKK03DGA5Mr4fnEnu4JC+ubFCmhKX0y09chWEEEgA2a/ED
VY4/QmO6R4Sq6P6FY8wrq5T/wzpjG/b90r95Vd1e+3b8uXekHQnQ2pA3mMbLpH3btnRf8+0O2iLF
/vCq/pzhza3xvfbDkqokTvaVHXL/kS935im7814O7oQxB/wmkaHxcgkQYKq64Cqd+wPkU+i4bqk7
DrnR3O9c9Q6CQ9vFIhgAxWoLeUolyx/Y43LKQyIRagO0kgqIuC/JnqtDptqRt7r/hiAH7Wx1ZOv7
EpQTHK1Y3XDertY5aU+IflvE/JjLY5A/1nrWY21qnLcHDG8bMRfh/9P0S88ObK9dHWjWMF12/nkY
dk6nJoBuqU4xoFS/njnIarG3l6IT0yXIwltzln3W6heGizrcn0zyjvC6b7umyy/tAOOh/y3yEPo+
KAg/LB579uXvw+8qB41oaK+SKiDXZZ0mHM/r559FJh2j7CuU2jc1ZeR9f9PIoQiFszaKkxIG5mrd
h+jdMmjPwUNWz78GwNdhmwdkL3ETypI7dM3qohuQq12Pm5OlYhOEe675ZByeKujy8ic+VwUGIk1Y
tpMNZWNhxV2hNNKx7lcXHSb4G7hnac7KyCkg+ZvfxFEX0svsIFwB64dHKbppf0XDPN04QuGSjkDy
IIZy4WQ1SGy6llVN27VdC0jlNmlOrDbcTwy6vS3BJYzzShKutGx+uw+GXHvUgsOlL46zU7B/Sr5v
73i8MXFXpqg7yTuMc/dMcx0r8Q0TF4HSzFDAzugtyAIZRgQTfgUHJLRB0eqjZdsWZj5U9bN1q3wG
j847Fi1FlLIKe3MKPGTsY2A6VLRoAEYQ0/DQRwhp8eHLGi2+UxOcC6pQZGchYYCMX4BU3plaoARo
yuj0hibHgEhBspf0VtL6XpDJaF6JuUXLZIhdocsyUeJGxkxXcVmN2/0perEFc/T1zJSOYB/IbcqH
/nzgCl2yCvLSu32U9Vz/W69WyK/+MfVGOllblDHowQr6TxZSPgkVpny2PkvKDcLGEx4VbKgcsBvl
13iuMWgYsXLUHKCJzotdr0AsKpN15mCEMu9tW0lwP9y9q8UUmIH/QZCS4Zt/TdmRxedgef5YftA/
2NkBedmPC5UdUbv9aw1A31v7s/Hqto16uM0WsioSsbhrkl+D2MfQB/EbR/z5EM+eixTrSTZbXtWd
d0nitIW1mluJsTm/q6uKACc7CVrZHo10+nkB9C2sCnW4huaY6owuYo7mRX6FiuF82KiTfKIkwdwV
Det9/nPeeGWVinrW5PJowA0n+6A641aCR9ywiYYBtdkqL0YgxZQ/OWItnjfX2g4rd5ogoW8JM/0i
LL76G3cMd4clC6pruXHNclmKf2okDaWM6yvL9OKL9R1botbUPmmjQWjXotaymiUr2A2vIXmfPIXT
l15oFtzwWfo1Y6j7RXuiSUAzM8iNSZ0PDLUZ/l8P9HTuPHd8YpbHSOIGhP820JyXIwpKr4ckxFcg
7J6H0KqP10L4BdfNAoHJurErV7TJT3/WlCzpJPqIDefWMmB1CvMtWHUj1r3jQ9LNJ3+2gykkyQit
ib47j0v+SVGcrmn1Z2+iOMFz+FfmEo/jqpCJXJLareGTOKrLmvmdXU4v39dPdXkd/hYp1wD6STsS
a6FM4EFbKRBeICVo+B8ei0C//CadLoZNDR8gpfHvgIlY9lNtERCb/c+tjInxBXG6pXXO3Ej4YK0J
+BjqPUWWpU0h6jcDIrnsPFM6KjQf4RTjv2p/FmJLSU9c/Z+9yYJg6Ovxo5qkNHgQ0J/2hUdXL4sl
T9xT1bi6Jbwd9PSVWNytsDue7ON/3OruRxPWjKIK137VjFWKHyFimOO32IZPmQvSFgeyQy8KFyQT
RXDz060qZDYRcYk5j0FZeF53Gcyz5rZamZxj9ynhHA0hDM/aZRWo4JVR3SDWB+qPVYHKRZ67kjmD
N02LVXh/RUpP38BmEU1wzVPTHGbIj8aFwc06B60Uqa5EC/zbiLUWnVdmvS+tFefqaRViFPmpF9lo
wZP9MQAfyXXNtRiHHE9D+5hA8h/OjT+uJjEqNJ3buaTk07s7JWHcg5VV9RqtK9Y5SpPjmSD6Q7uj
/qcmhOJqZooUBo/OfS/KTsZQiXErvb4F2x3+w+8DA+hK4yofN6Tsfqnnobz47j8wrEdc+PFeLLjn
3I9y2KB/IMBGnfq8VmIT+ewsorxurLspFBhasxAaCN3lJ7XcCAEI5eZvD/pHiL2umDAhLWVa0dM4
M2JA/05wJI/NXH3mp77RaS4FoBb2J9wdG8b/Ziq7U7hU+e0NXpLTsfxJgmZTktTokXIQZ4jl25oO
tFHoxM6ZEMyk7llvi2AFgrHQvir+Q+udd7t5pa1m5+9Lt/iuO+ZgJ+A+4gr+qW8xSQY1EEoEpASd
8q8OHvtSxE6LohPGB3E4HW9H0g10RKz9MEayYzuYqn5GlQdu9ACxbr3Nq5Jgi9JDvAqQZGKgxevc
pNkIJWaBaIP2mRdYEGrNpMe5XXYfPQFrV/sdVZmQQfkXHrELJ/LbO8CdvLwkbMOdwTfpOAvvRNbu
i1SoF6srgt7OgN0FGAw3bQoZnQUz6C9GltdgfGfyx1Gv9VJDrz/LuRnlu3TPXqyrSzi+/pDD8ZGo
vAR+N+MQdaxatDnPW/CLHsVUECA8DPmhwCEx0n1+tAJ2YRvF+aUf7SczrhIVOS6AYPiA41R88t/0
J3fgVWB65J3bE0w4YYiHMaNRg2OBH/cTUJtEOuxHi2Qd4emgc80NYcylwSlbhSlucA3+CNeMyAdK
rw1+xLAeTwcfp4IM96xC6JVUEBrhC3hOBYaWlUIQm71wKyLZQcIuoNGvE0lKLERwsx5IwijOXU9S
4yXQE2nh34XRjK1ygP8jp01k6hPqP2T8C0mF2yHsIhzbNJDK642eopCKlT48oxDC4INo9UsBD5bq
FkyfoR2wfojy6xU36m0tPZlDEzQaFjvVa5ebPvnws1TD4vy1KyG0wZbL1gkjdXPKCndvK9oaXxOC
JZYXjfhjG52g0Z+OUS4jlyDpGYcVLzh+gONyNEYj+h8AkGOkO4wuPCVpkHzoTqyei+1a4GRtpfAJ
5KHpwjW4UXFsik1PoNJS30SCAt25VChf/7DQGPtAfSroPGaaNRBbIcGtws6zUOzxUMyeWkxM0AnM
ZX4fAOHmYPHqjNHn3QRTohBieogyFVYlM6pxqb+kg5zRZqm5unhaAvXAGWhL1t93tF9T9AzOD75y
mX1BkqT5SLafCNts55RdbQkFHD9OSLMnxT/fjp69XQwoKkKzxzLbJO1RC4q4L3HD6z3GtDmo0Gbe
KJrEujk0/5rtgWPBGKpx2jV96TDo2awyG1i5mIkX/b9mTvwaFCcmVwEqM3uubrAIz8Iq+9eRhwtH
ofUHl6mcpaeXe1JsaKc+cdPmdV8Qid063aCAITg7l99z6OcM35cvTQjCJ7UGo9t7xmLjpXGAlysH
MgYmw/Ekzv3LtseT3n+xrRofP27Eo6SDhHRrcDBLPXmO2wvCIqcp1q/REzrxT6S9A8Xqwh0M8491
6njUbO+B+zWV4HgPZU0WUjqxjozhowF3YrWN3LuVubCDYWsni4gG3l6WtL4DGsNviyFiY2NQb8Qk
/4HkRCv34Khq3Au5XXGjw/xJAJx6NJkwDk3SNAJLTYOOTIdt4x5IPvMyRGTU2pot/imLWpnx/l7T
TUwB/GPV1bGYKdeuluG6kz0rNvEgspd7H3doUNFP3Bpbt3XFR0b8mEP3WrBaSyfxomEj+6qW4Pb8
+13FuCFvbm+YYaQs5cpVItzwmKEBbzFgHxigL5yvKNx+91TiL19o0o2mQ161doTDyYK/4J8FSZge
QN8EHpRwCWKbhkqOlh1UN715+6eAaX854dZ6vWzEZjUBQzhLj63YUiGUiZZ/Sp1G8fqfm2b3llmO
qIttTU4tKsMGBzDJDZv5dLczFpHineSGsMtTtd2W7BJfzn6c/Xpb5DQUpWpTaW6oki51l8Bqr9Dh
yRcyVA4X22CLF2Za2OJZCgZBNaeo6Ao75HI6u8jCAISjy0kakkbFV08xOPJFxF7+4vqrLCk0aVaw
4FFZnS/sCCp7CZgq5V+VCFVKX9svumGloZe54x6zbCFe96qWH75yhsr7B4WaM3ce50FRl7kF1Dmt
8OvYv4J3Zi3ndVYPE4bpFcf8v9sdyTPJjz1KyG0s14pM6LOBYjs2cM8ShTryIXyTfY78c+KBWPWz
eSHARmARlPJ6Dy7ery+0sBiyHKZZ/x5wsOi3WOBnr31NuY2SBGSR/8JMut6WzPDrTspNjxHW9xXY
AfVgLxCxUwv6T3/EuiikrdUwzPBnkZ2Njpu6FOFFK/g8h+pK8U5CRZODFri06tt+qosPdhhiQ60a
Hd19KoGFNrgUBEHlKyOKxdwHmTzzxdKJMV56xWQhaRZRaKKaiZTD6LcZvsjair851bjj4tx2wH8t
yYDHPZEJE91DJoriuZru0nSWo6L8acT9imlEAlZBU81r3JH+bUgT6MSqyKjexCksrXrjq2/l2QL8
jdIdHFlH9PLOpyWGjbvuito9NzmdZdk5EVmOFCfPRcXwCYIaf7dw4g8wHAxSSYH/V+B/jXnx//AV
RaoTppIP0Yo3kz7vxbiSNBWbraWGlfVQkwRDOicLwxf+S9IHKVcJhi8ABbqI+68zNCtw3UwQGbMU
I8etA3Afhnl8sf03KAmVPZUzVdSzS/sLQT4qV6LUlJHkVbr95Frz1VfApT5fX6zPfvWCyysGNyw/
v41Yugn8wkjzi6bybawqLHDoaNlunFYRQSORaWTvOtFfwSOln6P7T5Elur2Pc/osdsUFaDikOfBS
TibjoA+i5ynmmGwEcPLf1Et7u0Y7JvjOm5/toR1DiQkfT4NhkG8A8uGlpynzEfkrSfMBiAjCVBMU
uqL4m/BtQjA6IdwR+xW7pd02Rk0xM/el97Wl/3BF1WnUcndvSEVJd9TRyKCgh+LuFsmWVvHycJYy
VpN6pI/BPHjT7ccS0BfM8Eq4VNHTPyqphXJWaACd5QGsbxMnyWemO4gj5qYQEo8TuWINE7brs0MQ
4JAOE5y7ivNTjRqJG22pwubBNjQ2i7r5i+39gaz1Sww4Sl7CIQQPicoPuqPvBDp6T1lREZfAmwEW
iApiIL4S+ic5XvfNJ/J5EcHNYPuo/XVtKauTDR8luf6GGx5qxuYH1g0LluFZTB/F1iZJcmXnSJLd
SgYnKPqygWqrxLj4mM1l3yqK/YpDHNA75d1gUxDt4gRwmN73FbJG7gAQdhWT1w8t7Ri83QOqut0C
laD/vpGX88RB6junWyINyJRM9K+Y1rCKmRQ7wUjlTbgocdStpp3ysL69GYmDh6l72rncadr9hQlY
3EkRqHzycFeBt2oi1pqcyz9UgUtjojUh7TNu02G6WoGvzZ9TKhL4eMAYBbSYzrhceRa70ozAPYdN
u5D5lrKnNg8fdxgXld/StCeFePhqvtQtHqtOmTT5a4CqKNtABpRgPeKOK0z/Q8poDM6W2z2R9eyj
y5yrg/p3sE9CVzHkN56wqmKU2dY82eT4hawOhRZRlJhTbw7RjErbzwM1yTpqaacmGjuk9PaLLFd7
hB7M1SiEaclJbh4XmCTFKnzd8vMTUs/JTB8nEwFFxUeQjDPhE9w14lijSk/Ly68wrLbFLMtNjnWC
VsGtcdtpxUddbToR4YPRGScgn6CfcS73IFB7uflamhayD4O3worQXLClKOuuZLwIDI0IDpkc/tty
dO1SLhHmYf56aQ4wh0cJb0Xt04P/twBOby+lvS5Oa9H+lea2uNYHRkutujHkKO1F8V6SJHCPPhyc
Au6hLspH6mGBM916OrZEZLaghzpgwwlZbSmT1I2/QEjsiNZH1f0Y269KG/giWBdvKDazFjsFsYcZ
zKFsiR4WDutqbj4S+xQSrW/UAfThGNGTubm+CpfQLNLNamK5FpDeWiVfauJz9E67+xjr6u06Ycks
cRYwyp3EhzdP2PqsH+Pp5hAF3izSNpryfgUga1iBMfGN15H+oI7qoP0UUBbnbNzx5vn5zpjUet+F
hf5XZmGsDCEDjRYO8u90AnUwYfmkXL8/bOZyUqA1r9nFiZNLM4zJ6/vx5H7i5QC1MFxuvvIPasxK
Z63Tv6L+V7WWGTdvqUeQC9mL43CtYkytnxhF3JioCbJuzkb9oiFbcOyzEBqiFOHNvsnuz6b88fLQ
2epsXu6rqugC2ACS4drcD6EvWKTi4bNsboE4I3UaGQf9QnG+zP3ovfIKyvQtqaJ0yV55VU7rOjUR
KgpGZvZAQEzlxESokIeopU8C2m8JJ6Ev62HZprsJ7Ew+RkixQnG667Zi0z/K/JfFDR/GyJEiIDgn
HhMateZjuIRwfmZMi/6gIkNQ6WNJnA5/jaZ+RPlOK8I9IAzspXui8mnGTMGsAunbnll5wCo2fXjh
ktXnuTjOMrKh6au1I+CpYwROFwSmYKBD3/ETRm5v9R++/AdCaqt9N9cgYSiD40AMqF/wMQednDxd
8FD5iHQ1tBq6JUgEBwnRXmOn9Enacj/Fp4dhxk8S0KDVvSr/1iRX8l6b263YrOrwZe9ENvjU/kse
XUXes1Udp/C3NPktcqlpGcja3+dTdrLkvnoht7UPYY1ZHoKebIZwRGCAMHFHwZSeFkDJhCNOgrzj
tDJx7mlsm/8cRlp6H++FSY/W4Um+qMIQeO6LM2zS8TRZDDcKoPxlPKXqTmc7NBLCO8HIwnNrEdaq
YKG9dwh02NkZMK4GZxous0M/7jDf0HPnFpjBZ2SL/A543aOW1AtGHtc1wCTpDMZ7xtzFH9V7gZzf
PZIWvDX5gmf7ziP0bycDnoy2t8ThhGvjdKU6jaFiUvBSGxhUi5aeNC4ovrtpa0huKBhHRwH8LFul
fgYBvC7gEUpXzuQU8eBhEBWGiJtgum/QR0PR3h4VihhEE9Z+BXu6uxc6kmJM/3jUKoc+pY1SjFi1
M3UF1A02Qcy+vJ3RKiAeU36jreC8WftpEaaERH+vNEcNAdfwWXkGzlWnyHHZAGyDH2n/tRrJaPnr
t1PeYDaSn90PLuWgPk2TClhcsF8A7s6iQw0ogk8sC+tN7wzDc/4oKHVWrankFxwlEVaKjJjgcqcg
neOQd8VWBTSwlEvTkvMneW5VaMKZCnNJ5uEGNyF8/AlEmImLkyEmBkAXWlW5/uwPshJb8Bh0PdgL
EG5DBORvCtAC6ofRfM7SKdGy0IPCQHS3xR0EQfMnIkQS+/LFqjPEw46Bij3hcTw2gWYRBNvcYPKj
Igg6ovcs4P6kQragkjDNOiN2/mxyvKnxtyWY0Uyg4KOSqppCxS2fpmmGU3IFAAA8WvcdfJThMUwR
PVJKxlFuWWM1lParTTO0ZUqVCeTKkAaBXGupcf/y97CdARbnQGY45vVFopSQ/I0cISSIemph7tyw
J9faQUxaq+cGyPKEb4JfXdJ5a/O6Gf5V3caGyITJ88se13AjtabJRqURa6QY4cAeNsm6rAxF7n/Q
i8OBPazVjrx9mDYKpA3k1y7VrtF7CEi5eguQcpICsUJH/OQhRzv8D0MoTFPRE1ehpYFY3aptg7DF
T8O9kYGfMH/XszhCxJykhYJ5xwonDKq+Mnl6ErrK3bWZDKo1gWMouZCB/NaBDU8ekfjZrqH/Av20
SlLUvmYqgmO25uErT48EmPkhOgf/+JhZX+XhPZzV60m7y6hGw62Dr7wcSzgvXUCHSLdwaPBb3zVI
EwpZK+xydKvwJed+Ga1kuixSWjUkgWVP4M+uWViXS17e2wObQ/kWrjf9ZqYGcsJGoSUEZ77bVOhv
uz3GQK320A4aL1vrOaeSgsbDB9MBz8rk6AyJ8QzCh+akx16dZb3FQAaWqWqjuoCN6QgSeyf1K9xZ
PckR/U4QK2vj+kWk9IsUM4XvYhE4dFxbJvyxueXuBWKSDfoDj5/GAAnL4UtmHLmjby2JUsGpEvQ5
RwkVLwZqEg9SbcpodSAz50WQL+d/MdK3Bs6ASmcTlZ1pZlT1MbvZ/AC+HedtbAn341u0VN32re64
V8b5ABLtlgdu9eQV/sXqNN1gi1enviH4jUdXt86T6WH6OCAcgjzrzfN2V8uRjT67YFarSX/ZzMCj
kHrvTvhPvIKri3LIIG3eeqVHc4DcVvEbNoftfhlHV14+VAbYUABAP4EAeVaKwLj0DMCuSUagAm3I
hYgPVUQai4h5mhv7HefdG9OimcuyK5JE5kr/KblHzYuX2Xa5QxcvzBALcxlR90ws19aTcZGKDcFG
8EdReHY7tQCpeZwsTLuOiazI26zuNWzcQS1zsVeiLMfLNgOxhNTXVjTCndDOP4KOcJ2Vi9+kLUCU
NT9P8WaxkWOaszRbGXv+tys51LgpZYqxUNKXps3QhH402e3z4Cc0Gfv7KDyd7Fp8kofQv08BD7MV
elbC3N71Ep5YARC/1K/BWOaJIxDtKt2B4lDRGZ0NBpQeqj5ljwTyZe6phpLoNRYygz8kMVQmJnyW
JgcQaLaeiKFzgxxhTprop4kP8PMvCPA5a1XriteMiUa0Fr3WFNf779V+SgPnEsSVTashoJTkql6E
gRkMBw8Rkn9WGD35vMd/4yWynfnzugk8wkOXR+zFvm02ykJxmLlwKcXm2UsKUkZDCfISdXW4aKPD
p6M5+6/4BspEKbuPB06gkNdaIj76WIECZuJtmxMC0g7+Cq528AFPgsUHq/0OUAKODDmtEC/02xKW
p1e6P6xyTSQbwk3rrOFZsPrThbBVZ3+DzQLrdBtQMLcZHnGehZeLepz0diJ//X0QZpAp3Gd0KjQB
59pIgoFaOfp2d7WAS94JRnODieZyFOGD0kkl6uUbnoq4oXY8bb/jH76Ceac+3tg0qyedJn6Ed6as
6CCwygE45A1L2UFcrlQjGshUYaMcvxemzH0nMERwD4G+mAo+1Z1jbTR30Qg0uqLael5PVNSlmqdR
eq3osVyWFzfiABRc3dU5W63rs9B/V8GxqGEukd/tlLi+N+5Cv16iYgwFA+SztvwcQ3/j/Q9m/R03
0e2L7bSJGyZPdlcU6FjHFGZn4hrpN0IsugU2lRKh0Jxty1Wt9PYCOrTMILhKhoWPN8Cc8lyB18IM
C+4Rwxdo4Er+e/aBZPlmhgMTfwYRn9Q6vN/i9LvkBnZjlvGpNvag4HUIL1Ve1cHVi9URM+/t09rZ
BPXsbyka+FoQh8yoGTO6J/srsOff5b+m5piohewE0xHn/USgTPbfrrm309NYS6Ztl3foMi+6FtTi
WVNQGkTAlxiQu0YZwfB3Fza//CUYpO0tQLNg6Z2Zkn71q9H2k1uh9XTuO+xk+BGw7jYLolhXjqk7
gxGoOfdqig6DdMvXNEe/RuNBPk1h7Z/ptB3wH7wTdLzezBQ0G/q1z2jlqKnMkg49NB6CyNiH9jZ4
/arA2I4EhI5SqDBk8ka3mPbgsGHxTDYV0IV3nmPoFYpM1ugw1ve1ica2UJ83l5vniT1HGfVEVDmI
2QYYZQwg3exkneVFq/eskY27RwFLsu/oBy1xnYA5bFdhuyHbxp82ayOa43VELJv5ddHbHSB60dF7
v6W2lDAKar7VsnnI+dfIdRp+wHy5dMzg51DHsZ1jML5qAc9cQ7Hp/KZNCrzw4AbAyLgS+4V9AO0P
w+s1fqHaI9cCuS7RluzGQ1kDEULKBnJPox84hsljby5l3An/GeijuQJ3tRIy8iXQwqM8W5VN4Q7k
mZyjZcF36eweXT8a79cdgP0Lib2cfljPqiph5FzeMoQ97sxjHaWIRiPSXY/JcIueLzv1/nwZ+Y73
wvKCbtCuy7Ev6hwi9jP9TKD1usaBFbH9qo5eX2YRxyK7LUxNcRUuVXuIL+ecyY8hw0UIrPpJVvTY
2omHfYrb44YgDfrESqqWLugzw67e0z8r/1vmql5SIDO55bU406UJWa7zC/+PAd6HgkQ77Q4r3Ykp
sjsD6hMbMoaEIXYtZ1lowaEAC7GhsyAuzJI2Qr4eJHXa00QWv9986YwGNr5p2Uh04ls2s4FV+gG7
ByJHT3WkTSUrFkaxvdd5IO+57wUcvX3HNMb8j7EbNyfTSW1f5WKJjYMXA/9iwOcjNmhXJdePTP3L
1G2EvMuByhz/Zw9E6Mhjicj15YQoPb9bGcUVKbcjTlg8CbucX28xciA8LPkI/aM4AUx0deXrBJZA
cWNcOfJNXfGuRtUxzUXp/KR/jRQPCn5bcdBDPf2/eKl1lZxz865koib+4mUDm904VsoMSIaH2b0w
pj5JqetV66xJiR2AAXpSbPHgRotcV3WW81K6OyRWPe5F2vPMdQsCGbDnRMeR3urPkvbqK380Gpfz
YTArKN4LrkiS/UBmWTm3Ydi/YYljt1cAcrTq7TmlQU88j3feEFG0qJP1qjU7DWcwGH0BgbWAt4UP
AHTqjc18yWqAmB8dy4H2paYfBhCIFGIIaWTTztTqV3sM9kFR62VFjgYRA1DAWrFz+Zsj5kjPjDt7
ElU78/tWd+hZVbwbke93PDVtNXq1nQZdT8yCkEYZOIbmeAV4RPFmCFDcR8AQ+b1qG8VPLVi8srJd
dcjV+EoJd4AGskmegANuG1sOP+YyhmtwwEH7mZ0AFMw15hVrPT3savEi8R84rFNbaTo8rENisSYU
KG+x+y/SocSRqdyBaD7+2Gv+UINDYlvzanwUuxBrNpsVina2pNZpPVK6+rRkpyazu6TGRzsO+0y4
S77A1n8N+QJ0iBBDB+gTQKSJnCKSxbcd/BhB6wRXPHn/KWJWCbcz0kksoSsaDPCQrmOpw/9ZRV/5
wFPSAOJDbkys0wVRji1krn+J+plVnG9JWlHqu6CABxNQg3gxcFcbYq+7uP0kUCoYItNIPUm8vNqb
P6A3TVAzzOqqck2BD48xOTL3zNw7pvELXVWUc2O4sUmy0BKfTECfmaRoXPXghfIouS4c50RhWbX0
eCuHacN3Y5CKnyv08cYY1oIHopBfuhz92GzINfmrtpSIwXzrxTXofiDI+h7+2g0EoX3Kj3WVeaRy
s4W70z+ao49SsrpN6L5TT4/gpbiQHU2NCT0cWEfs8Tk9UOxqj6nDQ0oVj+HY5J/hOvymmoT7SxLd
aSIGoxHOvA4IARq8pPe9rJFSi9NwbGrLIfuV9SZQMKG2Tnd8bmxzmooSUNfI3ww5HQjxATLRl6wQ
zTJmnmNZe5dUgovfFxr6pGQpY9umJqZqXNzI+fgEfpHd76txEFbzXVj4icG+iMS0NFB0+iAntw5X
TJIwpMiEc5XqqNm0sA0jGc5AuHvoiG20auXQ/AhOcwTX6pi+rBj3YXpVtSb3Yb4S1hQPGscQbv5L
T304tPbYD4bLCuPxP51IRarkpx28MAZndM7g8z2sX4u3PPERKIxUtVEypH9U9KksnTtBuxqlKO3W
BAJDcr05WdCl72DClCSOytAOPjX3UAMgdMKWtZ1+sRl7qy/irQRTNtcTVahn5Wcewy382McN3kH4
jvvqy7e3pdNpJrJ818PBu3jkYTrk68lNWMpVkYTk20V/GYvjN/9mCA1xF2iklHt+GYnbci0T8Sex
kxfb1DicPkAXe15sLvsjNe7OwmJN9YVon6DMZUEo3djLlZYqa1kgJDOGjqQBBo+vj3ElYIkdcz89
Rs0ATI1Uxmf3xAvxBjcyUeXUtY6PzxpuCBW1bsrwbziDMt/sLINuxiC0emgdy9anbFjD3nqYbMtD
X0eVDkd3sZvy43qDucLGnHUrmUTLKQPH00BFWviF7Ioj+2IktZai31mJcUlbiWqqbLPdwfxOJlE4
HFa4ybrbL+pB+52dHnqRjqW4+zqG8reAVvD8P/HsYeLHfm9VO7rAUDIto7ELeYycRN2K2Dfix+2i
xm6enoviMoZtf63wcX0b/WxPkHfx02aCYyTm5PXf0IJ/y8vg/Bk4nWxtDfLieKj6JBnUWtpSJ+N1
IqEhzMvgRd4dib3lDcaAPr/+Tyn3M71Tl0KxDK6c7ZGDaJ0fRJ8L1fyihtK4fkT5uIkRoPcdHfSI
QoQVWbuyQkE1G+Zx9nmAUir5QFfptOl9yOdGhLvGAZh7uRDl73fwb2aoBkaumStfPfDfMqnxutwV
9oihpZL8Xqt9OxAijn974XrequIpQ1oEHk3dTp9XA7tisgU7jsOY8TvkRyaRbjXmfLBAqs17PGtQ
2OaCSe+MpjBAPINym7XThB8E4yKroNS0sKOkrQI6jfFenDsVctHQsvBrw5wAkmZ1V5XLoKsEoMv7
gAkyKXwc9KxaMOzlwmF1hGvCFZExSkRFziear/LfcmFiFdm3OyGAueLEYTOylytfJ97yey0qDPYO
gTBhWTlRGOAWCO1EiIrC9J+htSD06RjF0q+eDA+SUkD73Pa9rTJZet+ChrjCoF4/aPRyNW3KFDlV
3vxP1ZpvSBpNOfIagTghw1cTk3tODmobJvg8JROogWciMgZkgfkZtuMOUzE0vkvkNE4iunUlrJcl
zJFXPikbuQwUAZt75r3+nwtpOcdkzQexmD+D7rM/xc7tYvIdVxsh/ZF+r5mTUu0Swm2IIuLaAxDb
zGgKTnEhH5cbWvKQFld9OnZCLjEj7t0TInUUHjP/f4fWGMe/RTBeNVje4oBErmMn25/FCO/lLqkf
ZYPzBXKJYQavDUKOpSONsHePo0V8BSLMBLffWbyxA580jX+aDfoBwfSx+1TFYz4UThX6ulh7nWg+
pReiUlCkEDDVOUqW6Ks2wjNueQ7zObFYrpqPzUYZOkOZc/OS+okO78O5X4rhyTi0naykLIwm0S6p
szpqjqYonQ3bh/747WpFp4RN4GrTNXuN3QfJsb0R2bfEcZOGAfW/XOYc0G0Jrsqm3bcDWaY0JyDp
r1FYphpU7kNNqry5KTl5HLPmDkzfVDOZjRd5AVpsdFq3De+Q5tT7TeFxD92OLJl7pVYwzo1+sSoP
OYc+iII74pWaJ0c33nuQPPVR87TBkcf/q/F9Af5mEZbm9MFi0nPc5Ln7caT+S0hjE+YYRo4VIy5k
wvtONCV23m7cJRQ5DNkl4r+sbY+o2Qm78vUhYpi2CSFPVumDTf1LwwCKo6hf0YrXLJ+kIeAbzyFv
1WFeiZiawYq+DI0KpCssw1odaePOQVGMYpyalt5YXOrg18MKKkKtvczdD6sT/mGAK87QxR/bPJ26
xgi4lJO2zmWFGYdVRFUxwLTTNkMs79fzTIwqZ3eCvdSj3TEG7p5FjedmR2yg99suCD4NMb3Jn8n2
ekf4ZtSB2w1CPj5XUy/hr7xVpBvjqe0APH70vlPfSRLwzqqD6Yv68FAaEBfiinaB95qVlaqvv/3K
9JJyjr3KLutMFnkfVe+CYC6CknGW0ExMSu1NEDDTJvOKmI7Epa5WIZ5gkbNvsk+68U//Pc07w8Im
Z2tlsHN1WlUqnFFswiRsbwKWc7cTUaVeVaWm7Di61lCyNvKUeCM+ub8tT5KKyvBPu4hz2X+VEqh6
RLfLi8FD/sgtX3L5REqngMvFE25Q2NeC1ShUEM6z24Fvu6zugFz8qT8vvq/HKA/y68X0b+lF4fm2
4ZdPZryg+iTlwvXgXDAT8xv51F2FD8UZiz8uDiAp36LzMeJRpgvc+jyKaEBsuH4k3Zwp0L8GD/Q4
4/g6b+WRKniEGC/06PDWuTNY2vvZcA8If5BPY535zqkFWvVVJMwL0yBI8htW/zbwdCaK6VhCQpl1
BjgyCJUUKfHZsQ1UHQ5PRScGvE8+eiBuMatxGG/fblUBUavn1SASuKRSBsQosnwzrGrxpnVI3eYD
LwCvyuD6CvAwof5gsK+gVddERBo5UVDR9H4RDQPCx//ZQZQUOFjM5VYmNqyhOWDVqoK9XFUSmPh6
DjnLvB3ZBz4i0T5gEkpr3gsllvzsBKGO+iKRPx3VAZRdA0r6NRKF14jYgTisc6DJjUyhbFcO2Pgj
p1HUmBxxlZb1s18xXMMxwj2x3TRSxlGmLdW2dcxGgm8yqwJIeSgDhuPbDXB9nxuHoIyH2NMOKa83
8+F1ZJAUnzY1evKJRYzUQYIPtcjxb3ILKIqTn8GHG3bhWBORUAA8m1i7hJN+0y8bUSUhdqSmG/jw
jSukvwTBcWwNGXatwl/tDCCMQ56gDSsHuky8KTf2J7GYm6q7Cjdxk5RuYM0S3xV7Hg0QCSoclQja
etvfSeVc3wEqiQMBSnoJ/lpCKVl6tWodsa37zTUZuqxzChqZvi7V4HHnWrDsVLipQM1Cn0kVi17g
2PaZCpAc2UgtJKFuuWIuOApgoG1fyVbNQx3yz7MOvhHn+c9624YbBHqWz0iOLswdPqHmw88ck0Xp
fWyorAqUB0STwQpkcrKKOWkTvqAoqi29Ixlfee1JoJBxKVft55LMqIMEBLshdGJFTBZrIbQSaJ3K
Cf1a6fw9U54LpUoSdxAJFh/qMAahK1LfyWMq1iXqIuz4Aav/n3Sbx8qtpOIoGwQip8CcVPwF+9xA
8SFlZBPqV68Dfft1bdkssLKkB7D4OnHmGi25rwP9YfYyKOM2l2qwQRQj8OLSgb+26Yprxow+mgNm
80dvkjj7wpOr5BTh5VcF1E0y3vOQFcwIbFEbK+XCp1hF7JpH/2LDz4os7nb4CVtzuNaCS/oXvKoq
H/ZyESBzS8nUXLHxYeeUryVw/QOOTBipevBZpR756ybOqqT3+xdHVYpVhkYVo9FrzpercYXO3tiu
j0vSM4xuVWyxXQZyZ6+jDQTAIMHMwN3vjiAnOb7weClip/QBR4gZQxiK9Cp4JSgk5l45jo9zDVfB
VDNHA7BmameQ7DHoEVAp+xjys21nqqqjMGp8sn/q1dmFksRR0jhWoXUvLj9xEAzRaArUvAvOSseP
hLLBaiqeK5/be4JzW0oP8N5WKLCQ2sTTmV6DqLfAXEW9qOKgXaVRApxxf+CL+XOAy4zg7nVBLgjc
nntkBhEb3PUpWpbrOoBLHqvnS1b2VSi6Yxx1fZHdZDPYhYntgNgp/083+qHXysU/KpyGSXahNV9j
+uUcX8TRGPBc213M0TDyHuxX8fIwWFEfaH+i2FsngsUAJeRrMngoBE3v9IGeZ058jFZVxTzwuze7
lk/NUcoQVAFIjJSMkd0ZtENMTLUdOOHLMKiTzyrt6U1v3pHQTBTO44RQ5MOcslSc7sHJ2nf8LGUD
/Uw04w79NVROSBWpwk0MHxVBTAqUiHyzwwdC6eXTpgdH4e4BbmeN98r51eCfNf82WjuQ3B6S5Em+
/SFDdOc+KwieNmRsjUIMuUKudtfj8k2S//zN1BiedC/pzrla+9Qx/CswwSiqCpuanbDtBNCd7Kws
xcra48zKXNbg1aE21v8JKs/q4QT+qCaUcbD+LsZ5rlauz45QQKOnvHTLWin6XR3jv24MS+YRvRA3
EgmYygHZDdYIoxLTUB/N/wA9IyqH+WH9fhARDfCSTe/mH7SBLbYTOwTJtXVC7N3tDPsG854MGckj
15f+m5hz4YJrvVEqIXonlV2E5eG8J6cR8cT43Az6/vePt2Eq1ZZZFlGxAltJVOmYizQQ8cz9STlE
nRVZJZDaXC9H+a0ccB+RDH4jzIIbu11ic+BW8K7uzk8K7nRLnhEAtBG1ZOXk0XOA4jWWdWDJveSl
Eo271uo0Myhrr4ltkS3xRyiDuWETORE6XMglPBoICnTuM3MdnSroxeHC/S6mErmhvkuDGgxXKqEi
ftqMrbbjFmBfrrWG0DbAAFgrdn2ANj7nCwpA8kA6gGBNEyVjanzu4dwx5ZpRgD3b6FUn3nX7rQpf
mD4cg7ovbRqU1ijKTGbZi68FeqnqeGQh6dUlNDsHru8KrqZ0Qy23c5TxDyMAxtw1+RABk2bveVax
DXqSnrzTJL1QyZyRETk92OrP8WqXg4PMgsZRoL7XCJz4V2EZjJmC6Eqgk4FgUIcYwjtaT4Qvhi08
IXRtjIqSoI44YhMieqwADJcJM5zxPIS/DV1496AkSpTlu6utKqo0ILyDieQ+1pmUvA6rwWxoc8gR
ftPlntYw5dUHjgVVIcMhYtE5ZMZoJiL/Lqu4p+TiLdkXn0eJAv9N+33wpg1WYGRc/m1rrl0v2vuV
wfRpDeXPRXHahS9+6tdX+wWHARxm72x3y6k5YkI+AKsPf14+pEG1C5pFIoAKL1mu9UHrhQKoZeQK
LOBgX7s7kYIzCvtt8caTiVJqR+Ibmkp8QApHgIRqYfRMg3NOK+rcgVST+T8a7JraT9LZkmPiNT0r
bGTULFPk6RVKxbJCK+ToaM3Ht2uEHw9se3WQgFbSvO0v1wkgJCwYJ+tZCb8m8oGRmxRzB4uFDo7l
2+QFotigtwaqptRJbaHIqYWl8bYGBuWKd7rA3sMNrIJ1YNiSpbn7As6s5nP6lLgOFXmtJyJUP18i
NwFu3W7F8oDcjkLQ9OGGzcKD5m5VItkJ7SsagGeuR4UZR6gPPeSA2SzHsvULl6k/dtwVyIho9g7R
wOfEQJ2rLEtzuI7cG1fV1ZpvuTbR6mlsF7vXg5rl9jx7HZVsSj/GeDBw7sieQjfF91rHZ976J1hQ
zqbUeIR6su0szo/sCNogMP9VcHf8LYaXr7bZx9+xkpiFKvIJ4m3XwSJAkI4w3MgMrmKeJVhKI6vc
LfM5ilZtmPmnKyw50kc2FXoSHDAx1Z6Xlv9UbKvQ6eUaQjFG74Hci26aV7PNcNVdOeBBQYX2JDMo
843WNUTpdWgmJaYdtpn1OZe77R+5FAqQah7kK/3RKj07+yzMcRVKjwJp9ZuSLPRJ6uQPfx5t6Nzo
gI3btqjtmYdCQQI4a7APn+E5t/zyuWrHd/s54r7tUQqyeJIAZEoil3ONUxd7LmKW1kvjCHqlhz3k
G7W2Qo2VC5lHG3s8qFjfPMwunknWKlokomO5ofq3iuMhOI+u4JmtVItyvpyWvEpQT3UKdFbW82BP
AF5SqNvn7/5MJSHi7apAz+tr4Cwy9IJ2rlDPurKoXJbW+VKPUqZzsoju1hIGv0rjcl9Hr7I510vm
+w2+jnYsuOHZB0WjDZqluQpAbnHpaIzOUk7mjG2WM3MhJiPAP6bLw1NUHeTNCx1qJz90iJUstVV9
vqroa18Bu7sgpEufspnSa6sgTo3lVR1n5mUx5lKgkVlvgllADMI0pnRd5lwoFlBdZ77dPPXYwIwd
h7uQDbBx59fpPVVrKYyVG2LY/1iY4XvTRSQaJoza+jAZ1HhDU+Rm+ZpGxj4lG6JmwswEH6wGpvsQ
6iauHijvoP+tO4VPZF1cmEZbp4IPFGA8EKVEU/0XJnUdZ/qbuBGQg9nDcGchYzTZw6zNNDy9icZw
FUSZ6a+jnA2s6IfcxJoDNfhqDCsiaHoX16WJ0XktD1BsVyfUnvTn54gt4JslsQdoXgPXI19Hdxho
xLzNJhoM1QYorPjWzHK9yqWs5hUiCXI/fkDivRKms3jXX5+RO+gDFO9ylEatBjlQdGGsdriFTnbs
cs+qhwTdN8WkpWg4TA58nBFh6ESP5UOj57gdEeCtLOcJbV9Vn0WepxCC0hqGMn1nvzHkve8TFYw6
5vB4+ddhSlbCnFWyBQbUis2eKTLs1cUJZhgcYjlO/qZnl+WgXaM/7ve2Rlbx/6LpQWTSlAPdweLF
OrbZ5XLnhqT0WWzzuDDFcpETIRBGrTrLbV9r/cA8lHcL58eIv9IVDXF8LUl7wvlhTTsiN72uIe0f
0hKj2lPS/0rtMT8J3sP+a57D6iWQLeev1BM4O4FavqLcND9+dquH1kTllQ5v5KwRfJoWiCTyn3M5
H5uu+sKPxtwRDJfG+K/JSdb9aHB/9u8322FKrPLO+oDNMAfIRc3T6QhIV1YqBAk22iBZ1bhXRCTC
7/Azl0Dy6UuMQaFSF5gOgkSqCRSGv8WeU3Q0wGRKPQfaqz+1jKEPHF7vddA80rQPuZijh6Ueprxk
L+asnfvxEOuKgHCZyN7Xv3aajP0J6euh+e+AuXpiJDPcwDe+IHvp7eyyTOtpagVbKY2pzV4sIOYy
FNmysBo1CcHtegB3nDaZ3hO3X1L6IlSppL5sJ66Fh4gl0s9rk5tJZvoL6OahV/9fRJs6+/dgMxM9
buzDfr6H5ar5eSzb/o4zGc3GxMQ4hJmkRYVcghTM9eSOJSU24KFpqd/w27GvQTK0B0J+rclXGe5/
yegUghTxSfC312QcC+PSP9LXbheLcyjYz9sYEpUklukKI0KZ5Uru87YSeob78QD4fB7dXYa4G47Q
2eUl5G5GvMrTBtdO0vksi71CwsQsdyYjN+GBEAcb3O0NiqT6118NSh0UD/gro2DN4NE1r+Whxeo0
hJB3ASG+PwWUnyKdmyLSQAPeFp4cftP6Ki+AhPHL+FXwBXMVrOr1b03PrZwbgZX6dqNly/3qw9Vh
ACC6fTqXw2wBOVfEALf53Bfka/xq9iHmvSQiOyaGIOch+H9mIVXkbCObyC2NRLfINwqnekdqWQln
8ineGFhhOg5uJYbf568SgO2UXsOrPCRO52Vfwh/fEhmdYX2p31pyesNnx6sHTXDxC7G+6INRrlHv
YkjBXrVLYAg9EygGb+58vgrXBkyQ7d+9tDgBNouAgmIJ0JOwLPjVij+n6b9mMcCoBUJzuJaUf/2S
NhfbXyziWtzHpCk9F1ACJNe3fd3+MW1WdM5MHfOjRK0pLPmoskgczeRfa2DjrcHHU6K7S7HVB/wc
aJSclbvAhdbnCRVIauU6msJs5DBdqoj8ljKiKD5YW2imG4cCvkgIPx6V8UcBDu2WYuOwKogysgE7
auWA2CISYyDN5XjYgFT5xIDY4dD+mNgrsABCee0PVDvaWbr8GT6E7Kyo7szzqL3i2QH0dFnGO42m
vjeFfpM0A/u5vbibf++F2G2k0uRqPliTfq3FcS0ZW1MWhmyfBjcwoWDAr4lr44giLc+VMbcO63eD
PgMuR8GwkPZaYPoYDIdz7Ft2Hw4goYVoMX1nKlebxpPE5ToD1V7sPr2yykPOv84KwcJSRZtI+O4A
rPmwe4TItQKJviRMreLXJmMIYx7MTVZ/Qx5KqpRWYfeHzRe1NTmIVZgHZKfuaUbd4kBpFjAz0GXV
333KdSRTPuFmz2HJhYll214Kb+WRgkPFthOfVgGu4fqZVaMyMRKFk0/tqrZFpDscjX90rCaQpn2i
B9O3EYr5cgpNFeFalN44Gk+fZQM1Tz7YL+av1BfvNbVJ6Wmj25Ssd/mceHTnl6TPesjkIlucJSkr
Sx6lzo3RzNjVvmPdpFj+JwBYPphBfaZkXGus9XT5lolrCq5dANdzhcKISZIsgmap7xYU/e1T/oez
NtyOK+5hv/2S2G7dNYX6T0GX5UgaLhGlQ+w1RsBc4KzT1/TJI5ChZjU5qTN0nbxZNuuw/qXESNJ3
KRix+4uaVCZV9/uUsceru5dtVkiFoB91EXZCUbSgLZyv1+y7dWEUcxvcMgQkDwxYGxbJ0MD2z6O8
zwH7S6jaqQjV21G78+P88oJeWsAQRoZKGJPl2EY9t+vJNyxUwsGPGxYgC8SzFWBLHQxRmHE91y0T
Bk+EapouGNhyoSNisp8gA99fkcFZpd6FIg+YiFpe2Dq+4y9gy2TleBs7d+8xJWMJ/NnUgCwLvq89
oqa7Bw6HAevz++DioGlu4KObhyXzvbbfn/UTqgqlPpvK51tTF2Jmmo77pcgFIHi9TEHhVyinatPa
p0kgqClriUGiQu+tXiWDvBYqRiZ2QZsWLv3dg6WZ0dlHQEPWkb0TqVWlcTbi7lMqKlii0lGmuuHx
lrRb8+U9rXz1vcfnB3PBNPFwE80Lmjx0O9ghyzkeayFDEjhmPrSAkonFvaWRxU3WHjmUVnpnmW11
Hc8bBDo47jXjm5WSpT7zhqFZCHCpnm2mddH/BAZ43ExRCGxC43gq0qmMPLKMnWrcN3uX2OH53We2
5Qas/mSLqXxihrzWeP2s3gyNqDEsEfWLhWsGgJiZMYkDk3ryeNJRW9ldbpCeZtLYbzYDYibote0T
H4oWurnYAkeE3SKXlteFB4QBLVEqSHTGODMifpzTwRT0VHRmGNEjS/k+z72AOSMus1m/gVocpxsi
u5mmD6vw7unscIidnjDfS+ENhliVOj7GvExD3XjpNE8K24juyES+bzkmJkz2Onz3v3xwRBsKKIdP
scBVEDq0DQekOGy9hfzvkhNfCwMmafdZwrj4+CNrVCbnSN+1Sw+GTdrc5kbeSnS37h7kB9h6NuyZ
JQnoI0276RpCU34Ej4VEIKfLaz9nfpeh706R6w5seIVW4HqVgTIPNIZsQUe0SPNPOgMruiUc8aFz
psMLfEoow9nM5uTJhZK6t/qX6zb5vzP9DAHqAVzrn6BJjpFhVJpgB+u+VKekYXYabScxaFQ40AVX
tCECtcEL7dM2SJjAyQeAc2+Q/5pSPCuRmRThzmD0rKrw7NFNVioUi6hzlYBCsWA/pns6K1jG8p9Z
sdiS/inST7yFu1kJUHnNfBCYAI/41JZF6fedrEpf7ff6Vbwoj2J91kqHcD/FGULcbvR78kcrUa3b
iqpI0WXGCtXrdLGmVCzUo2vGiKWhSU09BdZ3vn7P5fYQI7qbBkKiLDI7aY7DhevaOwnORjTb4JAa
uhpDFvRwftLnkSMGl0ZDHqHqxNsQ4vVhg9Ea/X1s1WNFwX4PQdWo7wDEl59epDwpRiBQME13M9hB
gqFhAfR7n2CGxNiCypTfRI4uLVcJ/jjEi0auY7hjQNpX8DVH34rlIYQMns0Q+7nAC0JjFJb/Flfs
bHWtV0F+PmHy2oz/RgGoPtx7yHjbWKc4EPsf9lYyzc1HOzP0cUnPq2bsdnxuoNQN+QOY9TMxf5iC
yjpLyClr7vS3YoWk7ItLKFyhu4kcC3bhg6/xDuUxVK6sfEBwNp73XXgNChECmB0iX3+syrhWx2pp
/grF22OqwJJNf2PEGc7c9bkUBxik1235Kr9RuL/M6qwa2KBuAfw1PCTEduGAMI6T66dlV0T8IfGN
26yXuOPWGyWeNjIbKTpZxpaJs/jGjwCUi6HiJWYFoGmn7aq1Al+5W1F5jcmgUC2bev5fFkcC87PZ
W7hBlOy7Qhoq/T8isBEAr99G6WPM3DhykRMJ+vvW3jpUNUzK23f7Ss98dnAMcwITHWDSbkrmdmdO
JdZcXP/nus7XYRvd9EvEtw+qgOYwdaxY5eOCIz1QBxAGfpB9CuSkRRsYWF/AI8pdLSjCmahik4+j
17NjVphSd/UQhWnzg3rc2L0k8Sn4Nul8jZ4xio9KxMwXNWvEY1wEfC+nu1zYcwkBSLGJJ/Zn7cS9
0VONY8NMaVGRi1pC/e8O2uQoUm8P9YQu6sMyZJnuDP3BIEF795+AcLJrN5P2L8Gfe1r0WwnEGn8w
9/WNl5EshEb6SMVw3kFMDcv/wYkdR4vOcMnOcRZ+KkYKZQC997/NUBJJo8pnSUPFg17zXLrPqLb1
D/24MTya8/MlwNijpaVDYehZCU6Lw4I0+B8tAuwH+f5fy0zY6bdDRY+vZY4AOaC1mO/Z+P4Ys276
vchp8v4YoqchkPSLHQeIIZZYXoqLqB5cSldLKespF+HUQsOouPU1LqafirmDEb5+pZylHOusdb/8
jsPcH1hTWnPKnaT2PeXTqMDiqb4MHeY1gzoGvbNjGEf6ln2bTWsek2kowDBT0bDEpsg7J8MVqKOX
AJznOv5IDHDuE8W+IfrVIim3KhF3vSPR7DzT8I6uLh45J1RWYXmYMpBN4kKaE+d0XoGa90IP7I+U
0KL02tpRSoFsqaN1zVVfcLfzqTxMq2mIc4Ti7lvy0uLyz083lYO4WUpJETXyAqVP1uHXoJn4RQTA
1IH5xbu8fJalQauekwM/BmKkYbAymjETihAD6xIYkpeoBczE4f6KLdGF7rPSfJV5Bq8zeEcejhRV
6lJG4UOLTl+NzNlpv9NjiFN9WkO3wbxLAnT9IuRDhE1QbRxzm3BTelqZSlcIB597KokRNpjsNWaf
k39LIWPXUZfaicQnKvLPsGmzJCpxpn/20LVCiKHiqRcWjNtUN3rZzxuf7eTC/vYAZ5x8X4GVobiJ
gQAePQyfzUVbl6eEIcZLGjlwMSJz8p0AyltMJ1msDKA5E3MtbTbWRijQTpefq1jgyUbSHblO1DPj
zcm7Q9MlUH4AJWaoiGQvBuJAMYLmaTjqX7xSa7BDFytBpe/I4XHchRLuUaTCZmtzR9C9AWiGadqf
RPlkchwVUgSej+TEUrJl98NKrr0r+Uuz+AT/NjlqON3MALt7SHCL0qHQzHi9Rk+Tr6YiAaGBbwde
q1KZSH7kVnOkle+K4KoO8jyJBlgdM8fAWtmC5HM82+MyKWmjFG+BTvK1SBa/OGh7evvhnIcDROTT
mdWspMuIDnyH6guz/4i+tHVng1U42COS2pkbN3U4Kzr4uPUxcyX/HxvFLAQU8uU7kAuailiZ1CqA
SOE+6y27xOsnr33rq5+WRXG7BIltLS45zjyGvJco1hMKjIPDT/oQXXvdhcu8XsxaBxJDAotHAVd+
W8MrSnL/QqCllHRhZRaujKr1w8J2lLqGxLWzYwJG4kZozspe+UzF1ImOUij9SfCPLENF/JhH2Btl
WApxDaLZCpFz7YICm+1nKcaD/3y235cgGYsxT1vZQhtPCAEKyCXeAavKvdyH04cU6EqK6gzqsArh
bTicLUB1aNkY82d0bpn1s8X52DdwVzSCyjygm5xUAOn2JyvN75ZUg/6QkKXeKFuU4smBM0RABiAP
Iz3mLK81U009jg3t8ZZvMBOa9hHgjhpzFUN7qHsSr0Er3IZ1ep7DGo+MWWH9H/f1s3Zp7H73dqWe
IGcbsExBoUSdbz00TSpTEOHfJPVAyjvvcZJPjpZADSVVfUtjqnxMiw5iPfkvffmEnpfRDxZJpkSN
65kqmUcNaXMG5TXI6+fmJBuoELXVpQXlVmJvgzAvmc0evm4a9CWGbGXhAhMDJlRW64hDoidFfF/U
6QoiQo639/eW+m7NF01Ulrwg0Xh9zWMxbAYZ/liFaQoKyImKzHw6RJ7gcKXKaw3Kp53jUAPbzbbv
oqorSO5z+bmp5mEuCn5GQd+dpWHWNlNyula21BeJ0Pc72lQ4HVj7nHq7dvE0hMEZ4oeg9N03vxlm
IqnfuhAt/i+0FrG2Ezj0KVE1zKorWdiwj2p6xaXvVvwzXvTmuCUUtqXzDitPjDYjTJN6aztTeuRj
pN2ZfDTiCBkN4v1wKwDFD2moVX+p8yGVkkm3LVJB88n2SjteqRU/1B+s738G97EhvescwaQbSn0+
5ZArjRVVrNSlFOSEByyJifrEfoL64gPh6lBBdqZ6J9BDu+WspCvA/IcVOOaqMZSvHNS62at1WTwu
5dDNMSxJlPuJl86HHJhmPPpxNCJuB5yq239DNBsH5YmDbLAAPX1HNBUbPKzLDQ00GHWmyUefrD8a
dbHz5TvwtEq88FyyI6EvlW1KaK41uIUhw62cQ1K/0Nz7EdNQtE9kja/jPNfeyWpiSnPLHIoquU2q
gDowSNiSqvFOk9LZr+XLKTaGjQSyfnnCQKP8i7RX78dZE7nMTNEbsYsxzkLuB7jMSp8gmKcqUjRd
p18ljGINoT5yEAwcQCrkttsDRSmajPfdShFckcfozxSaLJA6IqVL83cK4/GguAliE3EaIKT6vc3r
N6UxvfyZOcTEBk9TLYdmfi6B3FF1Hei2OD4SjIMGCfPcx6eC8vDoVF9AnUY5Baps5jnym0eZs+bg
prtGCH6pFx/fEKZFlHk2t7MpwG37YTGMlhXBl4DFoYVgVuu+SFMsgV6QQmFIuY9i0EEujgYQ+EDs
h3oDsaWTFsOfDQwuYUY+agG74JCt9IC4Nm/+I0qbrwt2Sl4f1tHMms5AuH7ij0IZNnwdwiHxIR/3
m07JDgjALpY0GCewUIs6ARm8zKs5tnVpOoazesCOuNQHlL5MVLPuP5NdFmcy3Cz6F3mbhpeAsqIK
ItseuKVqiRwBL/e/OA9kzNJBmoPR9Adf++TIyrve0DL5y6K08tb5q2D/nIAlU7UbEPWCSj0Rp+Iv
s7qqupKcxReCyAnABEwxbdFJa3YQ/mtV1xkz5of2SokM4eEOEIAMTvgh9V+bhsKYMBoJZ1swdGUM
0FvF8T8K3Y673Vjggw9bwP50+qDkSFKPJTuMz8Mz1Z//3ZA5+U2MxZEpI9jy1O2/FLx2KtTCKc66
IL+uEQDCFrsHOzSayN8xOFyrdQNoycAv4bITY7fpMr903SoKwc3V5+hptI7suSo6+STWVgHFu2Ux
DTJ6G+WD5I9TtOanws3ApxL75+2pL0lnN4pmpY6Z7H0F14ehRraMCihuBPF8/k/g7Y/+dkrteQ6M
Fgfqfxq8MFpg//kIbFw7O1LJpE7yo9vBsTB8uBc+GaQl0/ALgHfEIDqpF83+kaPa7UzT62HOihCX
lF10/S6BRIOEkEd9W79neBQJqc9A6tey2DjNzFPDsrI/oWBW7kVVWSUhnqWoIZIk9H1uTqB7pQcY
IbOZIJUrO7sQ8ey5UGWvyrVKsW3yWSmscsVHrPpW+FT8x1uLX+bzeEoVijsJRTv3vrgWZaW6aErI
xbBT/LHc0N54SVCKbebbctbcfkItKx+7msW+FQ69C47VD0Zwq6rBKUoVsTRQMy/iCiuhwr980AlE
Z8nDtWYRoGyK/9e3uBc1UAWftU/vS542xcJoZsHl22vLaBg/IWohAMg/yagLIJkhLUOaLs858UvL
N3uGECfZSxrTp4vWPrFY+8C1HotYl6HJCDtHD2Ws2YVtJZ0PYbco/vPGokEo3bilJsjw/2AO4yAp
zoBnUP/47GTZ4Y6/Ljo9u5T85SZTWbI2BSSy69JVbo6EwCKbViuC5g07rEcFDe3ET5zEA1hXC3Yh
sjxlM1TxMUgl1ibfa0ZZNOVaWv8G+ooMI9lhTHBsbPiUb9Y3MSTIlu4WBIlhacpAurIqhe9kPbrb
r+wsXDybWEkiOc7CIqrVcLUNcIcCscDGirlTC/pW4R4HAqswKVRy7k8WjFCUX9DBdkMyi5yi6t7O
wayuN2ZdUHGKPTNs6+Ve1i4sbKE9sUns6mUDN+FIkLSgkbW3GAeZ3mYrQzTXt21c4TZWkLT+VA1q
WXksYggO9foGMQoMV+LWJoE6xULg6Xow38uOQyVHd/a+m2nCJBj66FdasjBCKBGGuJlQCLQqbcZg
3RS15s2gPyaQon4or9dLb/azdm+UHtCJqGPv8SiCVqt91IbuU3gA61skb1MIcvEMLY54b/IxHg6T
RRm5koLYVc9EOwB23hXQrqfdDlYDHQlREFi7XI1Lj+mGgrmkWzuCtPMTWZ8FnzshFYdDOEPq7152
uXnvpURl8heU6DqKzP4vMvjPbZ9srHzcykHsK2nLjnbcZow/zWWOr94Xboyz9ZtXw3tKFuWNCG02
0oXgoaD2G+0RiB3zRol/5K34T4aZW+RiuAi6krFp71l4pX3/S16Xbzwir72IZHBk/3k7sopFIzLS
xV3V6bRYOatiSXBaeE+p8PyyMq3nxVjAXn+jtNZNKsnQymgTJN5p2iGPq1LICbl9HV6+/xxLJkvq
FsKEU/Ur5V4I6dJ7+ltPITLy49QfN8njng5NmMIilcTVmyvMJRiEftLa3UwJnBGrrb63oHVwU6Lw
088RiB3zXB+AiDigoAPfYbHhMN2alJ7pGW51CBsX1GwtyCk+vi9y79jqnXm2lRKQXldwW4toJVJ3
fo+ZyF4t6qkDIVB2PL4tYBEoZfPlA/gn1swfBH4qWR2qtSdismD7MA73qzGpEExlX8iqpLUgjFFY
HGOgiMnk1G3uMle9qJCUjlI5stlA5Sp3QR6GJWc/uHmQGAHLYePy7MMJRxMjZeevWJ923jIeWR4Q
SEy/ifEjjW9isDtV4B6xN2phg9Qu5d82uO+FnV4NawVqenYUEUAUB5p6uglAB9ulGDHP+c40D5+t
pMEYH3n2KeV+Ex39v/XActKf/rzCo9NJgQnytUkR7V/YRpjeTUIdy4WBTXL3jgr7R67DihbW1Iyg
vw5g7EnluWzzd+bL8Al2lLWpRJWz2sHW+CJkdsYWjce9MdTjeGUasCOWgn5v8fpRmQTWhUQA3x3/
ObVc3Ci1FbFcBtES34Ks9DX5ciJvwngWRrRNSHw86dDFnAIcXBWLKPs85pGx30bW3O4GVungY1XB
mqKPkwx7Px/RggGS4rNfXsE2TU+1REWeymgA4YUEzOw+pibvfP1e4UN2o1K79m/iFkvdoLYB/t9u
jHK570/6fgwMpmN0pLMjMyOr1+k8qb1Znz3WkyG0hQEKnet2gEM3sgQP9JxpHq2vyoesv+hSzV+1
y30C25oKnNO20kWe9fjbmtP3/hdUOHHZ+XAANWx0GvaMAglcEvonft0zbbvG8ymw+lva1bWkUr+3
aBCiMpRD7f4AxOFvaVvqAd7MKZ+Pq5kaLAqm6m9Cn7m352vbc/0BVrnrwAgeLQfzSJBql9EsxB0Q
YUqAun4W9jeqflXkHhsOTlI5bcOrrdTov+OWT4QAEMFlnBLIh/nzGVbHHFtlTu7536ErBPPYyfWk
NoBrdx395ggdxk77vt+usZykx5ZPX2qlhSuN7OtCOkjeLgU+wkWcp5Ppx6S/5K/mLCsTXfAqEG+C
qxqxQjLJ95WApEMcd08bkUiPlkiP4jI/U427SHf5PucYVebZnGKQK+0OaGlT8mIi559cSQFgNsSG
U8ibbN16UQd1pO9PPYPmWr9Pam3H9eKeMk86s1nSzyFNyNQ/z+tu3Ne6L/lCuclGRrXS3c3XFwq5
tCstJYVM3LTVyKXkIgw4sPh9IAQVgarZJafZgJo4BaxMXsNCakcSTXdZf8rfYoAiRpfKm8JIbhm1
9zR3OxV/SOdcGW5/aYHtrJAhs64tbH+nhHPqBJEMUzetVWse5z+3LORNaP9sDRvA0hIvfx2a6Xk2
uNxbiW+UDPU4i8SgTo/7J2Vy+I7r8B5dd9NiQolostA56nqPQnhDAOA+qPnZuCnJuxtdSq5BbaFl
WUjsIMGNHVg+pSCLxUfeESbphfNG/iyqr/U338ElL/9k8S/wmxLtyV1QrjUXbakjBoyUzekluZ0W
H7LcPRSkOFQwrKKq3CjNfjRJO60Nk5Qx03D12+p8sJQwu8MVM2VNoW5TfSkIfNk9OCg3xP6bPEnd
W2baULXrRuwNsP1OBPPLw2oUSTdRFvg/H9Ccx3Bd0I47Wt9e1e4OVmqRLx1pjI4X/IksXIpuBUkw
CMDPuuQv8lQR9RvsdzeCJ/7CCiSsi8X6EhD1VEKgGPkDeeuBzFY5BVozrygLnyBpiDIq1utkQ8Ko
L1bAkqqFE4lq2kTUJZJBuUVFZ7m8VFG24hf5Z/BGq9F+yu1PLQJBTLOQXWVo8dJcuA232fArVwJr
Tnf2WyQJCu9WHOm1nJ8oO/3i4W5XQE7teJ5VBeJVZOWgPfT+yPX9X2P4bMq8eNsMjqDV06/61nha
I30W86k4JVnwfKIJzIIxUSV8a3qWf1hNoX3lNu/NqzzIwPFZ9g/eGPHL0HIA5GLOEkthtJFiRyMx
P4N/kb47aa4f/4OE61A3rlOkxKgxh+j4fQ8wwa52vi0B/RALKmlLKKWYevibOkvrXCRiiYBMG+iD
/aUSD3/eVHMtKPdvXXeScVbw0HIUzvix/lidLZV3lvneUeuiiYYk4omUvz5OU0t+nPMDCubKfoi4
2K4pgk7XcER/cU+V3K2PfL2jsiKvt8FnNUast+FVWoXvrQC7C0CLMxa05KSwgG6Rrted+VXGEtp4
kIBS1WWLj6k3b6W2rRFASSBx2DGdVLzCpFS83HoskrWdy99wOewLx4WPTyLtBfuSDg+BSCc1ki1q
fLRYGHNZaIkJowi7xKPs+Bu6zSM+fl4phFsAIhQxDYW8uS67gbl8H8mMfxv5RJN+4z6UcavGAZog
n42ZIF+ENG7o4im1H9lETKry0bX9UTmUUqVstTqSuAJXPIeML0tFahqzob7SEljuPkyXj8BOX7Uu
u9WhHQmwv5+L4OUNzqoOPkM6arUb2gILQRGOeHkf2bhWEj/oUwz5oJOWzpDhMkO0U/s2u8rVX/gj
w9POhJkXoSha3ViF6m/dtj0LY2cl0ejdgQ3TMWSF5dTJukO2CIkEKPUWzP3AQKa/f4Uz5TGiB6uf
Lpkz8ofBPbmOIn/+w/WlWN/HarA3iD0bp3SjYX/HvZsyYCJMNehOCA+tTV9KQF3nC245CkxWxxoz
W28sPE4dPaj49uSR4i1K7oLSClZ3q7XkGSGvOc4vbnuRCECDku2ZPtJvPR9hgChbCvBaHseRreaO
w5VZq/GIOT3D8T6M1mkM1oLPuhc2pWZAGJ+bpEUZ+jN8hs0649I55xy1bw5rFWIOgpa8eY2DKjFf
vT3qBpIH6VqXFnaAuXggfa1cPmFWIS2RG+JuFkJZl+r4QHD1G+gBu3pzsS8MCNjpUfhr1GzbJcZJ
SVmhJKhqh+Va0prQj4uPGILtvVl/CPNH2dp4nXOSSVLyRgFBj2T6FgreCCJ6dnm2nERXYmkKZFqD
Kr496zKOPAfGYjjl7P2u9m0jZjSyJBXwade/oRc8UrK+1pgy2j7fHsQ0ZbwWpfgF7ZCk3hV7+8Ij
fK5ulgyABDrgzVSkWnVz3AO8ykuUINQUgeGllFD2fKcEyOFtl/CQ8JWW72X+gl5gkHhIDVAvvnAE
P9TrPzN5YjULDjt1JEYbasEYzD4y0XOuBMHYFzB7yI3kI2izWU+rYTD2G3JGEvbnlKIA85j92CSq
hwBvo3+Nb6OfuE8MjTpHHExhwkIFV3GqcHqVIBO7TNsk1Z0OEQFYfAXebUSkm3uGOQtHOj5xIPGM
szGbl2dTLNY68kwgMYFvmhGDwmn9Fx2miIWXzxgaNEg6w+rJz2lmdsDbBRGQuXB/S/WMAHeatpBD
Pj7lIP8FjSa2x8MJdR7uToE7X1jXE4x7ErIirT/feSQ7Hv5mEDYLAVHn0und1odROOh9XNq7ujPO
6668SMnE6Tcspa4rl2y3cIb+rhEIkpJwgzF6u9z+t2dg9T2ntDs4htaoCtks4uNUlPufkOXMqrpM
g+vJ+mvwTLr5NAAwpfCanwrtvbm9rtPokdjQXIsG0O9eOPiy+RcM4gDIumZOyOhpV7G/IrkeBPtN
FCGf2qdIRJtnX0noI7OBY/TYqIq0cK4t8Mm08OQzfIVQOPe6XGGpiVUnsxlgTVt48e3xKQmPCqmQ
a4PIjXmvOLthUduDgJEs32BPPlxe4tmac66tVUr8rX/GAIczotoO8c/YP4q6apKsWEdrxzlXGKtD
US0ihNjha76I0bSmMxnC0Tf2Rhakqrl0BP7bnm2eOzZP2Cv3/7ZQNrhTTfP5VPA1RmK4jcQbfTid
g89CDd0aYdoD+xOYmKoj1itFBwD2+JiAwYhu+QYo0bBDVH572XPv0ig2bilywyZfSMSthIePBbB9
FWxG3aRCM4tpgxYNcC+KJ2vKqt28EkcgK9SHFY1IeKsuvdeRkBV1Wnfi0F5PRUN2hCQ4VbgQRusU
qPE9eZGYFy6IQVwiKWX1noR55cOtNe8fufaCjxuotNPbuKRYlzKrQSwKMOPIW/HVnRog+2+PFYE5
Rw2AlWPPxnXq3LF8hfD4L2m6pbRFdU6to9q7N6HhdmyO68J6LwORVFBDmZ1EMMojOx0DcwR+yvLE
Qn93BXRH8rBYaaLOGLiGNhsE4VEyZc2Yj9yTg6MkIVIM99ycG8HFZZYW8zNJn5BZIoYBp6nEszZO
mzupDWt5nOOTjbwfw7lStkGNs6vr2McY9/4+/H9vegHQblcNj6aHpXMKiwIZmgS0jiR0tagSYHjJ
dLffbTjGmvBBUtqcDCGLDMRd2xg9QkqdJDL7YmoYnmCciFzZNHHdJt5ci165/BsT+Atij7xzS6zu
UQ1r9kaMc1glmXiRsNaZgu2tP/egHH/Ds1koaIxkynsmcjooWrUJTT8pU69YU606e7fkBNTaUmRN
Au/xFcpYgk/c+GfHGY9KzGZKDUj9iJLYIYqjXFOJeAq5d+FFRjXwQJ5deE2r4tHZBuC4p/YzHg4/
GwtCVDSCwgg2wvQTN0QKgrnQsktrVpNc5o2B0TDWh0P7pnKwSM0uWPMp0JyHRFc6NKIjwxA3qGJ4
mPsSpQAXGZPupclDUl/hn554DRUlaCjgJlvfhT1Tsy7+US0eLgP41RysT1aE9k5Lbqb3QyXkI1D6
zyADe4gA3JZd7Jilk3+29RI52eOTn/sRazrueV7dM1zD/XfJYCMfgArRf0yT3mk6YZi15W5q+8lE
OXsMmlH9XiC10a414BFX4eRUm51ptxHQ/zlRhA63Yxa68kcrZ9EWd6ZtvwkUA7wwbxz2xbu2hfXd
7DK4KmwyM461FvUldhwzEGTPk46mdBxhD4XDWpiywKtL/B5LjnkbTqR0aO9dpLSamFzk9VquM3U9
tAaSFnf6mIIO+N6XMfX2w+WCKkZDmUOkjjoMrbqAlnoKB+lXPsMplBnMhQbiO59TRQBW8Cr/PEtf
aiTDNGhT7uPCQ6/x321ljtQm7o6op5kgao9stdjoWRiiENP6p4LBIR+uNw+WLm/neHXfjYAYO+Qt
3R6vqVl2A/evnpiRgEGF1b9+nK1aWqeEX4ciqlONEGDkAOSVq+Z86zZQfCCEyr4dgd4xrYZjLfzo
Zn46N5DvyKlqA8TjFO/FvrJ16ERHzvf7o0zVaZ6SZlCY8W3ZSJSeTy4y2Z9U5rW8GvEHFDEoylZD
6sgDsB04ps0BPxhXpPPLJSUmMNwv+FJt/kGecUgt6T2LnC6hv2dwC4lhiQukCFaTO/7SdrLrj6nP
n89GJB9lRKbQS7uHxHekIcAhQOeB4cHakdy/wXwHmPnU339FWXIqId0CON/S4+Gcva3Bs+tg/pPe
N1BWONJruqEWFtIimilZpkISajmhzh2+oeWHC0YjwRQ1veEUeO6NtDtRUWHZB0BwVwiEtdZfb5B3
0EUDvXm+CSHkSy9tbaWdCHwkKduKVTvZjxYz+m5qSfiTNxlxgCeUJthMnkc4jTIz4Adtk1RBjB1Z
fOHV6PHKekWH10dgdQmYie1Rd82yp6eEQ88c/FraBnhkZdrwzLrbBmKxTz067E3jkghNya3mCKYK
S0d5M1HiPD4Vh9TpBOeR0NlAqfneveKeNgoQaFrLajdsT2CMgX+z2r8wAKAT15mcE2GCJ4AIcTlq
S35nlVgN2Kf3AA4EAP26TpyvCAQDJorkmfclfec5kQsk6T8ANFgyVh7xNb4181z1v5S+Df52Q0fS
T60117jDp7VpP1j1Gj+RGwh+f6hxrtD7jqGuD2x+xfC/sz59hwJihxkyHs5oEVOz6CpVvg+tu4oy
qBDmaUFkXesS/Ov88YEJeBrSQKODPY03K7Xr+bJQwr0AIIQBQe8Mfw8rBAJciz3890brzBw4arkt
7AjBmmWuxD89wCzZGcCq7boWM/8pf8QPbyMjlCH+yNHG6jQyVGW+d7x20kG6t1CS0Oe/W8EpT1Vx
zJzk8LxYbgsq4Hd8tWcNmHaqo2r8MyHBXU7X7Nk75pVPtBvsWGWFxO9ef83ouATxUEqVpzFEs+LL
rYg3phUAdsrvH9dn0nCTtAStOG6nl/r5dBRqn6S9Fk1h1OnumtHg8+gi84n0RoDxXDoZPjgMh6GE
Bc9qhrYx+7We+KqTL7ILkQ0Lz5U8zg9Zp82PaFZh8iyHySQo8ffwPVGkvnIGzsASPqOCtkIY4TJJ
X0leSQOXEkInlDuawd+oYw1Us/2yhfIuTnWNbF9hxG6LFiRC9rs6CPSJBd21azrVkakh59XH+NJi
lMFwiKPFXiIdIRUe1LIbklGSNEvHCxd6WIqvuimUJpuQMrcjIAB7WEtFmvF+P7TN53X0tA/SpKJY
hic9MFyScN40xMytGS1Hkpkrl6NHubKAo+zeNcIo8ln4Yfj69K6v8Tuebk3lQI/ZKHoH//ugC02g
iUkpKhv0vvR3f7UL7KVeFwzZuijhvdxQyWG91C2gUnLmqA57zpGQ0JjzqvwP3C2D5xlkZ7A/tDaE
g/sR/OCqWh5AXW5TUrKxw1Ns+dFEaUEEZtuy2t5DnxtCQhkP9Gpe2CuZslMLoIig2hSlm+7ITFkq
9hJg3xzMaPLUxbBk8J7YmTtvW0+GsjGQReJxFMJQ8ntbjYVus0NaWYt5dDuHtfeY08Kw88Blm1l8
o+h1vioYMf3uanv55h679rnV1TYBEd9YIGZswOPgpvoRt74X+TUcKvoEDgHW/9PMhRZckHkTWDSW
3ABIDdtkWUNTzuCk1iCGW2WVmbgSYz+fuXdkWXotmXLy3I8FQuBlRbxtsfke6s+Ce7xSx5+iXbtO
tmE2wmISMAQ3JRaqgEbL0cIYhKUmCAWpdrXF2AJlTLqGovXo8qaWIz2KrZ2FcP8V7lPweUooi2X8
FhRrhVlaSeDeHmH7DyyNKIj9FON/Mo8xoi7LNcK95yOsS+yqdvHUcUTMMu3AeW1JLtaxzBFK2shq
ZC19e8R35jEx/fnBVem3bTozJTnSfNeArPfeKhe7fAwyZ6dEwtcJhhOlpWt1YH/KaA6xj9N9zNVu
4+oSBJgtYkvUTDekb9+B0Tf4EN3IyHyHp53blfeWGQmvXiNBFfV8m17zlYCTvbus1bGVII1pmdBP
pjuzsUVsPyi3I+fr8NBIpMb+/nqGXSna55H6ih1IAGPgpL+D8jI1yhiOQeTlk/mOVRULBZ51QDbZ
naWzedjJ/djwjZV7Ipupf9TBwyScwqmsQE96ox6U4V6+E+m0eNkP0gtimrnMhDkEKmMs3Bl4T1x6
GY2ipgKZTcqghe3MhmsmGD/Fn/BGsOVlcEwe6FJi3DwQHaJZCBCzYSTYhEVaqHGOIxRNydjIQVdd
ipycSLFikvoDqC1GtAv/XpOs6ZgNIJhxpn+UhsrrN7yl4RV/PO+eShwcYqiXficRYAQ55d38mAAq
YEvqX4XeCpPPDIyrqUlnuEzhpU+X3fnwiyQKxIjr5gCKLeABcq50VJXS+AQBknmpkhFXU9Lu1FFA
6Zev0HgIlngfrSWd6bLGL1v/g8IeWFccjpi67Yiaj6TJmjy76dx++nux7pHsPnkJB/NOFMCcSoJX
hH64X02u0Gv9oK61lNhes0RPSsrmbQ0Ugwl3fIhFiH+l4VbDYX148OoHNkDeEuVR5PzoTp324Z/c
Q4svH4SS63r70dzV9TMqzOhd1/iALCIHGNxlWZegp+do0aw4AEaVFQBMAHR36GqqAETkzOlTcUKm
ZSOuWgtb+XRpVy3W2AFjJmod06iuj4uS650mCPAKiEPWrw1Scd4t6LaFVzF8hY0ScyUJMpPxZPA1
qTNdC1Jsr7csEEkOJFj8HFgbKtA+bsOvdCsl6STWM6+mGMphlmQsS9iH4I0UGDBfbJyvt+kHRMii
b2TucTaAwHeAZSXMOq/jGaFzHczJPBkYQP3SOgQLGQafP5RnJaX1ykBtR/fcU5QQekXI82tQAhtC
rejl6AtrVE2zev1yevez8043ddRSGYInAPjVONo///6lT/Sto/tA4p4Hb3Bz9jtm1RhmgZQwneFv
nbi75GCgfPk9Tori5Bq4c6v/hBSp1IoIM3GsSCChpBhS7TI8kj8dsHwaGhQqM7U3vZ5JYVjy3m+5
jA/2v1ehlpa5kGOfTCyiEuoGDKXl6+s6uDIl8ccRgvUnEDyOLPfNVW5dT9OLBfa2etZaDipf3Pgr
lEFZPbGzcaGQ31P0iuLXW0v1Ynx/A0Mz9BbQTIs6RYE0uHAg1ztZd3+KTugzRbnD6REFuftcfPPk
Edl8syzEzN05lJRYyYijwhvrMCHEGom9hB8E15LLtNa1IjHuZEzEHU5+10TA3Wqq4b0mLTwFxg7a
YMc/fOls+IQgc8MPsksl5QNdi1lno5+diJWBzRJm6HAObhsgKSlPZLLbGLnojO7zmKsjnaKask5z
WiaRLyUxLW2TSB85KI0GoFj8VN52oDNll+YqSGVlhzCURpODu09kmUCcu6XPUhwy4m9z4+/Aoq4s
txROnX8w6+wyfaOFJwipaeRRoqaeJVBE1F3UjLC5NQJZgcfT8FZjy8SJK8qgBzvVqefj4nKRIlnU
/JYoDvyl0H/+FQKe7Qlv7kKfs+10x6+N85O/tMgOQZ5h1Cr2bJYhT3NjJDPzQPHCE06IO0Ja00Fb
7RkfcLmBCOJ0YoQOT5UVM4vPovDqHBdcrrOE6+o2WYwGXjn+P/aOod6qzrQPfCHZ3VTztcE8f0Ea
EVk4iFZMM9ebDTLQQeRteh/yYP8jtiSrAEIsIP1nwZcuG4UBr3WfZgh4JVEAHgYVYmUleSPLqNNN
57hxlD3UiLyVfjBMhPSXXZuddYOfyUlPOHj8ffpxiAOyczuECZ8Lp0D859k62BkTOnGKCFj2ZmLR
zSWtWx3OLNYSXSF/PTh0uYQvdfFTHzdyCd94HxArxyXOcUX4HUbmSNVHqm9nDd4+0iYe2jP5jAxi
CG0UXBzTx/x9jRrlScTZo96FbUeN5NzMAdcpWXY+u1TVOszJmFHIMFOevbSUIwzJ/rsbRe/1ZF6T
KKXGOGjrBuyvERtzjgiXUyGT9m2Vya8zaNJVjEvr7jCZ9yz+gm8RkJ1OA2TfYKQGTSUmrSwHP1rd
Fcgx173uUluKL/fEy4Aifj+dYE5jWKsOzGYBIDvoWcDfpoDL1C+s/Dl9uTWitlj7rflE0VArvUeX
90mzE28l8cHAZLNMdPWqrfVk+rJIDIzhFP6KayGfbEc4hh5+Axt3IXqa7+/kWamHLVLM1iRhJKJk
JhtvniJmTESwfk+938ge/l1Cip2X+8S2l5Tss15UUFLNF601Q4v6y9lcWw0h8HE1EKvO8hpORNTs
yobMF7unjoxKE/d42O4NpZyZ/A/qelSAQv5WqOmbAnsmflKqBnhOqHtQEuL8gUuKU+3uFM/abSqp
CusPFPmHaMY5sqjHKkyoHFV4hPkJLCoON820PKeTAjHXeUQB54XJl0Prrd1qk3E46NR/aWajLkcb
mPhm+y1yEQaNbvc0oSwHIvAT2ZUIeEPuLd1TJGPz35KnOcDAAqM1yV3Xf74uVmcPeqlXtpbjjDhd
73yIDUo8dpHI1DlPR7+kqdszwaYZoP401pLXPMjdR7Puyxci7xWZ/imH+xsf/7GgR1lCzfa8W5rQ
tp8abIDpMlJPzsCpJ47IbKScfg7SkWIulUbX0r2bflNDTvGNSa9xNIQ/rnTK61uyMibNqnO0Dzr0
FDYYoJF6aNE8bZ2iGYtMo9e5iBDgCVtmnzDRsit5NXIDQnSNtSuFMUkq8wbBX3oZrh/+YQE2FtMX
qeKrHrr98Fv3MPKTk634BZRyRuWNkpTaprjWkwk14mAYNPcGDBbY/xTGQZXStXs16qF7Pibe1cow
lNtSznL4I9jOiuznidZgcRLtKmsx+qYKY1nW+N+Z7PiDM78mmkmeiHlRj8fCwLy+dmR9EevAoynp
WXNcLAozIGeaCbccOdrFdQJcgco3pErB6HuaseOblH4I1gKSWfym6jyfeVO67oqDhaEgwIwPyyVQ
P4vBBvul8LrykVttomt0v51N/OOa4oWtPnp0F5iqmjkxx8DbJYn+K80AU8WEFh3M5CadjJAEt382
05B8rBGESSJ8mA9Psl4dB/6jV2h2+5VUA1vqjtSyj/Ugv5/f7hwR8ACNybTl4aPoK7pcYvpKApp2
RyOOcd0PI2gKABlADfNQykkK9Ym4lHqB+b61gfnvCjmcFIBP+UXQ8bid+yL1+BLFnvgS3ZHVtQ80
p3vpC9oTOy7KWKDBN24ODAOyRlezajWQgrTWuG9y/PFlQ9VjkK/bprz+GGGttpWQyHEZAYGU8lK7
Q5Wx3pxY/UZAt4AMTuU+fXBmDsEhNyx2bCwXM49n5Gh5uKSQCrb9PoEkKdWlNZvuctoBmL0Rfi51
7HdIjYtn6SxaLi7DVZhM94jTjyJWIpL+A9qz6M6ay+WBDDgV0SFgdlpJxvDYG1xI4dOMN/Jaco19
g+zQ+PolZq8HfxBy8ZWKG3ivp7hGZxyLdc3fDXqMSvx07ojO5NesfWfElDs7ekZDB5f+ayCdrRbb
AnU0UbnKBxh/8adpiq0XYAN9qAwzY4mXcO10Xbep21ugNxevA4B5fJlGnUM1ny7JvduuFWSNJX3E
s2HeB1t80JX9K1d/wMNVxpjwoWAN+3HngyznDKGxwZQ+52BVIJuddFQNyNuVPJElNiusdoIyJ8IA
eWkb9MQVK/g59VOCfX+v281vE+KmrFq1Zt2y7SapxNG+QsI7PKE1OPOwrwR0UBZ4yq7cK5Eay9EL
L6p2XYURaV7loMIE/ug4kU/aJYX/cFRLtps+0LC72DndyKn3GBr8vNjoHaJmAlj5Abd5/bZJVEUf
3tihOWB0HLq8RdniSJIG85B7ndTOSR6jgIN6oG4VGRVanVA/BGHJbh7Z067FZgKQltUxlNsFy6Ol
HPIe1cdteSsqCgDUapJ3qF9QReozQR2I6QMv9V6/qkdVIYxj/sPvIlDQeaQnuLn0T+4ub38aPO6P
fHSbX5+YcywwCCV03FoqC+O+K4I3OH5mgnkcsvKnmYNukVRn3e/nFQDlDPqsVxAYEPRouZvttnXF
GNAu0yVuMbtnWMEalRia5I/wWfsJAQDyG5NqQMBobaJIa7OTSKC9j6ht7sjYf7tVY2ugksrwAZhD
eVG+bDBZDZgWGYuEBhEphmV8CftZS2dxbWsjhXnPPeP/YXqtbCeoUPbixAuaoe8sy9D3BJzllpj4
0fby9s/otWR5WbVAvRVrK2MCSpU1eYTnV6A8Orv1jaKm7A37AZ6LmmCN3oxK+7VyKtJMDBk/xjC0
rz77w4/QxTjzSnUDJx14LUcXgFkXasHGVlvohmed0QL4fxX4LhIw6JPDqIG//zgp/Z7lfEj4Hj9Z
QwcmE3jkeK8UHL9a139cvQeF70or4leaj4fqcg4rDWY7Kw0lS4hkX/WPlwd1FvhHgvQDPrUJlbIQ
9SryRs725B7NKJQ088xqnYTcNJ3TwWkoQX8Sq6Mvfg7qSgOOTNQIWATE9As1B+2KOB3XKQUZ2JKg
aKohBUvn1aRi6dLyNSPxezUx7FMucxA50SsvJ6YyOOvPvJeJu76iWr62GRoeMSkaqHCzQZK5KYjU
wMR304Bmxji5JztUfwiWqK5SOZ7aBRnL+U1D5p8830Qc4dm4zhoiavv61yWYMXv+HAkt9YE8Jv7w
WQizB95mJH140bbHb4d1BAZuLVuC1BaBWPZagiZfHjJTFYx7tKqx/aTMkzDwP04AiDcTa09Ajc+o
i+oKccNuiT0096OKmuITkysTfDJi5OLcZCNn/cVDO/91+RQEcQQiZPZsXG/okqBGgda0oauUsRPE
u46VjWllLwXD8LzmbpKyJ0WDmCVhHZAx48JHsEreuHUEHsSAwvH8onmsHIAVFjZ9RgfM02VST6xV
1oS4L0wQ2VJMLucifn9pOF7iA6e6rdLJo7qGdfsuWYqq9P/DD8JVv6h2SQnbHk7JD6tgFA+E3rlX
eC0feSW/J0mXv2v9Fq2TpiPgATe5Bwr/xB6b1GE1qaJzPlNcSzR5kcOb9amkWcTeLnKJNsPyRmaP
hE64bxUXb2DoOQAdCOIdXMWCwMoUQmBttdmQd1G3bfw0l9RxQueiaLU4ln1YJ1baG4QKUShXRQFZ
/Xv4pcfjwc97xmq9zwncWNpLQkc3syyuRE1mfs45pDCvLd2Ej+URe9LM1aI1L6hulwKveWY68Rla
jV7s6E/7DSIvGnPZeVhNMU42qEsoDFnYS8mRDlPKsOb1xKQeW1ThTxpvHXq+XStzPz9tknufD/tE
8UZKLk6nDYFy9prRrC8FuEsr7gRlQ0qNoAHTCIK/QoEXw5ksbwrDDAwj/EKcj1OJgzjV6erq0FIF
wbo4j1gXOS0afYwZ+A6CI9bbkrS2yEGIJ5B3ryf+NZsDVJqadxBLB9/syGm1wtPLsAEaanePc7nH
KuK7+D2GgFesn+PEGWyf8fsoXfKahWaeDmX3+c9sBtJtScSy5eFDxiz4CKoVOxVNLOb5jUTT+PvA
7idUwntY+lxzTYzLdF4cHa5nbYiLehvNdU6Ly5nHFCt2Vr3vfK/xRxpzpTf3AuY09uRqtiGNNVhr
SWLmEmawEP133TiZFj3p/eM6xgPEpE1g/l/Fy0M50fSeGu00vlnqXGlCwfkYbRj2NUjeBW+r8q+7
yaSzWrDhKLaymJXMLi3FWog8Ev+kxJRZXd9g9gcVg8kFeAewU5QPX7Cf+bVKJUsr/1AjqEKFjA3u
F3h/YlTAVHprbi4w5m2nihvYqnk1/HvEVMP0/0w0qnv01MdiBXfPD4n+gh/SpmMN/mDjHg5emlLp
TsWLdD4AV77Dz5x/mhmqreVwN24BAzfGYrRq3Ow/E+LQwcOuEMhnAfcWcLD6FZZ/ZDkuQYWjnU3j
Qijmd43EuNVeKyo9x7gNH50DOAFmLlYpZ1q3aDESxcFAsQpSFEnDyYvpxlTMFhPYb9wUDmDCtAeN
yjYFiUQr9YgHmQH3nPOY1tG7e25av/i1WKkF1sBHu1ki6vnk6QL6/z6zkh6gZcrYC/NkDesT0wCJ
o6oEswEwzE3ZQ2O6xL2PIQ9b+nbsvA/nN/CIz2Tb+oEGrI7USvIhTRQeoygs6hmAwIDCoQjC84W6
OQ73Q7LQJGJo37xZ2MlVoa1sQIxhHLMWmOdh2vJrOQlUfjhJecrky4JQ8rI2EAHL7530BFE8B9Xx
uRKfkJq4CKfQG1SAqo1cLUUKJUupg0R74Q0Ugq0EZRyM2f9uTogQf/EDYhU6VO5qC0hu66DPpqxD
elAHtEQRVVVpy7AkFd6PvsCiMWNq/ZKC6nFp9SqKxR1NWV6T9nYw0t/N0naPDlDUxVTWSTD10xEz
CCg+wQudpp9y/C6oRCMjjlUymfsruxM8jpsCdk3WGhVYs5oiGvEeUe0x5+Uvwf6lWT9NEFLbzoXl
HkNVZoygb5ml/kSeXiwgOg3l9taOEDj5IhlNDddAy/5PqXKOHLcsAjJQWoHHbknAGx/MtgJVYAQj
BDLw3/hr3I+Vrwn8o5jgw9YeiM8DW5VKFHRN8rbEJIH96LKN9mjL4oXLHB9FVF1NzXRVZPkgholR
4HBVSWuJhPOTmck/IwznhpnL5xdkYFmxgt89LSydBDaxmQkZHrJARxvkssqJaIbEL0nyirOpnqKb
JmsoSVSLus6E9TgeJsM21tqhXNoLg4rVIxDZe/zfBFAxZc/QwXuNRq6Wst7LkspL5RSID/v6nMvb
RCrXJcy2cwBo0GDQqAZ05bdF4zCAlMMlDGlIke5Sro9bUjEaGbP29/qS5ncyHu0d+GGjc3F3Q0PZ
+9DN49qZ2h6kvptfyr7Jv2GbXZVHY4GgoJgIX2wKdHdpedma90up0nk4JJSD8MwKgxFcyJFgPngM
AuQpyGQaECoeuJJtcVASkaMHSsUHwuz3et3M5bqbAYPTgva08niKT4JYNJgoZok5CRW6pid5fw1F
WnskC2Dhqwif8w6/5JalLT7X+U5RnPMvnZqPLAA8Xex7FN7L3W22wXOFIgpBTy7hviXI/qgiW431
c1f47efZU4of8/STG3mLnTVpSXS9sSrmpjgGpY7y2rVnRtGozKG3qaexsTneAswZzHFwilfXLNdt
Ooh1MO0Q+O/KqTItVs0O5pZKlgVcq/HlbFwE4uM9ynnfa8S4KrrHsQJ6Q8j2djFK8QDsKE6oQyW4
ryRYvxrJ2PuMJMs2uzeAnLuk0B6JcLmHksI7T4kk7eU9p7XjAVM8Am2cqPftoquglQjLr7nC8So9
OOCNMW/FEKvX2kx0Y/GLSnl1+Fmlg397R+G/Js0fIugRHi4l1xuqbUT0m+XHE1OXFMBPUkS8sz2r
NuNHg/4Gc5lHxeDx4TVq+PkCFh+qoiGTK+Qpvzrg4t/bkjum0YdTsw6ny9EzW3S8mC1m56oPYyjL
iQdb73+YfOUn5Vpybn6wEhXAyuF4dQ1WxUSiGHXabL+0fWJwCOt3d+JMcbFw5R+n2FLj1IpQHAsX
4Nxe8A41Nh4w6h6I9ilwvV3+wCWrb4axoojNpnVa3bXTI+B9G5ojAGjQydqSETfIOTDby6aQiHrf
p2OJFdyf/v+43ty8B1k1VLj6T/aQt/6SMiA6LcGQJ357rrvLt2beS/rlpqoAA8yUfOhEPa7nNCmR
aXYz2xe5uYSZ9FsYp6MvkdEBrZQ6AfE04UTEup4fO/rw4P24vzrLolkRJld0OAWF87jklVUDwAsX
RaBlXhNvaYnwzImczGJ+af0QOYcTVSjVNztVtDwls/lboUX3+yC4v7I9zCE0oI/G2hgek1afoZ6w
4IR0fh7bOBuQysKndVV+NBqxRgL/m+nksDMUYqQPhn6/5rzKByl/FDgsOY9j/9hGFyfqiJRHu9i0
RYPZttbS+/BFRqlAhuafj/92ph4dKFcFKL82JdTrdTTIzCejzYp/mUazrnJ3x1cdKbTWBewJCPAR
7wtsDauQfbY4zMS7NzD6yWmbN4Tda30zsn42j10mpB21bgSZeddwNtSuOIud/6RaVOPuMKVu2vUj
x7voJXlWD/gFEvRHzFpv2fMVV2NzmPDzm7iaoUnPG/RLArrIY8Ebl5jNub5XYT9k1/8ksH59k2NY
aVgkCVnV5BsmmqYgQ2e63dhegO3I7YO4Rxng8KcLmjrUv1V/7mQt5pIbfNi0W/FWJWu/4b5Hx+zI
cpOBRhX/BvhcIGTKTzXi/rYWR+IUsaXuNzd2/Upx6wsQDMERnUNr8PfwOB9LN63W3TA30Z3/hG8L
/xJYkQR9ug+/oTV6axMg0IyslTGZMHezLBo5ZeM2382RwJWPU5xdif18VkcayhUNcn9pfpOFId5U
QQw4Bjq7mWR/SKoEpZC2eQ91whZ6doB8Jwoan47QbRgWexWVTFZMTAGTZkyNSbmX7WO35AX+u16o
WRyerODTjkoWQeSLCdnhrieqf7UCWnV9XvF1KnLZrfi9VGIl7pItU/Oh+T9ViP5hdc84k/b/qdFa
3TUL7nk5i/nM6bgq+vNKG1ET0sVdECtSKJE69tMKWHBAT8nKoIt31l/eu5ptv4gM4D4JLP8PrZoJ
8KOHi22pIySfJvSxpzSLeJtJmlwPVjusqggI4xNIbGsG8/ta57iOSPYWm/m9KzB49Ijkh5PyIK5n
z1SMH+SBznx3Po4jrV5U80p+eF19P+J+Y3tIlDCPAyOh3dGKXztwbu7hLvLQrFXiUjBnAyQAvkZW
icJS5hJmPUZMq+JbVpM8f2LvskJO6WR9e8LNQq6lHTEIa/253UIx0tzdSQLH591vAcqwEdC6p8r4
79zG5ppfqZUW4CR207zbUvM2RdkXY+Joxoz3hAyUAJQm3tlHyEBvIk+ZUD4J0BxQJcQYORDjeu96
vepKHN9zBpsmyUdKSZ/bQKbPd+U+WdCcNbDl9fwDyRTDA7OOby086m70kC3772ZxotCuu/u6iqdQ
TFtwTX7S7sE7sybM+i38t4kteiFlTN3rZ6nDP7//O+EyfaxhEW/nKLsv5LX4zJ9NxrP6ehsSp94o
AE0QmEYVJUCBFFeZzjgufbTz8k1nQfPtGTXzPPNYrxxpmNr1PhxJrhidJHolNJoW07d+y2HyCiUQ
p+6ZnHHM2a5mGG5G+yp/d/2yZcWDxy62WxemxHujijIYQyJVTdDeH7lxZ3Byiyveqi77eghPH7v7
swwm9Ya5AOGp44N6rZl0zgYa9pQA2LznrQSw/YRqV1n1b2/XriZHyEAuF8hhqXYxit9DMPMItj8x
CbUGXjt6RtUg8jnRshoyAzvTpPzrJu0O3uAl/DNvCEbz1sL4eXPhjUfybqsyL2fDMOtCHucvO2Gm
u93739fZDXaOmv/zGqs0RX5u9oZ+I59jsYB2RUbTknIpodtRB8AE/l8ciIsR9Q0mc+siB75kowTQ
0Dv7xw5cypv9Vt5+Z9pIEvmZP2FL6mb6wLKHV/5kCbwmBQoHdgYMud4w3E1Y+qH7hdzD+y43l2EK
6Fh4EQNbo5TbVC68FcvcsncCE49XorF41gQyezPx1pXd9EkWTublZHHHZjLe6mGn7in1HSSJKMs/
QION26HIJcPnsljTsCCdf5GlOo2H8eAT+wpAMsBv9FAu8wLv6dK8ZQIPYJczqnyACeroX0CPHDmP
u3e1xmcrmLVT+SRjNHThhLwxF+uIa9lg+/0FrV6TlOP9JodoM3Mi1jPDl3Z42rvyFodo/qE7Lgjj
DMFnT+VCc8zF4qj4d9ZMlNb36fPA+wgHA5yYmne4ne4buEWC+BFIhPp8n+jfnk1xIlxD7KrFD/WK
ZPiUuYi3WTD3Jslsu+dnFptXsZ7v+JuHslBHzAKhBu9ryEM+GdGlypW4VMFhHVciBfOBYKbGasNe
KD91HmZ9L3k2HLse8LI5bCitfZf041dmiBH3ruXtNl5qaN8ZmiE/p5MslzgYu9p5wMZSi8JbPqCK
xdabfSouolrQKMybO72S++H4oUsxGWQPa1rprUghe3aC/MYTCZwvoDGRK/+WpyKXyEbBJ3ZZ9Y5I
mpUiiemG6YZrhwtRm5xJXK57IMKvqlpktiOeXv04tuNs9qQxPk8oADR8+oO4qKAxzi16QjfpvjC+
6GWwdMzQIp6TvhZw7MQZIAe/J3YgQF2phs12rAzhaU4x3c2fUOpnEF+SoUZnNAZ3LO90ZbgjmZVu
/DOX5B/N4xM5FlukW9pgSDBfvrisLDr6+l5IbyNR81IbYkRh+cp+a+2eKRMI/2jyCvPps8lFBf/9
oKBZM3fgV7XXkE+GuA/9GWd3zz2BwdRRK3Om7LEbe8QcdKjxAkzhFDIYZINsywVickjsts41hP+b
XLaDY61eWNqVpeC7EBSFTRhP+oxXRFCH3Bi3PVSETHIo1DK69upfOjUla7/er5xSZwWiPzRMrvnk
rXfbxpusNXVScZorWOuHkN99RjTly0Op0mYQWf5B4UynBOCelszpHVVPGqW48lYL9YIaPiGEXIds
IVRfWoAk4zkdKdFGehNRiMP8cEfKZ3piSWdn1+/pEkd3+5Jys7VkO0xoKSw+pqnLr9t5rXsGQKFx
UsIz30f0RjIistHbV4vTcPHuNLjwohJb98pR9RCOdrl99eepGorflFhF8qxrlHAo5ugSSUbCKrry
smnHyy2XeqWjB+zhD2ocWR21KBYM8knciP3PCkjfbWkWWA5Ift4qneFeJEUwB90firno1fAO2kxX
Rdm0ohnTjvP9SGkD0dFNrdfe/I2Whelde5fk2ECyNT96+o5ENmAXtqlXuyLfWNe7nkabItn0vu3k
bd3yh8pG3UuRas1Xg81Gjp2EE0bru3yYpql6dPtge87yPRgVMLuL4cjXVY9ROEN2xZJ82SKfzrVl
Bz4nj7Anp89+WXdRjJdOrtvXWtWqbMNvIriaO89njl1XL3c2xFiKFlwHV2UyXsAVFDfI2UUbyo4g
cDG+Bm5XlPKi7jekd2LKqId2eeqG7tb9tIF9RcRXYCsRy+col2lT1yANlx3uv253aBE2exeKWui7
Jtnpdr+NxllMUIuw5C8XXfTyHS511QkFLR6l0hz4W1imMzDQEUWgK70EETH5VryCziTvWkHe0K9g
ES4MppJrQTMqp6Dl0aCuwIcEIkQbY4wS2mvZF1EQNN9L8YfHtq0dMaFXtItiBICsIcvoMZfVpIG9
BTlKGBMPXs3gXzezrCYEs3+Nl6vxPzn+t0Yr3wKgC8x49TOGseZiySfLcsoau+FEl2qMSA1KGOOv
AEipWJu/AL94SN7eScSeTtAtD/0Nb7eXWgStBp8XGjajqHhC4bPs/q/KemF8y7a49+2VHAYdJniY
Y7Xg+m631XaQZisEo5uKQIAd9nq8FBj6zyT5jlgshZ0c6SgKNjLjYVlxm8rQpWHPsN5s51Ygqk74
ieHS1/5h3Fe9lxbVzwLJDeM/QeRQ4c1dNUIrsp6rmCYLbKB9rOaVCPWJ+XGvH5xRhY4YfRM2rf4n
6sM6hn+2RHRwI/tJJEuRGfsjhzcjPulB1BuxGpoMffx1lTQZfwHI9viLM7XbwEu++V3g2epgB507
jkeXM73lHTbR6vQMiqXPd7n3lmn7/YhH+NX8FRijrDu7+dM0ZQ55pVPJgAOdzb1PKpqlweMQ+Qgb
M3zbK/lal4EsPQ4DO5jHdsRE8wybg0EnD1aMpCWa+DgsBYmijkWGuWEYY1PwBUR6StMW3unTlaj6
m5nK9KJAR3t126Kps0IjxcvyTDg6N96aaD1LTXrfd3A8iZkXYYSyRGrJrboTPLhWF6Dn1klOCHo2
MjBqfHJ1WuiM0fKmswcNFoFAShxnl8VNF0AgbWJOJyoq8Wf7LSZzDcmcGCDSG/3m3+eO3pnZW9n0
3b9BWx3KOsYQMoAfTfwtOfk9DWqvvnoPtvr7n8EuRMhxEuaZ5OXj3TCrPBBl7XwFORwvTUY3agr/
eYINDZ2LiPSL9v9RrY0KivLktnRoQBdVSTzqJESKeCbZwCeJMOMl4C+01mc/ClNkjiJYbI8AqdoV
fOlLZUnj40r3re6KGqCTksF56jp62j8fevu+vT6T0N8Uzb04NiHOvFFmipiqfqEQUViqkWkWSIvA
SSKO07XOin7E0YdJwQF7tgN56P43eJU2aHjxaroTZ4APg8ej/wlfQEdEldcABM0tcnaKOesSLcdx
BE6POn5zupRCIfj/NLaiyxGnwCfsTNGpNmO1wxeuZjKVVvaRcx9SMeWzbz43HjQQiq7kuewlMofn
7PIwiEBaxvlYT/wqCOJB4nDlkCA2yTrwgnUu8bDUTieN4OOfQaA78sBP2nH6xYduRDFuXZl76fVV
RAmjlP4U7K3cerkXgJhT0ggztXY+l+QkhKOTkfwWWNsXbDkr61MAn7ExW9aKDGYgZgIP/gMde8C2
2FxjhmdPprw6aZ6O1SoIRdlqmSLsWDyoybD4TtPrKnRk9237JD2e4n6JEE/rZMJaKvRWJ8TsyuLu
wiQYPZ1PiBnlHcWSzj8JFMqw5OaobySS5q3Ettu4POARePKQ3VmSywP2p1vXgTwQpveN4KfVTfEE
dqei15oYgEP7SDKQynmJ+kVjvzaK8DcpaVvQAMGt1e9V6wR68vxoZ0Skyt7cXxwgwsucQYj+ZUb7
a/lOMfp2pIQw4k7EXMY9OkD/Lj8+o86qMcgiDtjIjswFjqhoneW2b54ZBnv0bKfNfkZdCCEf+sDB
ElrPhKOb6ws16HkTp3c4oDeijR+q5iAsd8s09wDGtcDIoS3sLDDLBFLGDDknnijxbb47ogv2mw+r
wt4SkdZpq6D0PQ26PxjjJFoRXrSTevr4O8m23DLYpTT+7J9fNE49Qb0z0LuP6dF/t4gO2HRmFHJ2
zsg+9Jtzb93TNnA8fxUQtL9MbQHHphRBEQLxFEDP2hguTiZiWzz90992g8W2/Cc0kQV6jwRfY+GC
qtzTpK4Fwy8/qyxSMh23uIGXsVtIB+02qBQj8yuoi6ql7TMeVrwcfUZFT+dDsk6d15Kdzj0RYDFL
Efk+KgHf1I8l9fYALVK0q3tsM5mJJlMrUTpUITpc02PPxF2H453B4CgbUJ0Zqq3dDro1NEGLIMQN
9DHVGQkF5GQY0Cod9xjUdCmleQwFnjGEw0UB0Beu1Ad0l/skYTatpQhUDAg09YFCY+XssnhUhFgF
28XROC44JSoFr3uEH6r7/0weaWgTcobssgXidEYY7aLeDsENoTFUk5k9MxBwrNIedMRBdL21g3gH
0GqYWsML2sq+ym0wcOpx3Nyt54Vbv48Rc7aeQITpKv8paN9mGz3zI3Ujl/3U4w4Q2geRLSc+8Fk+
hocVv9dRfDUpyysExXw4xu81fut6o55UvkHbW0MNqnNzxCMZIy8iMTqCdFPgLIBcQRSEZzIDSw0/
NV1DA25o49R/KX0le33G+U1jFQfcSGjTKbOSoOZoW0/SsNp77uSUi/ExRGCvb3s7VxHQUKvxrMFt
Pxcb6eRb5/g1zRJtd4UxzJZp+1IXOS8nb3saUk9vMjdSLD+0yW9IXDstTGGT1YVvMO7/Iym6dUXO
SwO2amujJz3yeKAPvBay0XIEGJ9dvNwqOXm1BxWI9/YLsnReyBZbETTqsEXJx6UPnHkS01UrDXc3
vx8AA2SXy0jMWUclUKj2ftA4aHYjjN3nAjBLTGk9q1sUCegzzTsJ3fQec3KJj1DfS2/zdSYjLixr
/og6k86pUuV0LlcXdTkI1xIJDrzPqROkjTi+mWhfgeIcFjfJLfDGKPD/8vdCDRYCREOiQp/vWJB4
xIiICL8QH9tddHg4WZioZETv+GMIQXCyW4jPJdPG3QJHl7JsUea8tbjge/pTSSj2NLHaBJZpQepO
oO6C1biF7de+zQmwD5qX/BCh1ojRKaa1HYA4lGYw7vbzKlAUzRGjNGw+0WrUyTuo2N+Rm+h/6bDi
KLkShDrZucZmcW7wYxb4RkJKarFcGNtFhWHjBmf4GRQYEvrKrtE1beu2aBcbdGxFmyXuLtuu/pf5
h+UliVWQ1whs5go/Sd2r/iRQpiAfASaJa20iGS/P9/QhLjdkYbh7jAFqpxm8AAd9zUFwSll0RUP/
RD/dv1o1ad0t8UGBZsgMOn1ebw6YJwcTKt/qlq26oLtWgiblLksDGqTu89iDilDlHvSkT7LJR2Zg
DyIEzTO+k7PR67sdqxAd8yO+yj7uz9VsbyqxnbODnolW7+n9ayniRZ30HTA4zu01+hmtCrNbA1pO
RpxSp9cHVIAHn5f+69LEvC3PtGuWQcc2LNvyM5WxLZENlp1c+S2HrvqvPhUk8SaL2j2axPFXff3H
WHVW5RnLU79KnEyDHPS8wxAWKzCbnJlYUtYCJE/CabgwYkvPtFrC7CvTc/uA1uxSJPZZLJ2tsNza
B86kE6euLIXF4uL9RlVVWVAIqyJtnosqeo/8TuLiQjKSz7UXYRWeFm1+bjVk25M5FKKss4yhA8R1
rZnGZ4z4tEi09f6GdcB66SugULm6pKo8PaGwQzuZXGF6kBBy8dYsThuiCJeXPBe3f46pUh+OUnoS
LkJ9NDL6dOQYUv51V7rG2j4Vl/21q7vRYT0lHqtDqAHiA+YpKzdjNIHgAq3ytSnEh+FA2W61ryL4
1qv/KB+rsirfSndIb05qlFK145Ry4BP6FMD0bhF4XEpbGDHIwbCj3uYkLRDoWPD3uvsJLMIN0gYf
CsSnnIenIe6ig4u4Cds9KEqVnUFK8HsDRa14plxkiuzcTALAUIuaMHRmCsPk+npdpMxdtE+TI8e9
Ab0eA2pBZkMTlnK1tMLsHl78qDYHiAWlj0rbbg7Vem3U3d/WNVcoj7fwl4FnnTSxKOYORHc1DQg7
ydcEJDCwnIs88yDs1/sPMlp6G2W/d78g7zEog0xEbCI2T0oEl6y3/GGLwq0Z+zL5/VxRpLhXsGIp
LIsyfkAV55He42pCEfHuPZ0T07F5yPGcMH/CNr3l4pJU25p4DZHaZW3XtsI5lzkOAaxeSTO/kkD4
iya5DCE772gpLwaLMEMSvPsjucM3xMji5Np27mEyczhsJfFQOdyGaeLI8h9P37qLp+OaCg5OnuX6
3rpDVK3zMBSoc5Qn+OVB9cJl3Vr6LGE6y4yumKDG/Uwit+OFbc36ohKqFBNOuTNLgd6Ob1v45WXG
Rf764ZnyytbbtF4fKcQ+ZX2aepas3tg6parqoju5yL9YqIa/PnL56whYbRCZJLXQndF0LdIhL3w6
xDzJbOyNiZ1yDK8C/SuLsEdG9KQGVEvODHrxlMkm3LUYMBEJtILEo0pXzHwAOo+UApNwcaczE5SE
3JVluXI25J1n14ZTK6BgYy9hHjs1IDbpbUBKQ3kbJ/f0nw1eW6m3Kl+SOIRJ516ZxwYYkQap1ciU
Lj/ewwgWVYojI4i/OuM29Eo6TTQi1bU8gEAt4vVBq+QA8QMeXoar4yfZww4xKR0OQmHJgJl8cD7O
InBXAjEzNw24jGjMILfvWKs9On4wcqgof7w7/G03sCu0EOLeGz18uoWtiLn5fxW5NlqcgNRMgk67
QAyyQm10SGlLXjwt5R7NkKAYBK9RTTjl2+pVl7fO7Ta+3vKoOblHrh4Gy6D+izjf4rTfpaH3obkp
zTtcIfwK3iac2qOB+P+MSnWZC7Vv+ZnCTE1zXi8O+b6vDPDNgd9w1P9Qo1hvBUaVgVSwwM5OE9Gd
L1E8FnwotNA3m0Wdt3SZ2iqgqYv/pU38HGBOp6FaZYua2ncPsQTsexAvzX56cdeAxFFZxHWsx17U
evQlHCUsG8668+XFcW8UiNy/0sklvoRyK+k46Yc/XS+M7I73/gLJbEmfcmMWUv2eZFHFpB6fOppI
IyFHWqhM4sgIyl2Lpr42vdMa75nPUHx6HeMFVoGy9eG8cjo/R/hplJL2JJ95tn7OQtWgq0lijce4
jny94/1ILTa/j8TgdUIYiLCOkf0iqGgBrDo6WQhhwanFsyQZ6HpJKyDw4yyAWTQt7IRR0reBSC97
Lsk6oZ6uhCM9sn0RckYsAvkDgHyqRNSUrE5Ff3JBPI0gmSW+JsgfhpbSyT2mujOLbyuPocCFiYkh
JHkR3NjZi4ENWkPd9CH2ywQEbKguJCVulI/FIQgKy0Y3AUpSEQs3fiPGcDWW6AqiQsUpQ7iWqZh0
v96khai0tC9qxmiWTA9HhejM8Yx7PR3qATI+PiWP5eFbjVPEV78s8ZcaNdEtsq2g1etWJjjNKY2m
GrFvbsgWFBBxzaYiMe/LxjW4ulExE4U3BpfnrXfxcvNmYao+s439IPxa5F+h9PmSScps5fWJcGd7
Db6RFVYGUBidJ7viOzWUF3A/jMFmakfmGCgM975aYyV1r4uZRDBCeRmi/pRv13NR1zW64e9DDueh
lWYTY2zNr05VVqsb3BkAnSz6TO3rNyxDpyXL8OpMi40BkOpqp4+8p+JjcsFB1GNQ6n2yQ5BkkADO
l8urHe1Wdlck2Aq6b/baTfBtb2AHfNVOeu1SeVoKyrYOnhAQ9rFyplJbW9rWRCtpr4CJ7FLIP1l0
S+6Q4p861mUGYoP/GlAztPVjiOgQp3nvprKlj3NS7fDNm6lBbZdswDaeCrjqkwpVnc1+LbpjZu8H
pCBskjxYM/fZJEVBGMgaqKRb4bhRpc1e3PWrgGAB/8Bqd39BTGvnkoSTkkGpHo/3HxV/dylncsC0
vlgeLpu+p6iznnHsdcyFe0uowfw5zJ+K+1JQa0Ev1xmDuRPrHI6B5rYwj2/KfoNbxQc9p8wa84Dn
gfUgXrd9pMp5LFGeRyVpg9NOHxF4mKJPPSrWnVfLIVMdIebzD/5+SxE4filX0ulL9VqxCf+VBgGK
4eRHugzqhO+b9LVZT5olKawgeqhEKV0hwfKUwAFUIPr3DNg5CT57SW4rVItIFpvBQYj0PcXqiVgp
PMSXDpJVfHaCuSqJFhrtdjDLq6kydD1q9pOomWG2M7h9q1AI39cu54dz+zBKGGBy4UtFnbO5JZ5g
npidGJaEzN3+Ida5ASmab3QXdtAqNCWCNLbrF7rzDAaa1gyfipr/5H6KcPTDqnPvglD9JOWvoM6a
pJ1uLLj5EpczFHWcwqzHtvBfp+rB+8ess6dQuQjXlmXm82q+l8LprNk/L4bgOeV6ALjnH/IpPo4p
j2E7sd6lcgr8uEU0wFdxxlEP/+jZrz9eDE8LKrOjt2JasPVi5Qt+HcgpO9YWNFbXbiwonVubn4CY
ZNxl5jCrqYnDoLANm1ss4GY3K2F/onpyveAzsfF6VOIkLUtvUBL2gORWexpvOo/SPh7ntWuXjVuw
qRg6iD9PnllowEIG5a3rYFyNrH1b2jc0DPtThbg18vk3pVc/MjajKjzRhbqbJ06qyRvt7ef7mXJY
pIgAAXBVoYLjglVfyvk7AoL/oEzEYvu4j1USXE6EdXhohUvyLltauSkJxaGRY3UKw2oNduSVRLE4
D3tl4/K1uWga9SluTRdCSdTgBwQDG7/QgrzxuABcxkQCxAcyqZIjk8F9nxZg+mH3arApKhtbPHys
E1nED7fD20Epv4WY7u3TiqAd3wZ6neOzBL6sFl01cfQWJK59K84xRFEtJpjfgAVLb/FljcBjShlf
8wG9P1SWjwoKEbhPlR59ZesYvPFY6aaquCwje5rhfj938fOjN0iG7V7ovGWlbyZjmgD4WMlpzluV
hFk1Fs9FX1kPwFNH1oJfUw1wVTUWXcbO4LYD/ofb8w6g//bcmYU/BG65tPfGhFxQbtTrTTbqDD1t
UX9Z9Hrpy5f2wHCyKWKhl4ly+p5QwpTfjAXKbnKBSCJuHXObOJDOUMdEaWUd0AKezxl1gGdT7F/t
uG2/1hh6M85AtTvONL1yCl7rSQyN0KWxrzWRVjiZiF8C4dScFCvKA7Vb3X8ImS1XhoNL0drXukwh
SK6pQZZsoMeo/G4h//ZEkUKQvKRK7diEtxIpiByEPPyo0RoSSLoIrcsA1JWaZi2yLFcsIyz9fZWv
hYIWHV4Az/xFP2Nw5P/tdKsTLVrgRNiVUpGeK7pBQwUH70mmhZQZhvft/tAlQAP+A0pSVI3lMHKf
wscrGecVMTXWi1KCRO/boV92RTTAT1O1v3H9rZW3+VjVucB5Rh0Pv8whwjj8lryQovuVPeam8x9a
lHuRew/xRUq1pw3KuRShoKvNrXnE+5t/QbnMsK6OSv4cR1CacM/WmYcJsBVrdn1fPZ5xMsKj4fHL
L3FpE26tqly8f6QJlZ/NU/f5EJ3p3ieqDPwGfaSAVb/qtcmu6UBvaIWYnExZiUxWzZ553f1E5APe
SrkoQXNBpNoU6hDurkbzS3hZrhoPZ3ZacTNaJTwsYXY2cGJhjyPCU1hbM73PnhVEfgaJZ0vWzALW
G3RnvZKCSAX7lT75xOcLxbFr6MCcBa9ITLyjUmAc8imR/QuQpFQblhpkczkHGf+WwEBuGOq6H/AW
uERTcs1QX6Fj8Vo7E+5wM4MZCjQJToulVB6LGsPFnC/8ZN6Sc4R79XBy4HlRSb1UzHUkuqD8iGiB
AOJQD6gy7O2GWdoPJPYDRex+k+fn+OHr6jdyFWejyhTsq3FPAOjF/oIFH4kPw9LSy+wzqLOvqYfI
sF8GuasGj0drxNhtoT6aYC0mzNipo4OnJEpRz1gnHHUVouLNOmcH1QGPku/TRMOdvtpTjES6cOhF
JAEmm+7cUOMLLP23JEFwJ4XI6y+QZtYTNyWGQLZaGHoAuTFBFrlTf9utTRaQy7cmjQZI7YqbyzN2
xRyHYqgmit7Kkb9UP+E/HyUYjJtocPV4iSwIbPME7WEnwYKWlGLjjOJfX6B0JQdQ1t+fQ/+GGrQ8
wNxQe1SJQR/gkaJAtdcDGj8Okrll4jp1xv4KAWjJ9/DTqB10jfRFtcQOH2uhCrCKJAADqWln9ZpX
HtqwWld3khLMZC9wYSruhswq90Y2xyj7/ZDMUazZgdsyOvgHZEe+PE0g2qQHhRVt+zBtZuLf29VX
umbTC3BujN94uil7dAp4tCMbzI9yvU8x5/PUyTIBXbyYwqh63Vx5vzjMG8qSHa3W2TDPnHFITukL
4oBLX1tAbjV5jRwDc6dJdajzJjARCnjs0OnKHXzvczI6Lu8etWH9VgD7ylmcuziPlXtTgXRF3wQu
QrBeqpL24SQ3AW5ysJ5hhWVWWhnKRGO5soQtHu527ZqJSrsXe9iwvXu50Y1oYypSNw13xRM/Riec
/IvcxxG9VY7EsL6V0HPzKfzTQ2ufUBMiLthHtqCG5almhRBG0JNkWOZseEXZnExZjD4FuUHoK70C
OyJZfa+w1rmacOSDD7kXwbSGgFBIjGPmkjsWxL8avJNZt9gNlPxATQe1WzVyf9yvtCGzPWpwNbW/
Z/1NsOIEdAkhJCCzklO0lbcgRHxbSz9LjYyJK8YzOi4SpDp1bhXRI1/+r6ilL1V3BhL11T/6u23o
ygttt+671dXSO6bL8jRPp/KJ1BTv8mS+okX8n1Q1nhpmm0yjibSwnX2Q12KjWsLvYeV0EIPLOVGK
SSBeyDkf7O6U9UxqmCipo4/kptCJx2A60Bq1rQMj+AS4vMM3nE4rdnbFC9MVq7XVQNF/3t33xAxb
aAg9F1mNAQEREj3Q3I8aWE+Aaw7+kHYk9fGlqMvFG2E5osD5IG4Kq9fOdP7hcHI9yz4HLb1DexJu
//bwJlUNWCSjz10ssEeqwV0P6gRRbTSSvlJcWyN1eTGb5ZoHSOjfAvfn6KVNsbOc6VTrJsEZdAuR
LgEliKzASoBCQN8j/T+ld6KeN7p/0UTTssrHnEJ+HyGUqRv0I+XcHJEkfGgC6+WNJGKGiWKYP0n3
NkP/f4RvavILA8xRwC1PFd/WibuWFTFsRHXCOETX6Na9iMZu0I8Ig7t2Siz+lkDIIkUI928wLNNR
YdTFwyzke9WXkdVNbMlBXh0BpNdO/RP0mljGVc3dNjAbHvZxIxb+mSubYEqA2VShvJZueX1k8JwK
sVx4Tsr232GNID/9S5KwAZMO7mIXrDJ8OMx0TQKU3KYO0a+8GA6+OuMZb8sup8sQ7h/UvKVW025L
GDgo+/EmtCIC1RoF7jgJFcFDPTg9GOyZrRkQlJB4dDGeAEF/JCsYA3lTSzDvbHwQfda7eXloeAZT
Yn4MQg5axm0/h2z/XfpNtPJr8vMxH+eMms7uLyjteA7L4sbtBVIagnHzAAVhLVIFYiWQrwJrt3it
CjUhDkfuxDAgPCm/Q4hiqQqBRFipk9DSdrXvprVhs0fhfF5D4i2STNWen8VQRGH+PAUT1vYQJ4gf
prmALA5PWJQrYNdWMBV+e5Dv1KFmM6cygP9B4GB5JfR5OdIVElh/9Nq8vrgSGXbsQLzrDc/p9x7Z
9pwwe5M2m4+RKfvFK/IGv3Os0IKTw63E4Rkz6plOGwPmp+OWoqb4X1N4fwDtOGSxx6z3eY3VOL/j
7xZgUHPOuE57Bedblj2l7KC2eVoK+cvysY64KAjuLfyUo2gHQsNpn3rPyqoAJzZR6z+RF9iymkpr
1X06C/YCgszfEF55IVZ2a4iEw6C51SZ5iq6c+0fADR322qJnkRTkcuj1WnevW/URfNuboivrFO6a
WxzqcONOCYgNbZfqCTO9nO9f0goMCzC1xhB+Q+SxTdkzScwADzHcvjhchEC5vSqqjHU8bEts05Dq
QxymHANayIPnE4IgvUUnDSzsYsd1LXLn6iS63cqObg94kH2nZ72mnvGeKZYaO/8KP9jjB1RewEmm
GK6ZcNun6j8/trp3fculss9cKZb6mbKy71hI55YCNI39dJTQ1yR0d65Bl/YLFtzALPW4XQuRXM/I
6wStpnCNyW49ZhDZCJBFrYYaj033RtHlD4t2vnk4f6DS5j5H4p4KWCdErvjWnV+vEklAtYjzxQsP
lGoWsrCFgKNrLcRMRUQSA6qWazu9tVNeGosfJAc6ivyjbuthaajRIW6t2E7GsQfcXAA6Huhaj2ki
YQKgvnnakMZidl+GBZCqOijR0qSxqI3fk0GsNQu+NCkAwVDd3BGEmhg8jhHngHtSWEWe2S67S1Ke
Kr6b1d33ScoPeYqFfzjto+/89hPw5pvF8jB32fVdwqjIizCdhKs5ponsaLpP1QxBP5PqugqFgtOi
uSj1unEDgPP4lx5jrgwM4dMGKJRWV0NXLT6dXCqZO43F9pkTYrvN7rtf8gu8pCkj8+TdaR2PwHBP
+Q5JVBOervgC8inznfaVHnSaFEJfruNwKurBLK4XKCnRivYs+BhtcYWmpjXOjDUGWbXDRQIRThvC
/iJCGnQR+TBaEMfeOzpi/E5n/8DgI0K3I4mvwE14NrzsrMuMcC1HAnbeIWpitdNS6hTbHOhy9CPS
JPGTT5Jr6E+092WqUrYFFazbMjNIs3tDK0laq0MbTvXXlQqR1W7ml6fS7SWtdtqJf1aCFoTvYs7P
GqBQ+AxkWgIiKQpBtLcLCkaIKkp/lm2bVoDHSZssSUp3TH9YVM4qoHFKu3Ec5ue8i3W33W77FHSX
Lh8XgVSURzdKWZSTfyn9F9eywE4Wt9YgyFJhzUv4Z8LmGqkgRIAY/5PgBu/0rz3zVWb6fll10Yu9
QL2gePstAmAgpkF2rJJbK9012jRDTJHcvP3oWlXzf71TmS74v61ILsQ1EUQU0XDBcTZSC+A5XYkf
PnsNElhU1/S/BTZqLmW/fXodyYGd3OJm0XlAvJEIX35bDYoPOzIlt7+H/OoAngmj9HcbTFW3znrx
rhQsi40YhKQ3IrKdXkkNfRlCG3r40XOvRdcSO+PeARI0PcXbvHHtEB6xJ/l6lhJOpJSZCNsfTPyF
86Vhb40F9vmHuX6iC3xfpo8xu+8GibH2zy6f+3EqVFFiTWVBuCzAfKGV+hBVMYKjW1Zeth9rlpi/
ZJyd18eLfzNGPmdelFNn2irUVRqmKyQ4Y8GGPH4O7jKlvDpOUwWPu85gIMK9yqT5NIhPSCC/gC6y
iz+TRlYoyKTcS3mF7l6oRB3dVC9PKROLAYQmXt52VbneUfvKit7yJVmaysc1obx/ocT3gCRCmypw
7HgoeAFfaa9P8Zm1Lop/hO4Dm9e51X9zMJKstuvwkG2npym+CHEu90ZEOEOTKqMV5abhfRFCvVMl
a7nAkLKttfebTm+i1CQHZMXFHKCZdbiWqiyeO7T5Hn44I8Br4JWTCipza/W5kAHaxWAhs2v7SV3V
09C/2beCIZuipcYzJsaURfd9UegYo6FZzCMS9CyVxupeq8jaHDXA0JofEdHvL/AFQZTAsJ+wOhyL
o1fd1ARmNyfEFCH8HN49VAUwNaLp5fZt/Ccr/5RrfxcwgjUbFcQCAT6giYtUA5IFqH+Hz9gTkIFs
InHsiamyEyNba6DifzB9+F+d3DSeOlBnc3zavXm+rUOYe6Gu3i+dQ/82nZRuSCmuvy1T++NOE2qR
xb2aQb+dZROQQOr62kVQEJi7SgvkmHA6+ttugFwBy3zoLyzJVHbc8ekeA769EME1M92bbbxszsA9
taip1e+QOf9LHTM5IeG36NsdrSTHj/amy29SJV8KaGDvtVMLNqAeyfIv0A3ymVho8Qj3RakeawEU
DS3dVRg5QWoUulkgEt2geHp/lzV0ZRSJRylXQOkqeHE0nrZOSQabE4JlxXmTWZ52ZNKylwk5CZwM
cd1CLwYTBoZBFb5feSaiFK1TJjThl8+JRq+fFGloR/iLojTaLBH/n5o5MtMhWRfHtirUQ3O41pOR
aj5VsUQm34LckTwKluOaeiktFKEhgskg27JMqGxA8bRtGLWgqo92Pyk13IuEf4laURfNpoFP2EyQ
eQYsnkGRf/JkJiXkTPE8vftD5NSCl7GsYYS80UGtIDovHMwKS5wSe2QIf+4zrGjg8tDbPIsrE8ld
EugbdhvSisBHyX8nVOqrqOMdzOJ9HYGOUvydwjACDc09o+6ivgbn6FuTmlhlHeIWGRNGh31EhFBP
/fxQ9aXtWpe51bI19ymgHTC6Z2PUhH0T9BoHQO/KEOol5q019SbBpNKse0lP0OiKlXYlnZjKDED4
tFn5zvLE83qLVMdi/tHmkJRFV3QQQC2OvruMX8x/cx+/Ya9w1gguZd6MOjBXYz/Cpc/rlpL7A3B5
dSKPUS0rEyiHtgQFSRa4TSle2L/2DRlSBY2QUQnxUEZAtTdLJVSxca/wh7+j7gMqEPKRrmweV8+t
2IJRNMv3Adln9a4z4ng1L1LV2zdWR4wL2EAm8X9867n2T7dFfBE4OWqhheAHt8I98beo5tEOr68w
WSgIMB+oWXosYfSJeysdxnP6hMv3BWqPO/iujTwV8gDPPNykEMOwHWONyjvTltGd85DoWzEeh34U
sQu5bUEyQ1EuWinEcKTDINJ7Twjd79kxaXd48dOEk1MnWMABwoKy1Fj+gN7YJXRuNbSLE8rGLS51
oA2ctwOSzZ8/Y1GlfC/TNxVSovtxhLrKE82y0fOK8hIPIfysK57Ok3JCamAJMkcC/zR2HQ5zFsj/
jTvJeSkilyl9QR2JB6iz39XCG+wlvg8HiFnSYPWjAJCnFTnxah+SN2ERBLk01sqDuyOr/KW5aHd1
9JYXsAoqugErYK2I1LIhvFc9x0sXGZ+zRY/5NOo3D89mP+Af1cpcQUSWntdoJulZxIEDRjH+sC6I
HMJx3Gj9u/EyKMJOc6Z3TirLVc671YDGjHn1Iz8zkesrNH0o3eBr3GCcJTAUQVmtNILW7OKdxcyk
KbtEe20O9Y9ZapX0PfT67Cg5F2co2FCmJkAlcOtMxuU+kOk49bJxn+d7fmFMiNjCK2gmLKVYwrl/
IJphpkEI2Vq/xELf5jxaNnGovsRPLxPQEEUrbPTqNefh/x3bkIZkMmIbI4vtEXS9FGwTI5qakBUU
gWUYnsiSB5BTMW4mWms+n/6e53//F8q1JltPxozbKyrMysRiIxfD9gAjrXld7EsGhqiRUrusI2sr
mlWKXopFta4zzpw77oYnWsR70LXEp+Djpyw/yD7MIOqk+NHax+xuCOfNZW8eLXrF24Mkx2EP9vuZ
BNfpNpgSbIQNZcAsI7SeI7ffY3uPWGrXIxeFkAstL3tNrbMXits+kUVzlLG7q370qQL9RXO+zM/w
9/tu6BBdQJ5Gnurs3U1Yt9yHnBnQHf7p5/MpXbQTRTB5Ov/MPHQbnEkuJ+oMtwFJ8pY9mqI+Et1h
1J3OcXTA4R6Hk+V4ePhGwJzAjKGA/RgwhDDL1vabDYc7eqv3buFcQ4H/hEsyV0jw3VtJw1xwdIlf
57BOV2YuBxJrH+rBNhsOACAziswXf+qFn73cB5jIInPvaQo/wSzJEv0q0NndfuDneVPLl7ewDgcm
cPS2bnAfEHnOikMX4EuiEzYStaUqrL/wMPigLarBieIT6BPlrMG8pmOeoqm8wDWiSpFxvsl1UKvn
mxRKMIWvMQbJ3s4KVDw8pegXgFTSY2zWVxRScBF2Zxtn4TFkiTYXbkZN5vqtAsw2ufTpEtxJ14nU
uaPnfXIS1ynaKZL2PgaAdxY/YFhSZHOCsro4JDE6urjv9vFeLFrRCjqjUcJpyoVf9uyWQsdxXIl6
Q+0ZwNuScGpvCLSHKF0RLZTSUonwCwQVF3TU0jV2snU+TxrjmKv8jbVpKVjHHd6sZ6+xMJ/L2wFw
dY8SORfSVGkkNFmrwqmsSWbVsOkKPn+ACnniYSh+S+L9xLYg/Q/8XvGYi+ppL9U15+5TTQkUenUs
pVE+/wJ4nSEhIabKN9p6NjBw/UPZX2KCQ62OsYjT+hKCfi6lC7xKJgOIvn/JmapxgQzSw71UIkF0
v/wRr6jDQ2O81Ne/HstEQxX0ctmXM9feqO9bmASUTLMnobZc0HOgAar15g34lR9OSbRR3DWJlSOQ
FEoSrfIRJaBgof7EtoM0Y6TjJo/Nz3GNHttIcwc/xG62d4UPXSp4vWVgVv16+Ho0KvLIDOM9wsnI
mtEe9ZSwIWWa93GzdDOnoQWozC3IataqgCT3GtEuRoUykv72v9mUNaLkWGk/1sRvLW3upErJ0Ef1
H9KnQuDhrhuQs55JgSqZCdxiJF2rONWdbQ+Ss1P8wSF0B4p3gToT9LXTnNLdiyPq3DNYhblEr8e4
V+pXTf3mNnoWhjYKsa9nX9u+UTOJ70Xo822JOzPs4yjdVzE8VSKkybTOHQJWcgii1Kurhnh0uGPM
EzFYijhMWZ7neF1cFDe9TIE6wsuO6e/2avHa/9vrBBRJfSMjxU4mjTvbqhRozX4MRpPpRm78FDuR
79SzvlyQ0o4blawQLmql9ZI35/aQfpxqe9uzq6OjY+5Y4BebteA59cQvCvm9r1RhUZJpKhSzHt3K
Rt7r1wvm30992sDkRzZiJRpoxq9HzhifaoyU1vhiLvsISL3H1wLSSOaPLpW0EA9YW8MX2N1nRqGB
GDIEgQoa+k70mxdpBnVfQIL8GHLS289Ti1cJkAw0qOTgm0sUYdr3IIsD158lJnkdiNwqbwBr27OI
w1ByrC3FiZXA2txwfnlJqQMCwIRxUkD9ykPCKcS3tee9kyVoigsUm4zwxkKVplqkDZVn92D+dmst
i8oI8R8GxBf+sGG45O3NYsZk3razB9dYADRLTyNuAreRSFXGBsj+uQkMksrq3xD4cn6U9KFWCk0Y
p8Ov+kWmBRh4IQUgumI2NA4qA0IQUakbnuesZxE4UyT7HHdmVDDoXVgAUTV/jZLYHTIrKTKFI39F
DbIO45iMtedGck/0O6j5niG9/ITqzoQtNqpkIdMJsEzC2OqRcB8DcaUyLr1q6ZxOBecCbclmpElX
7RZM+7uJqqJmpJ4F5Psj0od741+uZuY9X3BuuyQrR4vUjoFnph8piWbgSI4o0hk2d3nkM5p3Z6ho
kbwjBaTXUlIiM6rK/2aB1k3IX04IfYifY0AdJhlOp0XQPcWl3Gpan0UYjkpKjNNLHR1n+NZ3lgFg
VFNx1MfugasVGjj0rWW71PJnCa/U6sdN2KHibsyQkQz34l6wBPMkHDpzcXCSUJad/Ajdt+awffz8
ZJwkklYchM9V26fm7iFx+z1Py5TitePMqnI7G9kKR3c5dou9lVNiWTKBMzf45QJaR90OqqFYElWG
JLDQoOm/qNZkmen/N9QrzlwFuzFI+NnxN4QMGnsggaA0GheF6avA/hbSTm/Ik10ysJ+nYNlsPli0
1aY3nE7nsQvrZIeeqABtRm+mn0f0UzNMKdi8/5Ibv0/+kb4o13x4oZIux4rA1Spik7YDTNnJLu4E
Au35WvJRK+EMLdqAg2HxSL3y1d2ZgMI42S4LKE420PdN8GIRv4lMebS5T1h2JkpmqoWukBa4CPz7
6OZPpwgsNciAIfZIliPbyZuLMrCpiIy398ZCpdyrDcTbRaOiQ64av0K5C2rLCmUJ3SchqTgDrV45
6LSRgohVwRmVIQ6Y+YlwdKUd9Oxi6SrOhbVZtgZEdOdDMPtWh4aofOqPzbx2UIevHSjW7g0HTKzL
PjJpxB94O62R8jMilgVOAus/BysyYxnNbhZf5/Xrpih2v9gSyiKdAHLgRM1A9rOxR/zfe4+/AbNN
unU7gqyoLHkCat0Khm3Y8eI03RQtgFTas958eG3SQsiq02eWr0W0jW83GGMx12AaTVn5rs40fbgm
+NKOOWr1MYdt4+kgj79bXlHUNknzcRFhKzT737CBHE0vqFGtU8f9GKz2CTBcC1xI5lBknqYtX+qe
EbBrpGKfD9wAcRqJAn0mEKxU39vV0z8ZCdF1/RB199okE7NVsZ5EX5eHoL4ZS+rs417d+nA1J40h
USRTKuSPUOB5M13gWDnUbasHBHh29JuzRUIZtttN4XV6/wisCB3fJBG2IdWgbosI+MBJjbVKuQ3E
lp5gLwuLMLtImV7S9TASFQOa9VmNrPClReSeYsj2I2HTAvdb3oLwJhZ8JrXTOgcGwMC1PT6Awe3w
jk2VLJ5wA8O4MMMf0RGB+BQJLJ364O6qERveiLw8Rc46psZdesSeETm4aK1DBstJkos3NWGtYrtz
lqWPGMlv9+IAg3cGXyM5L3LqBbYb+ouRJHwoTXMDL1MY1chGyMx6/VamF+xldCNjdn0ww8nEY5TC
OuAUiBXx+weuCdl5q5KGRy7Uf8tiDaTpihiSpiu/QT+5TZNRYsnGibxP5T5shvnE8Yi2V0IdNMUa
NbO9DbaIon5Hi++XUCxWN4w+tOUG0GjOOyzeQvl1C+7+3G/x5OkP7mgzFqyTu1mTD6e2wKlsUZPL
F2R9exjetJOUlFaZxDCo1yyOmTvzmbTvmSpPlIr7gwL9o5RswqJI+deC5RjsRVV5/c82tj9C4WX+
skQQ5j9NOj6a+h7koMcNkbYO/2oMpyDi6ncUlNZaTJpytsTTd4XQcB2QeigNzHOSRN4m4tOp6wqD
KFgbfo2YU21g7Bf82Bu4BZAUmYqRYybyZhCAlYBepFKvTysuMN7DYyJkO4HWoNq51I+rnuhO6XXk
IajlK4/M81CKEkcrFrgCxO1RcXAOUCLqixkC3pBNGLdNyxmad7B/QFfRIw3nN0uvwNkO83k3hZy7
Cxuk2UBghyTjmk8Js1S7mOPOvqRl49YaXO2uo6++2dhe2MMlT4PAgWT9c0sXkn106ztKsQ1Re4NM
sWV5iNGELtp7sRjWOWvBhUX2+/eUjA+Y6ipfh0osZzCPuTuNAhHAScL+dRej5/rg69dZO75LMyEy
rY97MNpP9FQtqZo2b5l3oZBv0UWv/ZyBxoJ0CNNhmpr3V8+LB1JpsivudyJqczOfLb86jCjdDT5V
IfQgEThKL2KvgNzhJK6b9jhMTcPJGCyR0wsIKm9o3bvFo1NRGF84XLNbN8olZRggZmYS/Ib4pver
raekf1nv2JXpwJ7f1KSa8jFpXO4JmficbxrLjUtNxw1DkaEGknFhxx7HRApOnJxWcB1t5eEOniHU
Vl+t9bcLgvep2RXmc9oBGOb9aiXEGBCY6vDzz2Zd/eH0YaHwP6UqQKPcm/3TlKfyUWxDVzeKOfd4
UW0RqYy98GvGqDFqcjCRvJ4n5qsYMzELhy12mKQ7+Yid0ae+2W0PJ/aJ+GTywB+NiXDxEGukj+jm
tQL1ZVn1gfea07YtcquCIdnhuehk/R9hp4VesjokwK1z/exRwmwcUrOsezmh+ql8XYH6NLuDq0uR
i7kGn0JkvIGz05yldefKnuJIvZ47fEzzADRiDN6/IqBB7dJeMApLPKT2hlTFjtUHiY5/jE15Q86j
0CgEAIZAHyZrdNhsG+EOMbZdm/eBvDduMuPZBdjQNQuVu/8b4bcniQaMCJ7sWNgaQI+LTJ+ILhrI
MrYDtZCM17okIQbfr5UW8ZqxunvuI1aq582BkwxHjwab+UH1sIawErSXzgDfrop1EKT6U0nPG2sy
EsOxScHZhhguFPpkkepVWKnoqR0GKRvRPB42/hqR6x2Kot4H/SaaTdAazK0mPqt4FJxQSXZeaisY
ysmDQIA3Z9HyIyAMvTkEVagj2VAztp7NmRf0LmP4V8spJLA5Sg3oUtKvMJBbHaTtiDdR7GWOiQwP
86q9nfqSQfLQbpLtMvsM8tZ6FJME5BFRjw9raVVRCQ/zzEVmFfjQu0AyxvpizafDS0A3BHD0trkt
UrrS08rr5BLom5A/eLcIEm7G/5E+mBUyoUECTV7lvs6J6XfGwKpuYo4VNRensxvYpY2Uf8FTic+I
bNT6PIYlNTtgarf0lx3CyxibkotC+G9trb3n1P5RFvP8MT9W+Gif9fto0ugRZXRBsnw+7hjHuyPY
i+yP65zUbfDSP4YJ8r2KExA9zfSEe16V4C0unH0Yp5coDxwuqv1MKxkvaFZXwA9JSCH7odLDWufb
BJJpUlTfh0lDVdphXICBZm9VHWfPSJWIKndO8aNmsWHxbb8SjFM+bp3ew3PYeTk/OzuG+PGTRn7H
CPwYANn9/R6UUUfPj6LD/g9gzjb509E8nnV7SW1SjJxsyD3QeQN6hqXpwV3JLIG6t7xv5n6Cd7jo
gMztLmmszuCLpTVYzKHUvt7lRc2RAMw4eMOl9Lrcy/dmpgyVQW7ig6BFIDPguvGd92YS2cX6Y3fb
mNXry4lddikNfgjbh3EckUjZ9MEDefXYvjHmzMl45c2GDwOB0lfTXuynCqknFk8ylMtNCFuFytMu
KKJXSnodE3p9WELQt9GPXFvpmrQjw8rqKArOCG9dlH03NJqXwTaoKXUVN645GXLe7hoNhG5rACq3
iOccRFE05CzyxyQi9WnkQDYWQfH2TZRyq8zdFWsowuO6lIgsJsWTuV5HJP7/GyaFrcP4E445yOkT
O4n3y4TdHdesXdMSZMpuKOJFIT4gic38JzCZ0H6gyyOMG8KOtf4Ur6tiG5ogk+bTlDXZzXe9g7a9
q4qVH9W4S6AI66ajJjQzCLMmL+q7CieIOBBOz8MwQ6LFBAI3sxzXg0So2ZvekuH0dYuvLBxbpFHa
K0WMnXE74mxle6L4vBQnYBOt5b0KWWb7/sR3C0Dwcjs6SXgYTgA90R0IhFRjaQFn9hbtwULsCOZv
DnRBDm1RoBXeoybTN1crc1QJ0Jv036si+36wagLWmqxwVtT8a0GtxDjX7dZT9n3KE0eA44aNDJXF
FBQYrqQ9HQSwLIbYcdZFTxaS/29elYfvpBTscKwLzCbALaiOA753YsdPJy90FvjDsBkuDeiytNAE
aTXVUwV6d0PKHBPanapjz4vgrC49an2FCaMv7zzTxFB3FXjInobZXp6qYl1yoe0PUic6onUv3tTc
TLAYxNew+05jpSQ4PdXdQ+nxfwSPVnHsJwY/q9NknjDDO0kbtKZKRJg0qLCKtM1Ebq5VI7d8xpi/
bs+CUh2dmBGeq0RWHB8IU+p5ky63Fg50Mv/IzrNm/5vmggvUf5HqPc3ri+tr22v9l8fVUncoKppe
/fTFnwXkwxNaI4TbUzhF/H6EGBou6GL/U4xCBxvN2b4c3Pet5gTpqvhhN6stSkF1lOv4mFLI8/6k
3uFmolHg6ODNQqqcq2bF4Tj/iUJbVo9GtXTGEOPz5ImYzLFa/n1lxLJ99fZwoeax7qu73UNZC2Su
YT4LNe9dcp+xrBc/EagjdGg/OmHXmOi4IXOivLJjBhyxBCuKq+1M0v0wn622dtKlta13oPt55KQ3
B8qnbLQTubHcGisDyazIrQ6i+u/o6/GuOWoRsLhua8Qd17V9AKkB85rzdzoFzYkhob2LLkJYufl0
0772lTsRF29o2KnY9Mt4fuG6NdOGBgqAwO1BIqm9gTp4fJAGItSBsjnTVvEcBxf6sXLw5NxasDac
6J2cDclW64qS3evbqY+7wuRP7h9sFsTZcTyUy0bNurPeUFT8kUAu5OYzA1jpuEX7NAL6/f8TbvZX
1cQI9MuOq5ce1JDMClv1eW1ZG2wTs9GvYRZkW96D/e9xLObyo/SK6bBHDtnRNNabxRdynDDfyOwo
ceM6jVDw2jwMOjFVwoIROLUXn4WEtge6bs0zGx1WObmEJ23NvyzNSeJW/oVcAfv23gNwlJg0NH3/
9SStTfR6MRPZRwEDe61a5FEHGCKyaaxaBVgnGQjwiea/yhNgb6t8MLWDR1vDRs0WbCCXFWMxkE0J
OnT9m9LFj8ld4vGZuT8q/DAhXdNsG2SRDcypkIeMDKWLnu5AqVqr0jbTcQ+G+NznJZOsIMuQUKGw
/O6sVYd8ViOBSLs7ATLH9Slq9FXPInzG587uIWg9XdR6rDN5i3GQhOa7dB0hJaZdhb8Qkxfj6rhe
srkErEwva6Tdq/zNvDEXimUBPrJg0maLMSSYW2SleXKaiRKWAI8GL3VU/5Hth+iISwEUqjmGQ5IG
t9V7sdheH9D2go/1J32cZygRFFSzt35yX+mQ7jlS4U/LV6Aijc5VYG489sb+kMjpzun7DNITeWs/
rjqMZkErvQ4KNig57IUDMOwh0jGNtXSw4LR7MkbCQfXmEQWIiX+doGqyLp3ujIBD8lbc+TTkud3y
z71trVjMegi4h7D2ojaUHF/Dfo6YQIt5b9twPYCe9qvIoDq4GVXHGe2s7b4k2r52a+rd82Lv0tS3
RDKuMTO03nwH8en4Iqd02BdGLIer9zkLMF/3Clo1rVjb7L526PJwCx8EeBjqkR+T8YnphKFcaHwe
uE6yjgm5fKaW5ETTCgrlJiV4NBbDzZvOXGzuSZb7CwIkB5XMeYn/EB+XoUjf6CA/+AvVCfJ7TicU
Z7I7+MoO83JJCJCOTs0+hDuJuOx/7OMh7qpR310yN/yOnJ8Qly79QKGnWPrvMZ0gOWJHIUyAry6l
+WaSS/S3Eq+1FBE0Ld/Gx7rB5EdxABVQQ4wfMb8PnGRzHyZF9hsaUgT/KPTPC0kX70wcCcqAHsKi
XKwyyZzCuGvJFji/NxxE4Q7mkLyIWM2t1jMbRPcElzXDc5c6FX/POEbE5r7hpmk3rXGxrMJKEIUX
he1bqNR4P72xHVJl7EEcATL2+pSOJgMIWhzS2HfNLm72YQ7iWJx1Rz3TunbgX2bJQz/KhRElvKP1
W5+J7OSYAPuu9p7KHHUleepvbywOAlhdQfXXJ824e44VUK8VgU6LxsBN6kDuqKUHeFDIedTfEViI
yc+MZUJxY85nOASceMcUBrixfc1KWPBqDV2ObYCYI2LC33UOxw5sbmavabtadHMAbMaiNp9noBPr
sRY9hn3qEMucM+C0GGgeiINqkmdFyY800ad+OCeN6tNQHfwY5yAPDHn9zzHOHnjyY9neTE0+DWHB
DfaF5gMV1jzf4FWFtrUOVJAYtehdqI85GKVGE8eS0UOmN16+lEydi0oLvBedLkkb8vi0oUtoND2e
shPvqXXswpEcPccp/r65Qi/3oz6F7b0q+QfMkMtbsl3V3lFximi5SN4HGqPr+LtH+1LJZYZ0dcQZ
Xh2anLyEwCn46doxhBFmhTW8LzBLILjuF8hGIz4HX+d2a3IUy8blblnzlUz6JUuau3pAYttXnvL9
dOMZaYSlxsj1ShtzstY6SHsYTKpcAKFkbG1R08pr3k+xQvhXIV623kEdFwhXVxdZKRAdR+kmFfqo
grzimy7G+ZYAtRf53FExxRIjObuIZmpjvk7/eZq/m5tP6z1VgWGYtBsrIQNimZv4EMBFn31pDvFq
2BHeayqi3lhrRK4eouOPPjlYqjnwgYca9coy0r88oYNm3ZYHjZFaxsf9bEeacJQWmHnfHiKFLhl0
4p3IBqPNuEzdGM/mUUyqhlSu4iubNugfW0QkB/uWPXkZjnyjiKBYf3F9y36Pd6uq1+DbGvFHhVq0
n5TL2HcL9ezohNvNYM645Bpcm8PCwH6AQmfxdUVkSpDY1lSWhIOboh3Yfag+YgzEN2bHcLpZEXjf
xA3AQdQwSgEouU7SS8GqTgUMsb43yTvu7ASU8YuSqFcC/cuZFhjMy2/nzxGccAk/pqVw1S58aEkK
tWi7L+32qJFwyILpiID7ahquVwLnuQLxUHP0suFieCgI+4dT5icxfI20k+w8ZTpujvgdJ2AkKmbx
5GANfE6lK+r8E63uy/QQkkmIQArcRXJkR2Kaub/4dHGurWDiadceOYytr/8llFCkYieSoyBS697L
n110VV/Un4mhsWpU06P1MePIA1/1Jf8uylIuVwAilPgfGeDStt+F9CU2Ffz6SrV9BiF91OPIRSIr
yQs6Xqm7JYGHCWAhYWLkcyyWevMhcsdqc0tt0HJ70agTKuuk39HM/DF8z8DNDZx0Y4hNKUMAR0fC
oE/HvJS1lt5HP8QeyzO0PA5yxRXaLSRRWHDGynZ8ZIwYMV1zUKQWjc4DBJ14OBPs7Edn2AXv1xB6
jPw+wy5jL0l/wozR6MvZbM0nGVPBVbVWHFWoHRFaSHCLpE72jKAmiMAv8sgYTEYRHjeMzc5dql99
+MrDaEdxmDBbU6F2ZJzhmT87k4ZIjMDMtQzvZPCYQ3MwdaxuGLMDWMNulv/Qt6NaO9loDVlGBxla
pszeKM0+tKRbkaeF85Avf4W/vL/TKRCiofEMC6FiyE/ShVTSb9qyz0w4s958XghpkDqYaALIBolN
78LDoZi/Az3ZZbH/yncWSH/H0AfpndHvt2PbPZNXl1HBhcb+epQ1cKAOA3tj3F9UHH35SgqUXxIj
1rbk9KfRG2DP5a1zE/x7pSqSoAOFs80G1hFYLgb26HpHhL415pFGfzdl8M7Ln6rF5Gw9mpA1gOGI
DaXcVj6uJbp5RnBESVPefD1NeUWouRuPypoZxKLL36ec6TUZZfSAmYKW7amxRNBxg7m6Oal3kgko
Is8U7G/Ur320IxrFbXPVe6pkhYE8XKsz+nIadwwtBqHPj5stJSMvYmDz0GjKaW3nVQCFzrRZKPqo
d2S3QlqN4pUHbzfItZO++x+XYcF77X2l/89ZCuLvkEWPXWUTHTy1bWqwuHNjAhqca9vGRbjIoPnH
Wa7vv11cz/GriuOO5CBHHfzBff35UMt3KPGjaZ15y6/85odkTNDtwJMlK017F68jTUC+nWN3EDDQ
LMiz0tpqwk99ZvAuDsjXxNAyLIzdSYeGbQyGhhUgUz5QqQgcoPLHrLuvpaW61gzOZYSaktmH5Kdb
bD9F9CGFHfqieGlsAHTMUrLY6pxNQ9CXj5hdI33FkXH9LFa1UxG9ePxmUpi7ka/HKLUan2yRXsO/
0PiZNz3xWfhseGkqb5AgYCF3weDah98hdqD2M5N61JERHiRxpSjaZ9xADdobOnJhJ2tYQbPLjbDe
1JKdHSmkgB2worbFxzgH6mV7GNwVJlfCf0t6KH4JIMKnsIERtOk7qF8jfPLsDkMVAEehxiYU//7f
AZq1ChrVt1ZEs1kYaJWZa+jJEsKhuKmBJcChqZeXYbkSVoKnXWZrWKp+BYao1ItjqksHcxqp9fM7
b7knWC6qah5ffOkHqoVY3bJE/Co58l8uaF7zcppzKNgdCMIj1lZ+cHc4Z+FcQJ8ytaqwmQdJYAgd
I23M9J1A9d5W7VtI9okd+BELP2u9N3V99mltjmuEqWDhIx9uxHY+wEQGZrY9vt4ync30tILcYUOq
JKwbleodl1+dgZzaoeWZ2QBQrqL0FQSccRtqSY2wo7/j5AxOkBxjUy3X/nMHZRp0QVn9p3pP4IxJ
vOF9ckl/xuK6jk1oQaqXvRpoez4vkLyi9TXjD5PL//GGAyNdpIb5nPAcIH5pPj5I4T+ons2HjU0/
ISnzwG4kZ8DsKiU1DSFjTzQk07ZC1J4xf3cgprknO0OfmfoqPYVLGdHWBzce9fl2vMy+JR8+vscb
y1yYuzVQPFovZ6duMWEM7QfXd1d+606mwML8X67wR8A6hKxse3D4yPizVwftNFUYISzK9lsdeOFR
fZzDwCEHtatMRR7hEgl0SFE+asMgT6iqSlWZUqJoEFyMfqbDqilaBL1ZXC67CPgq6lgtQhGO3RlJ
ER/OL18BJn+2w3J5xEVojmbDQyANG9DtqzTLSt9PVSMsx9EuJgGVDd55IYOcteffxhAyyvh5AA1w
P01Ez0D3DWnljFxH6l4csr8ifMR9r3CCqtOZBE5YaCxg7OgpI9wSoOI5jQwS8HigZUpxVw+XHkYn
X2jSrSBCBW4+6LI0sn0IEe1jOlFc1Lv/5mnD9nBWJSbyKHWnSR/gRoGxKr7Hi/FlILxJBvnOG+fP
RO49riP1Tohde7BG89yP+sfXbMl5GSeyTMkXUTlARmVxn0Jbte9oZcaF1P/BRrwvqNl9vbs8jien
iJyNWRJ/MxnIViCaNcll2j3zsiXczocmOg9Wgt2PDZGkowAocENQ1wp2kQPS/eGB2qvvjOO7nkbi
wcC6ODk3Jp1/vQgc9btcwDB9+RiVBGnNOrMhy81mz92A2w5vF2j+Gk6jhmBZLm4ZhslmZKTDByJQ
akN4FsWfxjz6NQFf92d5o5eoIeR7FPM4GXnO0BwNXl7yk8m1x1YrT1LxoHff7aOT2gANg19AUx3o
GzRLM+TBWkT5+TQZ1xmaUbbMnevZ0bBjsXlnKAmiNG78S2YrmOI9vAWAKlzMTwbfDGw605oFEvCX
fLQ3fREuiNiV9IAcrni+08/puhcrvHK5BeGxiAJ4ZQX54iBF0ONslvZN8Z8Ek9nIvJp/yR7k9Ys5
GxTjW3JvmACoQOvoAkLRIO02XLIV1kV8NXaBNMizVkRYPfDGiFAPzh+GH2YHuUC1VeuVWbIXyJwG
U1kJiedytj9DLZMVIdbYeiIEuVHmTGveJQyXF2zKU371rCjJ5eWqhgB5iTTDnE7fh/kyotMGRRHd
YCJfSYn53MIWdvhif0/pDYlgcKiEW9fOQNfdXeoakyjkZogRowtqTVGJGjx+RU73mqo2FDe3YUcM
a2KxVsZ8vvNeHXiSr9Kpo3DYf80KlheC5Zno16ewBieG3MGOGIbojJ16dVbc86FGcP7Es8vxpkq+
UH27hzxOl8HtLx6NgTNXrFaU4G6IgvXJp5QIVAi4fFy/+/WBJNTvUtHgdCe9886GD7ReSJMJkd8L
zPPdG85ARJQw3LHca6QxfFmoS1SeHrenLnLyyfMjb22ck0i3Qq50XUsUHq8BEFl2/8EWEQLUaqMu
6I2pOY5rEj6aW8eKMd4RBsll5e7BMnk9DS7GOUU2Bvbg9vqhSfXqlUx1kmxN/ZeR9EQYcpRaqlry
clEWzfHBMu01U6NcMTFqRHhAEww4uMITV6ByeKDDrE/GrMDF5FzF8+AE5mHWz7a9wLGYv4o5s9Og
nuN3VDAroLxlWFmGsIlZxoPOAt+LNM3M+G1vGUHU0yVtxExVIVwdaBMq4K/Mf4tCarWYjFeoGwjc
Kfd/nSjq7JV+f92MoFo5j2C8WC5XAbLm/eP9q3ZPKI5vnA0rqbVHW/iWS47B1td4dxC6Ygyl4BmD
TSLyUM9z69LBr+i1QKT8JcgDnyYeNmtydAHAmaxGDPdzj6UzIuPXbiw/UawyJ/avlezXne4/TTUz
+e6OJjHLt3lyYYsm7UmrIp4mN9B4vEVaqwaJPf3ZM36bZd52p7Ki7paFEKJS24jPpPbIybze8WxG
1hZk4ZOXq/k3oZsyGonsPhCuE0gw923bWiEh3Wa0ekXN4mGzMr5vd5UPZl5XtQ4g5TK7pYT5QsvX
k47bZ96NlJC2pjTy+cTdbzHoRg0i7NyHD7HOErnhNLbT13ZscDTtbZ2hsYnu55zceSX850gcPyCp
fGxUEYuIXZVCaWDJsIoYc7e+dt6f1zQd55+cJwEBSETj8YfLVsHTd6fQf+rmJidYwMab172I6o5o
FqMkYWEvQvuOBDtz/RRmIG7w/gYBLYjXEbbn01YuaYZEuoNy01bzLQO+aJznuynegV3fuxMtIaXZ
yLZ+17/CyGb9toF6Yf6BGZIAlaE07mMK5w3qWN8nWoPXcbqluIoTo/H5n3Av+/MllbqJckZMFujx
QzNhoJsOPd2xauPcmJCRvKu9515uKy8Py6/26dS52xqVes7Q8GE1MINDdZNtYjJcHrY5unlo84cr
MdKC14EXZLgb22/0xAEkKNJitGmPJw6d37NMfNSgkSBiRuJFDeTmHdR+i2tL72r+doxShVmvgbGh
kYXgaQXOY7qMpFKKe2xCYUE2RnjygFn6ZAuG76qjKccqH9m3yxplhLUeK6TUE33D3GnwuWakK+zq
/uyzdO9pJ36uvdIz3CJ8a9lSjem4EAsCfXPTIkw8hUlR93HTOTMWykyoxiQKDvs6xE2ZBck2u3dn
0Tvdef58Vc5xXjI82fx6SgjTJWeBymw2BetT8oZpUVklPT7kqe2v7BZ7eU5PmwA+q7WxCmypzxS+
e6gmVJzjjvs/i0s/VEpJuJIlIR3yj/PW6jBhCRwuJcyUWycTPcbRm+xqU0SXBI4lN4ozJDmP775S
6O7lg+G9Owx/X/ldv39mJsAaR+5WMGXalC+CJckByTFDN2aFXdNyGhpF+xWWLfFpG5a99zc2z3gi
YfbKHrwaUCfPSNbWGBQ/M5laQhvsbnEkbgqOTEeJldYuY+Zccboy36Wuj9egKfHlX2NCQUh1x29L
9tq8sR+Odebzs9XwT0f3x3jKLpvWhh2/OPRViKqZuHRkgLpDKLXgPpAqMEQ46zTD2++UH6aYaAuG
SAgbqaemhejbpb26Gp489ibhBgaWBmZ2SOds4wd5i13ag3msGcUumoWv7OOauzcl1wOhqYD/l17C
vwqpoYiF1/f7Q3s596WHitO4SxmKlfacauorWdXb8uDzghOAiuw0Jh1ZjyG4EblLhy/sewX5ORdI
8y5qPUmpwISPEMEuOgAYirZh2FVqSidJTsQ9KxV88qXtJB/t+IHEnf+HkL0Z8n7PBIHJuMHg5k1X
0m+zdUj+PZAo+xQkuzhz1zVDaExKEbcK+IjwRCwtbg5qseITPzU//nyHJdpq6sIOvkJ6Obecp7CN
+nNA//ihltntemSpkmaMzzxw+pjb+RzW7WmiyrIOgyS6AVxLLgLPJj+aWu23R608Iventx06LIgy
XMdWO7axAHKxqHJNlRyDn2fuMU3X1YToH8K8kQMXkJ3FNbc1iWntblmru4O2oWTqrjJhOthlT6gN
K+dlXg5Wxnrc7tK8oROPKANR4CtSWXUnvffhURghpBcGI0SYznsXihdrbXrIYZxrcfXTJIVk4Z2M
IsrWKaau1cE3rcVDD4q2mjhlIjFmSEiFIALnzCaNk0lzKLvd/FMqsSdWjnoTWpnJa3cGhBtRadiS
5wnjn2P7TZ82sDiZgXsAeM6/O//DqUKyDP6VjJdc7Z6VcVoB5rc2D/2VFB4ia5+XdxIWjAiPd+gr
HOyBI2+MOMsDRuge7o38rOQ2f5T/9AEv1oiKvhc8myxzf8tRZLSIcOMzpk1ZOS3Mc0OjlbUjxJVV
0PHRSSU/52FpSdTmzNZaFJWuHmpNYcFzPIWY936eupcEU3yqdOlqPQtPx0UZPLu1LD6MjT9/9VJx
lK1l8WZiziMs3owP9hMc6WjdGFWfB/PBL65jUreKVjOkugowI9ULz8JXfHx38u8eVlPjFyJwniDs
tqtCE4PgtKbd2WuoFtGhX6Uibs3/d9wGTYCx4ZHAz4rhirAqSLyAVmqHl8XfFSOmY+4N2H/+bgwS
4CbzshgU3bNeJvcyWzCpV/CgpZJUG4aRoj5eM7x0pP4BNXBfL2GACItk3buTprUhoDeJwRNtdTEX
b08DfqFQlHO/aVbjATJ+FNz81XWgCYuGSh/U7Cd9ywpvD/SQTwswqexVe7hfq/WWYWSXDF/X70/x
h64ld57LfhdHAaJpJ8WkU+SuS8idJdG5AhLW3IdPYMRmxAsdidLMTJKRmK3Vq3NJwH8eVdrl7eNA
oAXu2Sar5xJ4LJiFlnZ7cAryzeKezV8A8N0yWuDNfJkU8Guxi8sAe+74lygC0a4RnAPJDFQxpp+B
fPeLmU69RFxEQMGSy/r3Uvb2J2FlUEo/DP775siZ/RWtXpjBP5VoAOVHE4/dyLlI5b/KtuzKGWhd
0I+Cs9uvOn1rkpGj9JEltLAlv5iNNdXI+bCk6bI2DKk1tFxTDEkMlwDsdXHKLBB7iadTrxtx34hn
O5Za5Pxej5b8A2gQl1pv9Hf/AB0MZKE5t4Em2PVPSTvtOZmO9sFnJMIQnVyAEwrTLphXqcysZrbA
tlEKqNyfqYCVpZnjJ6eQGNOtD8ccmpx2ucStqhFb57xM6gS0Uv02DpUOeWQthkC3oulEY+NKEykk
hn5l1hNOwLhs/rTpYfgBp8HGKBGM3qtGbcCYohyaY58gul5Sik/QbHkpAkkhAkUh8Is1w/F4ny6k
qCgV3fIYuULIQcf0mrSafPoP0pMEBsYM9PN/O4RqPpXYhHSJ094isH18ZlQEHeG6dfEsSuQmcKJy
3pYPiftDFULB83GZ7/N97hEky6fvuKBsAj67bj0cXxQuOZtHAKKNoXd2lE2MxhC7T1PjYsP8ZpUR
8m5LDcaKJM793lw1zN/jyyanRAxywzgC/FbxIeCcD7B8vug4xLvUETfdZsEmzhMtlpNKAY5aZKHt
Wj4iI9lqtruVJ7nUNAZesEG2VTxR/Id9aXZfZp3YUlGxq/LvqoWvg/18OQa/xEuiOQ5HLX3qUf86
j8BoUM10C+anEFi8dyco16EVIlfxfHfMnAasfrxoQjOs0YbqzOdLgPfEVXpErWRjzO9h/Xcl2ZDz
fwxHsGV3aOfYAs8Uxn/NjRIcuPbemeCvfi+uL/LbPPxjmD57OvWnblBm0hhoux7MAit9KoxO+oZz
PrdX7fd8nsIY/O50eU7w0JMEL6M/0iMzWU6fNQjI6gIA2C/dg6yLpO11ZNeviuJgvhgU5G4ic2dS
+Nv0BRkxsfE54XGuri6H2Y9SXLIepd3XLsdD+ttWlVHVc53feSQzJY8mpTGgGntBWkYQ9k52jeYa
T4wJ5k8IrlNwzFxUJ3kGUf4Q6nd3RJTqlULvAOnP7agcsyUT/vuYlnOao+SuovjL2gj0e928ORb2
FyJGhTWa70zb4m5uvVCzYi/1ikrHY0sjUld0k9z8fh7sCc1YUK/U2kPDKl5JwbW0xRXUXIPfwX/d
okWlUKF3YiF2GWibJWsFoVAR8u0Njlr7+bpuSpixfW+EIBb9jVNOfGwkgQNtE/nu4s04Oz351Xg8
QW7QqZAxDiY74Zl5eEBR6ILW/4A3apE48z5SZdpU1k5dd7aY+sG5qKBvHXAokNdjeaO5sjmFVJOH
TwiXuCh7X2LhTlJ/DHCQEfMjZFzk1+oVNwYgzLN8A1j6x/hklF8CzDCRagd4E/UJ/f9lGoJle9vT
HHkYRIZXP+AleN08ddp0yvhevXChi6WxBZFQafZRCC/ruSG6PD/EMZwtfzkEtDnEccrXadXUkZ2D
czSppOmk15JxXyTqpQAa0tbvl7fAqmnYsveaJVrTAZ45Arwj/mfbCnFnYI8gdKrAJq+ZqNGb4DhD
9x72E77P+cVEFvmu9XgQtww8HjGencAIokjgsUEzIGXEHn+Ntee5I45iT7M2vMgMsobUMDMwWOX3
uRhfaHShkbdhrPWwgHZ+OJE9FdMaSMomLAGoKzmInAFu92N0jaZIWZOBU1KtzWm4cQ/pwhmbFtxN
HLWjlCjwfvF3Iq+GzUn+F0XSlItORWN+qdkwDQCfTQxCMd4VDz4dF4gcpZNU7Z5Vucbl5hCXWMgk
6pUH2OUyHkisDdimRfhPnFGcnLHcNUYeWee3Mq0rKKQG6OLewy6HGAo5wPtAcZ5G4i+0bkodmVHr
awib2w/WG8zRIHNLLRv39P/jKQyxHi5mGCOf43SflawVD3j6XfhvubXgMVGDnRfu7otZ47IDbjgB
bdFXxMBPXviIc50iIbd2uAXk96b0XcPXh7nkSZyBE8azv2NiuypJjkZuHWBzLqg79DlQpuClOUX4
DoL7sNfORG2cGfSXtAJa+ZLrF+723vOo7RKbboRev2gTYgU6cxcxputpAItN+Qd2vyJuY/dCsRul
64qSlOQZNkOnwtloJ2a78oppB9q9NxxLmJC8za8xL8UgtCBBk642krfjMtxeWDl9j4eof+T0Rz+Q
Ww+TarfhA4iKR3TMlnPeq3E/rHEn5uIYRonNVUV5upBU9gnf5rNWF510WS25rcoQI4R15GFUGbyO
To0m4wwwZvqISuCxNuclP9W0zaHAp7xqkPdghZLSnEmwomt+UHqMdWUgWFC5rU4JKB2T9iC/tj47
A3s8EilXEk2yR4XehjYq8KsR3EgiEI7VdQ7/niLX8wSXZ7atD7YzXi8JnvAOxaRIlZ71riJKI5Sk
9ekwy2I+qQo8Oa4nBtj0flgdZ51LAb01Typ0VO7G+GPbfHL0k0AwaPXWmz9KERLemYXqajoTISyD
VWW5y3QQTldPu1x7fELlHaQrkLHfLCMJwML+zjrTmSuOkSDglSJXFTtAdE5sW45AyU5f1U4p94TW
uWItrxHuhVV7arz4sgoCo0BT6oJ416ZscqbrRFE4S9ZGX74f2ttDQQRBZhlxEnmh76EKAfzAd2Hp
HDJFORV6AQcxC/MwQ3tfg/SZWF8wYoB1ENjfzj9zkgL0Nxcvb/0IQmKUJYXRnkzXRu5UDLlWF/f8
G4/sRcuoSS69hMt9FQ/qPG3+oZc5IXX1l3MfdVD2bq+znmRpAFFNFNpSdVkihBP8cSM0hdBfjBN0
4g4dpv/VSGYk/WSzZYMTyrkP1XaUNkvadwpcwpVvrA1jshayLg3mi6wSOdGDHzsCFKh7KUahDmMU
+N5A/cwkk2xXVVNULtMRV7OEsukJTkndn39ZWVmFpvbh4al7m2+vcpfloyWBHLadsh1hS6iAF0Ag
LY74QxAwQnroWxtRhO19iisfQm/nG7yxlKlnVSacJlX2Oi642KUESK+kjiBy8Jefw9OwuEFcR4mc
UGIpIIJgKpwsF9fSZNQYmAC1jldUfz9N4lMgXgoCItxlpMCsSCbS3jBWuqtHRoFgEy79IG9SI6cP
qK7sFSUvfVq+jxgKyWwvCOpsD3OEqdWc8EMno4jaWlSSNPOwXQVvEULRKHqaXMm17OINJcojC/ai
tQ7zhVR+PxXeNt/i8q7r0KmWpQRmw6G0iVXIZguUQnv6N7NZB7JZ5Z2dL91m9xYbf+bJ0HE8yGdy
ubULhjaXhbbPe/i9kIWWBH0rlk63/gJnKmh5pRCfmd5qGhBls/mch0XBmdYZCoz8USyluA6K0Qpb
GnKKhTckZfz46asHYpRiZavjKC1aNj7CtqOs/4nn953aVNbkijes1xtmPwdjoEs926zWeQy6NOP+
jRrDjVQ4y2XoOZeZw7Z8CjmRSmbEI579G7BtgIO9U6yTOOQH1rwGjYyzUK45ZMpLx984/i4Pxm5F
Px3ETsNfyyJkwp4piEzn2gcpQNzFx30YgHEKqjFIcIV1twoY3J07KcoprBywH9Inc79XjoZEhERZ
uKQhN5bCQjA3O8F9Qpy8XiSpoo/LWHrOJrnyXX+ehSRzmES37a/2NKGBUFzhD2Ii+/WDwBZrojw0
RKSs17GfjmbTf5UpVIwggZz9oXP4pa9l1WsRhDZG1wHUxxr8a9cbXtXs7RfGFcB8F7RCq83jWytw
fE2mafvEcTpinuXQQE+OQfba2Ys/l+iVdmNfxCgFoRAJAOYyUcG/ZyOrzEJFasr9cR29tkEBmsZC
8cru15bscNw3aaVXBenT01xXL2XLge7YpcceGmZ58NhmrrHfV3NFqCRlVGh8BCvE0H19+QtTIlXx
fKaHCScDglVkO76fipURaBECN6VrSzwhJ7tx+/TkYudU67M3t6rukiN27u606WWEEz3wCfuZg/jr
/jcw7OxPR/47+IbgKP9Y6lModCMlND6TiUF5EE1p2pHE7Oi2nnh0TqmDp98uSyRlMZyGos+Y4Dz9
lPJqnEkiyN/8iLl1mW494v4A3afHbwa/m+CvY1u692HToqu5y/Z28cH01lSESpJLIsQ7Tqyp5iDG
YRh2RMalpmJcJs5aZToFnS0WG+TkZOotSbpkinTI5TjYr2OTP+gthqfoxfTxmOg25kKOc0izo0b2
70M2HV62/K8J8YcBJrTaGUmVWdBU/kSYSq0rFd4/z5y2PoVkL6ug2xT7/Sw+J69QgexTIz3U9upQ
hj8WNafVfOv93fyI2cX97VHe99Bsq3WCHAkItVd+BMxtV18ESR1jjckgRGdjuYR2wb0/ENtw2MGM
NqiVWsKeDyrr/SOXnDmG7674Yr+u4lNbqWkcFMyIMFzRwdxizp7//K8V836ZEYyG5Iy3NJUwVLG9
+fKMslVwhV2XpCqRtNu6AU8pgkm4YI5HQZ1GiwA3tkCW7vNCJTEUJ+eYocOtZYVBj6pC3/Ji8HbT
EC7PikX8xezx/ei9BEnJH4YT9g30PS0tmIIKbx9bauQdoa5Yq5dGHeLBT7uRdltovtkX/OpYELuH
7sdrxYlsAMuUSGjd7+Cq1d4NT0dz5OQiV3GGBYOhYBKgaTRT7f/ewspxC4mZK9KxDd0XJh2yIrVg
YOECou4BhK36TfWGVa3vvzdGAPd9dmktu1+HiVeP+tUjDo8w403arYYylQoUfgZbXEkRn685wj1c
tEOLtuOdZPq9AyRDRoSZTpRfeRCAUyDR9J/+b2qnETyY9Qaw76qIIcmr3DMaVFtiW/mbBTxpFhmn
TDuyIB49nvQRtp+hWQO4CZ2RsTubIxant6dAW3SgdzsM0LsP+CPHDAazKY5+f9ivcc9p+fUA4QOm
hxlvYR9LhtAtcvNmizQEYjW/ZANNNlCrkwKbjyihs47xkoFQ0Cprp1N26De0tgaSH8fhNtJX1OJF
5ccWKqt+QbxAGehzvcqeeXj7oH1qv/85TW6hDPn2dRDcbVq84BO/WbO16D4hJlT9ldFIFcT0xagu
TZXfn0l16ybSgbYdg5upQ8ZmNBhMbhrBjFYjdE9axlyCDifZf8fqJgwoSi3oDV3mmHyHY1JhhPEw
P4zUrR1SWvZwS1uC6B1/X9TPHcsNStdQw3J1gdOT/YnEKv4jpZ8sMEd93DnAMqsKNz3uKtJ3/AmD
MMCUjm9THjy6U5n9UB+3fpHfOsfo5JD0lFFCAuxBHTnsS688tiXvD7k8iUwvUC7uSs57A8tERxG7
afRWemxkGMTWl1ebtpzpjPEWrK7aXmOzHQXH57nLr7ZBuJDGVI80OMEl62iNMdnpS5KQI8BJiDU3
k8FW5jFReCoxzG8xkUjBwuWnxr7/OVonccXIJ5L6nxVNNc9y2J2jVMQDCkZZ6Uaapc7Xt28lZ4Kf
LbGgQtoGkASY6oS7Ub/nUGnaQb/RgnrFqv/j03rE+vNx10uZttrNVrh+XF8gJXF8QQaBBIdeTvTz
gIK3KN692IUFN96cm6I0UnNr/AAniHxcDnFjLSkYLHhRl2dVZK8Jz+HFuoyiCJJcb/CBjAb2dc/C
sTZo2zU/OhRYAYHGcjN1kMS4EBgFnFd9iX1zQi4Rowwsl01ajBoVvu0EE58tEXlUWbI9QUHNvAuX
ASPf1JScm88bqJbQFYUoa35xeCnsq0KIAvnUssbC2FkQMJoQVtcLeRLs1KtPLJYxjhqXKWkFON+O
PZog5mOvX4CzEUV07c6YXLiodUICLUiHuEokKMX9kyBx5VzHD7TolfUN+GXg+nXRa2SbutjCzBga
0REBgmEAt6zQonjLKXavNI4xlLsm3aLhLd9lxGoriAt+ckMpPMWE8nDf5gnpVAdsxmguvXya6dbS
OdmJqLPP/YH8t7AuCZJfkv3drDKWA5O4clN6K7N68YfUtP16Ek2hh75BiFePKhS+DhqEDBJir5EV
UjXPgSAENfV23B9I21XEYDVEiTPTZ2iQg8IDZqSG0TTnF4k+pQSBveEHJYy7fAIyg0x6nEJCM9GL
DGtw/3mfev3kQHrwttGAMfF2lh57bytL8Ppr9SLzCP10256Ia/N7uuJ6ygG0BmDjIIK4wdZKR9Am
8WJNKHPYMv10hvYsoPc9VQN0WfBhqq+BjOsdkM8ULaoiTa4Xh+sLzaqvV5USkI/OLwVrH0KubNfR
75zRXNHLjlWrttGIRKFALbhTHm1k6vJlL7O4KdeawFawwhkl8dbo3TQTIzAzlbVWKerserg0DQtY
MuS4Zrx+YQkOyQVUSJdYmCQqn8mDjbVuWJcHIL39S46JgVTnsyNOCCA8NnyWsoSyt3V65pTmRnyq
TBpUR8CFm3ubzgAOQlrgNXRxxikKUSk277YwGKJ5RMFufcSlEDtFLFWWJvZ+c1aqV/ObGuUeH9Wu
CZWZ8N6/g6u06xuLeq9zl3oFWIgn9PVzp6LQPkEx3f+DSvQjY5IBKlAvc/kQegap25CdkhWjFz2m
6F9wWc0d0+w2ABdN3napzKRrwlydfxZi/yRUgLk4X53YT9ROgx8/eM5nYuJs87KLuwSl7Oj88pgO
N8ryCKViMTt2qjUkv4vUCE4xDYbNg6nu8INEvVtnOAkyOVaAvvVwFzL3PrjGBngazc+ukXpMtOsR
BHwQ1dXexpuo5bTO4EcQ4b+O/EGGoEGLDifaopnQK6xANUNDi+SfEBOxmvc3G4Zm9VGI0kV+rnX/
uTOgvGFyvWQ/2qsdUwAm9Ca5Abmye/Kx/gJwgEI2r4k35ZeEbJighJCvJPWp3hOk71QF3uEGUoon
oLD81p3avyy98A4kOSGWkvgWkKn1QdN60TA7qExqGaZSwRsHSt+VHTFNcM+FIzGSRiLKbNvBUJjA
7vIwAHl99Sk6ecMzw8KWodtzbVVCIP/RsE3a314aJMeKeeumI11J9E5AZcQzF93WT31ge5Xakbcw
bdjWoGSblWbWM7O86c6X1sdWxkhFVrO9g0DH4Z5VEdVzSj5YRBefe1pO+Wk66gupZvQv7e8q0kwT
QcAJDHs3HjtAlSYxXcN+HQvfgW0/fgNSHcgM0yKt0j5qz2v5aFkdyu+haiIUW3sgx3kX1QbX1Ypq
jaB3K5Q9RoPPN6yObjT14+E8vx1DraQ4+eFoJiiVuRPvoUF05LCCqeSwPCYiDEot2YiMJ5/YZGh/
OHxJLmhHRYVQ6o+5wwiwYENjmty3JkKruwiWnOQD3k9ytOhMuffjjdXQMnHHEenPdE1MOLCtms7T
CFSkXEbB8H9lTdRmrx9aw0bIyrL7BBlhY9dVdKw/4v0uiMiGGEIgU0lKZNGd58PQE4c+musAfd5R
m4Itq+T/Igh3z/AwVSDxwxVCCjYjpI9S+Vn6MCheqmXmrBI5IgUNSo5/sJ3LoDNEREFVRZ+HpqK6
Of9pLGqhPHFFhcwfIHN3Bi2JWijRERDbmxB8jnp/0hPjdL7pQ85iI+iWehRKZk5cJZU7rIQeTAQP
Q4ss6Q0mlPekf7Z/i+Ppn3yitLMk3lrEhwOyS001f+RgqFBM2RrszbB6iFGAzX8W4Vv1TcZoglvE
ogYKO0273Q2JDzVdORUN+SvuoO+0t9ITYXuhrgBEWTX2PjdM043I4FSLJ77qFlyAgmtbIu6KoAh9
4pV5PTWCAFT6d3uLF+m1Vc3yypJlrm5MNlMbpWElke/xtYO0ZgNalYuY9W164am6UssknSBL7OBa
6xR5AlQSLSkjBmZ2vrPDovpPGJ92GE0Fd+LTnOD1TlyjzKtZfglmUHNrbFoH2QsyfE+b9CryPWX4
2crpIe1UIVCNFf1Vq58ZDcQWwa6teYBCQ3VxrOaBDAS0qAgDBqhhEoQwNuye5MxrlA0+WSEm3KPv
ACCV/BZtk8BrX65jgk7XZkhAOU34snjt3ITISdLY/j38t4VWdcz9JKpXR/wwEkOEk4TY8POpX4wT
pzEfdzd/wRRmkJdM14k+QznPfYlK3IRG6t0Js425u6n7maibHkedFH+GU74IAD6LOKygaJ5dBgXH
KBnNEmMteAlc0drZcDEoCne0cEGZCtUKqYks5nnHBo+yAdm/FJd09gOdSNCCXg79vp+lNN7Nd+vO
zT5zIDfOeylrm5iQM2fcziW+PJsNMiE/+M/OfE3rO/QExQOXnyZjBrFIA3Dr+PEZ6kO1ypK9Nu+h
TTB3bgQvizwa45v3D0yGoFSefnv9a7aWSP871fZ0VZI9AK3c/yiqV0tJ/a9pIOMd2rt0yxWC8MyR
234DyNt1TzXt4nS7AMVH3MnZOyypWQBzB3oZisDlSEosHspPodtIw7c79mvdWcoJXB5JUTUrOKhl
v4oMozNYaAHmeAPxMvXk2Y5mYHTW9QjJYmItpjkwJN/theJ08VlcND+VsbbmZNvorjVf0qtLGmVQ
WcAZv5xDIsQ1iNz1mKV/s0euMY2ZOMdjVIKniUAGIxyyjDUip6RkwEItdi/D8P5U/+wTXiJASRXL
ZKA8oXPGx5H8YN3a7kkqNn75qRtf3T0EiVsQ0icZfjyUIiV0TFvG6Jx5mesVwa1Y9c5ozCoMzDOe
3K/54xtsByGJ0lFudMf+cci1NCzhuQfZ+eVx+WZeNspDPmKWVlmR3hPtej8Z71sqzDfk3sX1hrnm
RRyBNZjLO7qNJwUDPNMcn+PLSmCaxNVwgryoB81T4j2/dd8HIggRNMYT4eZ5ZG0tMB7h+stgsMng
bWdqfRjhu7OqnPMOQZ60wDtsfqV0M2IwBT+bQwdzGtFg2hFu7J7IfMTiXkJ7Fk7/khCbbJVhavVg
/bpo5JKnDc8zrDIaL+YP3SRHEMeHCmheFcezBNwKi5hjrbrhYkJB2MDxJrs6c0GQdUT9OoWTsoh9
plQQo/XDivPvyyIbDcyWzzX5EuJ9QqjsrmB5+Q9yFXyWW55nsGJkAx0ilTVuDrx3DSN8Zrze14s0
Wgd770qkZ2PhyV++8Q2PuXcPet0ACvoUjXl/P9kWgWfPYfICW7FC8lDZT74RSbBPaj8+CwWtOu1B
BD/8UYKmr0yVmt6iHrilRiT0dUMrHfvR2GlPWU5rFB6Jh8LcKjXW6XHTdW/NosuyYK1BqIVxsAmK
yEHaPoqGOetX/er3gAB6oL9AkRADXdegcRdAeEmkRlC0xWZbU3v6Geno+znId6pV0LFJAHDl9xWd
CPUQd9XFJvzt8vxkgSHLjJGLFaVO+xL4rUWQzhWdH9zJoa5MgPFQDVHa/lS490VzdEL13qVW0Zgc
leuHNoUDMkiGsJRm4kymGDsr3UIBwaJCBDMMyXgNs/eVWBTdEOlXH/Nu4mEPaXwCEyKuN21iHe1R
VeVw6AtfEyKuF2UNtZ/FaKtxyoTRTGiS0N/Q02WgJvbvAvtTjZMiekIDiHgjF1+3n7Z2faXuRnap
pK4KZieJc4B8Buxrz5KdivhxxKEb8ggiSEKlYdbwp0X9Lr8M0oP7fNDmWTVAFCWGBZ+effD1NUYc
Ma8dMiLU9pZ67DUqKIFDdhhjkfqtW0pE+axETcrWXS+AWurfzDbRwVTkzad/zvmKvZ02+G+LdZds
5OzbB+xRt2rN+3crWqwHWwU88TURgUSKqG27RyaGO0O4CSSHm+FJrkXZt1yKaROB7gwnGx552fl5
DEjA99rocmoH4x2/e/Tw33ndRHpUDek0al/yu3oRzXnHwn6CRWG6RDynVvvn+m8fnKHBudAPai0y
Q+GcrvkgGu6SpbAmCiPrVp6Duu3jlk8Ts0icne1rWVQgEXU+02Mu+8HTqckhQsPI0wRATLFphlu8
EwbZY6ryCdxfLQJ5iMWmY+WE1e4HPzmE69MW4vdg60sZXfnkW+BiVRMGF+UOd5iUwo2qRZQ1Nac3
vZ/Yi1nEf7fnTHs6B6ycQyn92FWbzB6OaASinFHATgkvzcsRjSmnI3EkMHTmuxkK5AsT3oES1hYB
7YMMjI2uwIXO9r5bzxyQkJ1Tga2wsmunKNNFJnEQqPaoL/oG+jv18yewTp7QMuIeCBPfEBBjiph3
e+XyuLJTmIrEI14bSDrwYj5XeFhNKLiI52pK7NxywXA6ljKepTIG6byzg140aO646ociFu0deYKU
QtHcuEjkEG9cdxxe1VXq7kQ/n++Ms4ZeqqJGp8Xfys+OVGDOrqyBZYPmmPM5jjCtQvH1aqLerAf/
Bek4x0lEd+7bWycPObYQ0VZ84x9/Y7y3F7rireIN7Qgd7er0FygvRr1/6EuUXnUOaXV5Xb+WHheK
Tu2uAmaB1cf+wNyLsBcRjIk+4W5Hl8pdtbRkWpGcaBASOxkFy4rU2q3iwxbuCnY+vH6vomxI8+OZ
1KSP9Z6rKzYPnuovEJL75d6BbDzDc3t191pyYFu7HN4Xn4IGlc7MlUQ+mJjLhmf7h1EqR6I3faa1
ojDBv2d10bsZYaI1r/bGRLtt8kYCdNA+uKx9EvAVpmKmXzVM3GReGU/3feqDJOBirbH71F4Ul9bf
b7JZpbUivMDqNso2fCyP54UPNh66auvwG0Kh1l44wBSeKWDZbenG07aZJ/2yjtzO4P+YblDsIjg3
07v2JlhuLDNwbgkVgtfEnG3XZYSupG65HOOzrEgeTXjWf2xslsfwLXPR/WnqUpIKPhvbFAHzi0Ww
p2AqFB82PsE9aXhObaJjmIb+VJirO3u81yB5RbvlzknFq1Y0ZDw+D7pjXaUXW5wXABWCkcBAsisc
XRj+tM9xD/pdVOJ/35s5JXHyEb4hODdcLyY/Fi/6WZLEAmaPaWtLfhsxfH/IIeyNX6NFMuCuD7ID
N/VVSHIDWBeVYA5NtkvMJpE0qSe/egVn2PHjRX+SOpI4hDXoTG7nFDRZ+2cx05KWP1VJSRJnNVoR
NvRLaDRMhpk1eyW9R6Y7W18RoOy0GHow7xpj31WDlccP/1tnQcEP3q8Mv/NTXxC7Z3OlgBbBziTT
7UJeOz2iBsoCulxZr4x6ccDFpBkHukz38exDajOgabi2E+QAax/QagJpJ14vF/QyWMZQoSynIl7C
aymYEVwoL0GzdcFhR8SZlgvQAnExoYvOzgeEJE8xg+KJgZv0YQ22SBUeGUw6NBzHstm7q896l+kd
YkOJeyERY9v9iIKLJBzuxbNrqmynq2lgwdxhX+4rofDOulr+FtY7K2j/JaHYK9kLjaVNfckwJnle
WQQdyMh8YSGpYIJsed04z7JMayLKHd/RmBVLtLy9fTCHwh/1sPnb+CaR44Z+ACqNy0LlGR4KoXVB
o7UD3ULC6UEziCiGHpOClEqHZ/XZ6748mDy7b1p7Ec9Ut1G+IAbT8F55nTAiLgwcjTCFtkjhvpLr
iaAU0Wz2NFaDJrILPd0j77pymJQr3dOH+h/U+RNh0MkF0GJlnRCz6YjNKmyEQV2mEPabpnrI0B+j
ep1fGoHhoCA/DhHdi7EOYlAGPc0z/v5izEcMBALyv10hpHr1IhbDVFUNiafLzbMIZdruIEZ4xur8
1Edz3aJMMrerYFYwLwDJ+8UaR6+ozx2I/jsLJnIQ3LcamD52xyupVJAmhia8IkaYamnDjQ0uoI40
l2mz55PUydM7gDMAxoUk+0k8hRrKNI5rzrIwrwyPgSUsMxgx9IFb2/ReEKmdtUkf6EorftQRtSXM
cSs6Qh4A1wVWJTrjzRTCN3K0Pgu3M8RmeTUMjk4h2IAEpb1NRJKr9upfTRy/B0mYblyLobCtkJAN
ycr5LUx5fVoraFgj5QHPYpwtlGQYuZ515E/mt0ONV6H63tDa1qXdS2879Fd3UZdmltqiumK+QknR
17GsFcP8z0lgmQrX0bYXR5unIhMGfO0gvhtP/lwf49mpQJ65qD0RD2LGG51L2iIzQ7mvUJuqeCGz
nNQspv3p+ix5X6rxoN10OXZOuvQldcMaH6TzgNSFh+sNRzClFRExQXIKn4O956DAMBj4WuwvXvvb
VvdONuVd/MNNNMr2AmWMB2otIiZvbgVe5XTjNFLLHac8KAv/m8yUKS568DAuw0UES/j1Cqdanc/a
+LlPzu8odtKoGZc6nXpvRIhjaGgx4I+ffKzaEQuxxd5sJQO/yg71VrrfmiUKHn9LdeLyh+x6ltwJ
ivT4scWwMe/zD3CXKZlsF5g1G8a33KXywursA+l+mUGjYseQFeVQVeIXfxYDi2GgWoJCB0c7lMDG
A9KYW35+R8uR+h59+BgBYsW1kAZM9wt+hLb61rmFMl4gd6P9DX0oKwjjU10R7gnGzwsKDPBQlcO3
86puW2r5sxO8H3e7aJH2qmCcHGhyFnMw05HdnKzd0YkB6sQqaHO2h5lS4iO/3PRlpUGsG+ln3fm9
4Mra6qM/OA4F4q0wPz4AAi+LAeHL0/kupttiFkiXjkmMnKGdLYwN7t69PwJfYFWvBv0Hl0VQaCmN
+Ye6emgMm28oaFZ6rp7H5AxyT5PSKAd0jmHfh5fclLYlvRwWP21wyHCsW6acnbHWTfTa8XR/JQjT
tpbHghvqSVflHvzYG91kknx7KqdTkBj8Vs3LunSp5GCrHJVcvfO5WLavAedZ3UbvVofhcrnzW4oQ
XPfyUTh9xAqRCjwqxz+4I0jR6TCyWl0KpLQ4jN1hulK4P0oQjwSpG0Nbxxsx0KC1wD6AMFmTYHwG
fpOHG3WCCWabRpe+WhiITKo35ibuIPYRwjqcKekp3iEL9SqLmbZ9Q85dgImVQw72FvzKbjra4s5u
BuvwHpUxPreLRTnxI3Dt+jSRUDWp3LX7vu1ZHLhWsAczdshyJMux9Wo6I9IIiH/j9DlICSSABVvk
X0H5kV/N07SV1kMy3U5ehC78P91JrfJa5xEtw/2Vzx6yEVUyppcfDU9Ao+u+IC80yXKltKvxI+UM
GRrk2q7+PurznCE/+zCK5y2bIGckWwczaSCxKJ7nwr7W6VXp/OB0BKiD6uejFYP0orhceA2J6XA3
4jWxuVOWOdMy3xSnTuzkiB9m1BezPzVjC/h8M8tVm7KB2LxkMlFiVDlsqt+SBgoWt3m1eGXipN3O
aVGaae5VNN9L7Go4rwvkMvqRXD63bRkHwAKw1irYkoWJdI9pwJMYOML4PQgCez0kmVRbMz3Gw0EZ
B2A/kqfTCZ3kFvmon1Z/fwrwp6jakPD1JoUH0SnNE2KuKhAie1N7Hjq5P6kPhrmbrjVM0xorsM4d
E88L/tuv1XSUEgrp8Ftocp3nvjZH2xElhC5mpZHHBTvRX4DRz5U71uQunskJd8Poaa7DTdUevxlw
h+5O3/PO0Ow0ZKyHGwmOAV1Q1NWh3Qb1spT4Y8inqAVjYkUPa80YIV2vDC4voWPsAgxxGPUFHMGg
9zmpgVH4YoaUQ0j5tOXlculQuYpxIO2JK2hKw7aSFLAXIcXFPUo6EcJPf7JbysL0oxbQ///O1v2b
2lkVrKJRQP1xN3tUDIq4/+ngjjOsh/uDGQcCrsmdxEsELmyCBGCBgHznOzI3YOe3ECmcMORZWZgn
qC7uEJy+8CYtgSSy8V93WFaqKQS4bmRhfc9Xx+x6ayn6ilYqhUZxx+choN1gGvkg4HiWVMk1gsnz
rL0pkof1bQwWA45YKH+mJ+TnzR4VLqT5sOVwT3AYor7zjTwv3Wwft9TrAQX6lPBTCiTYZ083GEV/
gUQhbUoGVJxouS20vfYPNzWk71VXfFYGKTbdk5MBAhzbGMVTP7n2IyHFhrwiKtxr7v/jWjuD+0+u
nYWjI0qKF/rroM8HQCDP5/GqfTeixAJOxXFTNjrK7mtxGnCpIa1lkP69h5TCWKDFToTstRH9ABMo
0Jbbe+u4ibcjljmY2rbmTsbtBEjpj1Z8Gq7YFiAGaoWN+Ifl5tn+7EXN38oGY+EG2cmnQJ4qAwoU
UJ3dlNB0IfHUOaAlQXjcNB+p7oI1q8a923Vqlo6DAAx46YU6UGQXvD/rrliNRK2Ps58oNvifW2LE
DNNMpzATRXUAtUPQhWGxA6mmfze7ATDMlSUkm50GNNDmvUBNOWEhPsqr7m29vxWlA96xkOVcWw5W
tvdRa36nLHDKUzqsppFpgw8Uc3/FdNcLwBQ1OW3l4P0x3yQAqAqkypabPEyBTLF16KlZp8dsY+zZ
0wKvcSJCgQkJSymZJlSUnBcLvHFuiycBlm7kz4gxY8V8Jjhw3zNHx5PX4exwKEFvBFqGNJhKUZto
m4uHD2lviZ2uN9gPMVeF3+W5F5Ftp+SYSKsyMW0vi7qgWpmb76SUQeasWNdD1dKOJ5Tar3oKvHd2
Pftq8BnC1XD4dk1+cQP1JzH7Tk0z2q3fSAlsKeP/NiP7r2TNRsj5/VM4IXRAPquFulNvtnUug4j2
4P3E3TWts4YNwcx2J3KNeddlbynfDoGxn/W1IlxJ+hG3GtXD1enZsnvTtpo4e4hGaWHvnnf6SiZz
jiyU3Lnr2cGP3G7OxalnvtefjPPEr+DrgvOqBeSG5KLKohRqM95yly/GG54PgkbDIM6LFskUybsg
qgQ+nC6ezt3r7jtXN+CD5nKPK4qVA5jm1w1NeFoszd4nJcMakO1KwalJJE04o5Z43w6Tx6Z1v9i6
a7sO8jdIpYcJUFfw2c4HAL3pr6OFqeRaao+AIQY8pgXzHbVrlUXbaMIPQlfsUwHOopugEX8tvAqc
7gyWR6LvkQn+FHsZCyb0p2NV4UmlCQz0OEfWMrphtKjHqqmPYzCUDYHfjENFU52J1s/XDkkxeDtM
LyQiLGHVQ8AyV0tOA/hFhlDHx3sFyVRjEcU9Lix6MG76Y+cDFheTee3Je+wLB4ghNOZ+1DRVzTyX
OYLQ/qUoKxLL+0MKyanjG1IHPHWSTTZJK5bpG4/xZNUSDUKbwR3XAZPN+9Sxq4B1iNVVG1JxIlUO
NN+U32OvH6GaR3XCeGo2bnCzMtNUjL1OUDXqeEZGOK4WB9GmAgKLTdwTYaA13rHTTZh6pxkrpME0
2dmR+yN9qtQvWMztoLfbnm7EyXeDrF+ATzXwWZeYJ6xUDLGj8WgFHk5br9WQdbftI7uasOZUxpqS
uHL3nQJzd2+vBJxiAE8T/iTYFJ8d2XiKpkOHUWpSNEgAAGVeGwEy5B56iBY+etLOsZB72+0ji+9B
p6nGVIDXRGrBCvVGtUaWhQxJu1lW0oSiBmrlA4JerllH9c/Dae3dMDNr8f5yrR+BWK+EF5L86wju
pH8uUCiOTwupZm6ECy18ta7GDDJj+1rfHlFEJAmvbvthr60EIlNAm68mUXgU+h5+7WXGprx0FT7W
n30tGxY387twWpUZk7Dsj9YcPuakAUQYyDfpooiJfMGf61RQ0W0N3Crsfav/muzQjNUhnNYDxr8R
altdVeAxx/yWqU2Ex5H41hRYvZbllvS5bdAZ1yy+Kio4olInUdbF8PnxVkOkWuVe0u4i8K9m9qEE
6rNWFFG/+4zo0nEwONZ7oFfwzmBv7kdP45OBd1M6/aLLjZ38LilExhz02tpo0gFOI7hp6k4MaXmB
2UcfC0ggZFtNYOFnDXUHruYFPYlJwYjs+kMXxXNL6y6ru3+LC/yBeUNv2eTGPhtSNLqhSr6e3gLN
HfJ829PhVe6VjaiXkWAQMdO0Tea+o7vkUEDoJYvi6Y1h7yCl/rc7FnS5878KC1D7mD1t7MU/PV/0
o7V6KHeKaHXa7DSv/mAiy42u/d/wx8IwKfjQukmfqIqF0bwlQ6Ym99SBTUHKfLJZzBAN+kPfmh9L
h04qWqcbdPOOvnjdenZip3MGEvNuGQ3PaahvSNA8QppCbWWOunm2jaREB11ETGi6QaVE8amD2kHF
FcU7mhb5T07FfI9rEwSH7FiE+f+Fr1oiQbcndDBC2Ik4598BJaVnSJQViQcS5avSQWr+22nit7A2
FzPjwwY5f/GUwT0OBSHGPikuxOL0Y8xhZIhDDzre2vHxLgcXuBMmWLMZGno3MhPEz0xKuJkeEgnU
sla8o3tOOoQSTzeObHiYvUCB+ZoTSWgPovVwjNE/9I0Z/xvkeCign636ti+EDLQFg4blrC48DLPa
pyX/zW0JgE+Fr0f/KUWMwVenecFmvPKCXe9FW6BEtHjgWl95Y+RNhYPI7THumfj9hnzOKk6JWNn8
guTj5sqczxeYohAcz7QH9/3eWrxfEMCRn2blKr7nVuCvk+O/lTYWebtv6M0cD0RZbHmpoAHG0Dh2
9y6/CKq+TzzYSj2Sv4kutUhN796cNng/JuIG/ei3pfoOfN04xyKWZHQ1wZ1FoCJFnaa4MH81hg4m
xr+CHAI6SDfdPCpzeCQg1Pwy1XyuDVyzaO2waOp55NiA4QtBLIoVffad3m8uqV9oZEZubNLiqA8x
x/BZg1UZe6+IdUPXX8n+P6nHtqk1kcO7OBSV1sWLOZY+h0fhFPRQ0QOZZ64N11W5GfdgC2IINJf+
gzlc8xwN9y/jWCQJhUU2xEze6VOvup2thjYRb5nxHIdLs+KgGDsc28xyO8nPCuWeNZCxAWbkLRbf
Cg5OURbtOk/1e2gEwE754Ut3JGinFkfmEGM+KakVcX9yxVBrT7kx/ZCKp3yC7EVOmn+VCyJaZYuA
tEbzzN6ZFbVZ5/0ZuJiSaUqM+0le2BsYenuytkjm97bEatJEwNa89s14Wgb0ylUpcTLa6z6YX15X
Zfwz1YRruEQauUHTGYyyRlLOmQdtGPVRMBp/R+DnnYm/ukfImxsddl5QKuqC29xxRmXW9BNdcwOS
H+d7cVM5bBINDEWrWAOf2kUKC0+xjrkLDy23qENKTr7El0mgT3SQwIoXUGZ8DmQSj1JNTrk3Jtcc
ttW9aVvwmAZE623OxGEr2fMpveJNg8yaPzSYMiOFIB/bEBIY19SCB8qC4nh0DeMywM09qNwaCNWY
1Klk7xB3vRIW9arnq8aGqNB9cXmLYDjKHmWYsIOIkifGtzOjdRyTIkn6Ip+0HAeHlWBeW9HuUZUx
Me1LLc0RbX8NCUkleWI3dSOO+A5Uw2XZ8j6JrdIy4en7YGo1V4aMTzdEgJ8ariUjaeyeNTH4Ps+3
34IHSBvBSEDHm0qXsxXmNU+/KmuHEUCDaBhNbndJaZYCn3Vt9WTGofViczgOk0aT5cfaXcUHZQg8
6UWe2oLemaIYnCiEKfELlQD07PGn9LZ7nI5RIuFMtzMrGrL+M6ljUEYc63zDB0hwfIrTwF8gPU2R
orQQDU8YvSQrKkYQPp+ESzaNAzuz6ZJcdofNPXsDLXslINXfmWj/K+r0V6fnREguOYcLaXMbyMez
hCI+aAxqooB4YLOoH72+JzUo8F5oDbVeR7MPfyTWFbd/TIOsaLRScx0tZ6L9FBml/xWXA5pb+V2I
t7nWjSMoL8HtwlKlqjo0ur+U4fBmy8oSMPO0dQQgGJbe7UNyue3nzXt4mXaag79Uvlh/J8TUGABl
0Qfi729dD7qeNpOMvCILs0W0oQ94kyTCtZlFFh5gh4dGgaWElQTS9vvhdHBqezVEMN3KqvjwXF+n
woGIkuDEaR0xrxf8LM0t/3J3o9DvV5ITU3OJF3KdsZK+oE1gCAIheVTyTg5AShORN+gQpa5fW5YL
VWnOy8JhHnlUSTlKnmn08x2tbRQAcMf+cJIQnEp4MYBK8XvkyBAocCjlkxZypHStPc+m9fJKr+5X
zpXW4oP9lu9rdbTGd5waHh4AGCPEpILZSoUQsgMPuAkrBAecO/X4+DYEhfmcXkYkQAsE3ukzgxGI
kGQq1zaLG1c+/YjQOAVrHBBiozXxo3FfIIQ1TiCmYLvEV/Mm84UF5PytMsimsBy/Osk3fI/S9qXh
TECvpepwogVKsSdHs50y17Ps1tSHlD28LvmTFvbxJkFdSrWrFhNtLNW8xXDkihAVwAPHLm88to9z
ssWlArTYL44uZVvZBEFggT2logOz7hNXeV/yWmVcDZiZwW4ceecYcwYEYKgP/UolwRE853z/7a0Y
RJnsyse/MlShSbZ23Nja+wxBV8SA5BXvv73KqAVb8IDI1S8UuIJACL1rF995do9eE+/b9vtEIlpK
U8N150faAPcAt17ryS3hJv5Da/yGN9VVRuC8BdyRGZPzrY2EP8bRbkiog5/1kUrhpT4fbH0s0IGI
5Qh2jmTONB5QoCVkyPGLPCzexDVgLkfXHzcgQgYRN4tqNuuVmyumAsdB6gtxheOl/KhyVFeYdzT3
HIuv4ujhnbGgQt1NvRADb7UpiJt3oeyfnYMEOKZANPfv2yV/Ili0MkUlfzUtmXq+juYcnPbFjXCe
RD7b1/0Lm6E5hBPcmiZfAySO/EVY69rmawRrC+vPx6Ywq2vYCNaGPZQ16v5FQQC9Tai8Kunf4E44
LUNdBsotRIauQs4xQq2F38dzKfo/KpCINaZqByxZCIX/FwzjvvCVgZvlyXDcEn4OKb5pLxSKQEwk
7M5yGTQbWzMH2awFTNGyYn3rk7OlbzGOCTW4byMssfGBEYHB/N+2tWHZFjFosNln1S1gUHqBvaCG
6wvTC1wBfuGzgASwV2IYFMTr2uNo7KepXxWN10y+ucmiW1xMT6SF2x4MqVANgZkKs4v49+gVCGnA
xXciXzbDsGom0VYUK+oASVe/jnIGf+TX2s3QyhB32P+K4NAMV0xVlgQPj5p3b09D8Xi7u2ctzsjB
Peb38OOww69sPy4B+4wsttrsjZBKivU7RwQ8zPXkeCvJyfNuXGlwSOEMRQRLaDm/Ove/NORYr4Re
2ThVRO+jf2IR6vIG/0nyeu79zcqUvG0QR/M8oL0E8YRAbiX42zJ+ZPDq7OgEnQbxWeA616Xn0V7a
6tvGbI9+ueENn5SiR9fWvOTS6g1Iuejdr2tc+ZjJq7mByYokS2fcamAU+Ci4IE2MmixQpLIqiSQL
L9+oL7QN1knDWbsXc/JdMGYbghujBWN1XS1TJ7SHqUrKQ5T0DE0ycYCY0GfU63zqy7SduNwMGWqu
kwkeqqa8OUTAQ3rE1t/ZabKVQRHRpHn8ELGOnpLuUC0Yb273dsKDpIZfMBRnBkBWniuFhqfYgJKD
cXWysWLgXHl7jIhE2RbDCPjGITvDTJyIUCOvhWyckt3mXb91UajQqWiVKK7cPgrC4NShKskTqoJL
sRj+yT3mfyjNtie2O4s1hTs8nIfoicFwAdXLzNkYnBHPuo8CAvi5yjaK5nAU6RzwGwWviTd+vH6M
uqgIWl3J05L6fjqF5UvU/ahCyLQlgwFGr2/WhAFGz2OI4roLUaC/K6pmCrVO54tQMLFXbe378Tne
NMu2CPS7on1wUEHlS51o3pso71uO1tpkPach5aYErOI8998usunwOmbtJ3tgdHdD9SSXdIvqurMm
FpIN9kjtdEWigMpRjxNfRJqlmUyBZ/TAJHT61QOH9XFSvPJ5AZ91JWEZ7x4GLIoWl3+9/s2YPsCv
Y+VRZPi6rD3mzIOIfY6KFA4yAwi9SqTX9bMXq7j+xEY67NafdVRWW0sFr0x1Yj09U5LA2t2BLQ/j
WNTGr0xLMasKxaACuHdta8F4rmYlroLWKP7oiShZ7AJRcOc+qvg/UXr6Mxl57Ajr+peqkflYlkkd
rhQAQTfsEQ569hcs9Flux7Rk/oehR6e4xOx5adZenjuNdEZGie5SKmojNLa9XYK89SrVPPUWI6dd
66oA3H75in6ssZCEE3nD20FF8Fu3UkMEdcxD1hXUm+mpdnEpsEVD6FRyFngFJfsWKdALA/TQUuJH
OInxrYqVedI3wdd1vgnR9TBK344OkbB4gMy5AdqnjIsYCgYPGMEYb/cQ0iNpCzHeniLg65S8W2CM
zK7Ly22m4fUeT0trOmqPsncfgs6qfqJ+eOtBj9V+0HRqNB0zeTtvVggBrugr0PH5KyaJyQbQ2tf7
hSz9cLS05n24u3vubQiLwyUAZ33b6G1s/Y3DUwSCKrqQuLTWP1u3Nbjkv78Q3cRDZGsZ6Supf93d
b+yLgQIQClPpQSeNE3a+NeIfV88XvsVy93Ka2cj9b/Lu6KWawonxMBx6Z8Xs52BY0l7lt6StnI2/
tR8P+xWRjtEzJfBrOwDnAivdOXqzClTs/FcQJSh443Yvq/OCs7HazO87wQ0704muOul+YpiWG91D
w3IcorlRB5Oq0m390Ksf6b1ew/KGwyAAlLPF7OrzeoWli57YqxVw9+Cu/3JTMTuFIWVYT0mmqk3C
e1R2bCKAAgjoKokGxa7/21cNQSQTiU9PFAazA3fm5Jz8Rz3pvC4CAThMNaNbp/0D4IgsL8CD7Tq7
fxJCnvefqeNGpoCX6tXYPJ8uvUoJUnhXF4sNUzPTj0USvJgryzoMAN7pkp8++7CEc6ikV5Fewxv6
g0NMab/KtsE3FuezzVs22FUSR0x3C0qbkqJ1/OgueLFqw5+uWcnZgIWwC/juK44hHMiSJYX+EAjh
Jghfuq4v/2RWnR7Y1hDSXWsFchGmXEQdMD2G9zWmJBSf6ck7Ef4jNmWqExrVTO+biqJl9sZA5UeW
EVzGcj1pySuVwF1gUZXX5wryr5XURbw75E1nvg5nqU/auAnSd0XxfMdDb7NE+otv08ksWzweuJYs
GxWeCVSH9NoY6tLZbAU1z3BPD6bTUllLWZXr/CFg7gv7p+Eq8r9gJJZo6kGd4cDPOVHN1YmXxxIe
xCjdfqGfDzsxTYh/ySMaemLYNWJkBtg/CPi8pS7ml3QFy65YuvQKiEb3qSgZCkWGrKFYfUmCcOoO
S1JrSNASFKo6yDB2vntxplnPMB/uEW4Q2ljIaBt+zGqrI1p/9hJl9HB3PPxfNfsQeHNL5aAm60Yx
vcPsIWKaL3CeOPEsSgEN+MXB82UwSjRZ8XV+7JOpfJ3XMzyN+RIr+24IAsrRszZjCVoielPCnUSs
gKiLnChvxAaxr/tsl8YLeDiOhUI7Bkq9my4/UTonbvd6H5EGBDFQg+Q5eEgzLqPrBwlL3NCVvuh2
SJrsQyWMc4Nwf3SMbgrOnaoCrYZzjee/8VaPxxPe6wopMCQdrFMBb8kTEu2HK3KxRNRPOk1TPz7Y
9E2vqe01m2P51vXf9eQIE7+KE9XnYkPV1eZDhw5u7ZmeTpudvK+Wepw7Q5rODNmzAaiegGiVNA9L
TYrjXMl5KbvLqkMqNVJIBzvLT/XCMpZTjO2MqBBTIwJqqlui5a5FeoTXm9ISeoBvKtlTy9ETXMyD
vEJMUahSYuWO0bKzenAuY2mP1b51y6TgyIARgb3fjyxy0RyL/3KP2eSbWumfcASLTWYtFE6UvMKx
L7zHdTaeEQGjyfNdko7ByCMcHLArlIyqKuxTRGnVPvfNzM+8zUL3CyGOXyAdn4XHly5qXns8qRzj
ZphBHj1kzi3hWHt7flXml9z0KIrsxpIZrjqnanW30tB+Ne+zBpcx4EewBIUY6l4ysmqVIO/WLWpH
kxyit0zyIkrqaCwy+4Wix2f4il7vgCge1O363AMMyMHvNnNyxxWoZ/kppMYn2AmmUXuKkgp98gUy
ZJQ77PU1K4o7XmJ3SaSAvuAg2LG9oCD2QnCPc+ToeHm9vGQJrM8Mj5+Zdxjbkm/2HRXTsd+jG1P5
wq0UaT6gt0VbwuQfSINXiPIT2Y2YsWN2XNV5hBBJm2fPz49RGk6NKIp4XmfLYCoV7rco7BVD87Ub
DErO8UYG2Fqhacy8GEaIRzl/BwqJvo+zEWHUjAWZ3SX0t5zsCkan7ZpOA3Vv0Oh6H6g7QNcecj2h
lWsbctygLviMC+xgkUqlnk+gWfWYVE9xaWTAsRp0hOzK5BPECjVUPnX8jIb1mdBtj97/hansda2f
vgKFfB0s55VVfE39h314mG5pS6QGCYbU74asyFXCxnpgi3wCoHahichpV7TQXVwctKKLlOvhIBBf
EJiKatxHBYkliho+3bsq5b7UMdhw6HKp31h6pDfy+FMT+AeBCx3qXbqjXVMV1VL6P4p83KjfKAJm
rvj724TXDxfdRr8cx/IWg79h9pqIgob2GmSHjn/J+8///MHC1rC230TC4/P8MWUsjoS2W2eb6N9G
hWTXolQdBcaAXoUB4VmLnyqp/2r7i/wIOZEtQJYNW4jBLkn08BWriFrECE06hprR7l6lYok30k83
g/cPaB6QRyezVesxyzl6OMVLH3G2018zjDeXTSDs5De0aquZ3cM55nAPV3BwYJIGonCpx8pYh88T
OrV+ruyBjrJVZpmCGVXL1a9Pk/0M2W6lwVYQeplN5lJ8NSxEyJHWA5CAj6tX6L1XxW+185/xyYFn
LTTjNxEhOe4hI25cgBFUNB8SF9gUSKdvukd+RCqK0hq0VuqEIyXex4Mb1ovPu2a1vRIM7ypakjuy
v9j3zyPUNdtD14ZAz7cvl9g6zGLZVjytfXzFr1wGCAhQ6vYwNT3QLxXNPZbKf5UCQvyV9nqL5N0C
XodZvjVMcQ3AiEA678MYqKAXyqcIxwuklS09XOea5vahxOirw2ZTc/oi5L91fa2XKhrpVlZxlvhA
oOLtxS1M+U2WLv3BSoNbqf3RY1GgcHDv7uVGk5VzpXGVMutyh4AHkvTY9623Zv3pgoM7pUk/TpIM
Z0E6wFYPI+o3G4kbN5xw3n6coo1xYTlN0Yhy2HoCvNFZvPjeO8/+2PaAqoWYzM6PUgsnM9agMhxT
qXKUMw08i9d/3qvgPd5V0fqxRbP4ymSOtVUGingUGP9NVmjQJOlEjZh1ssZw0wOef65Ycnax0lMk
onCNaeILrPh8xHwQgykZPGaYspS8iBtlUhdbwc28Qy6XVlqI6uO8f1xUsHaAT1aicZNGQAvvLoDS
kUa+ESezhDEbZlLLUGDnP1s+hv3gzuS1EbTtPs7xcij5NHP2/h+DH/zpM+mS0Y3HXtkssjVQ5IzR
DHW0s92Q25jNEK2jWBqw8JeL9y/8i0sAATQyAz6aXt5p9rHkKCV5z6LB7mlYnXZM4F2gRm4UtJut
Uje+Fde4I4XoysUwAPxwel90qG6/HLr+okscUGRUcbtvueAnD4Bo1AR1nKdZO9vS38GljKGOv6lh
X7f+0bDZGzP5a3aLKpaT2PQ9n+wiIvcuIuiAmL+bxYO7p/sxBN7dsTG+tGEUzJU2v+VjzuipGBjf
wy3uHjrMSfFwV3lbxlKDR2Feg/NCCJRD4mPDfxqWDkGQwOxK7l75YubdqIxprI4vhAjG5i1l6esO
GwCNUTKe6Glf+FJIk1yGF4ZJM0CneAxDxIg6QwKsycvAbJDSlnIMw9ngIIjdh6bE5LxtctS10RRO
dcRzU9qNWYtTcPts/yDC4svQAPeYP8xe6OwoVePZIiAsKbmU4FBPA0wtgbbcFARh+5k7BWvSzlj3
t0Nd32kOugEzN7EZKs48nqFRgbghzkVzom/iPedbhDNeGkIlm4W+z0BYdIteIBBA6kX6SJu97pAW
VhV4vFRXiQaPe2QaWG2BxWi9ZpetPCIqFPG2v/cO4t21TT/JXvbABgdI/5FsFOJaLWfi0xzUEaFn
Jiz5B6WOTFGo7vtCxVVfZGDH74pM80r1QQFjJRt3DZ9qv+u5IMwtkMlHvPMRbYMUexgKn/58nmWb
jgqdPwsZs0un3GQ2jGvlrf5JCbDPBclkb8WidEpkrwPqeVaRPuuhES+O5NrDMeBiGCpxthnpV1Y3
A+GKt1V2SP/DN1TXh5rMr/8islucg1HYWrMtj7FlxtZRpXuQ4YB4JKrGBLRBcvz0ozmgX3oisCFV
QU0XR3q1d/kEwwp2kTgL1NNsg2HssCRCTvAGVYzcPz6dWrN8y7/KuoQ63CnNXXUdF/7xnZCspsBy
TWOvWXfmqb9UrJJypX+w39IDWDgV1nPn94FjYI1KR7ARnBJk95OPqG3X+E2Aa1mh3VYDu92qQS8X
EUHr2Xj2/r7oxqEPRH0B/wSSmeo3CcsOk8AGHsSI9vyGMl1IVvVqJH3MxQELd4KMkvSUvVagWYeW
0q5IbDng8ClaPtvLKeJ10pCNrZp/obyB8cT+Gjx6JV9p6W7zJBSJzis/kusoWQI5GlwCNc4m7rHE
3SMhTnKPRSunYoAIhTZkoycLcFc/P76SXr0tM7x3nL6Rlbm2w+n1/uUAMIbiokpu5q2/k/XPZiwI
RPNJ/S2enoWadkjmyFD5DUFHIqweJ5KDVqo29IBFQSdXEPlkCQEMu1bjImJHhL4UWAQnOr1s4qvO
f+/pX7VL2TTuwVoR5vjO/08nPUt2S6Tgs28bjdVoBjHLN1d+TVpSm0IPEHq4q1XNsGQmJXh94C7h
OK4Y+gFCD37bnYMHvV1Q9eh7FhqT9mGmxkhcjs9Mr0SX5UXUv7JIZ7C20okYoH557z8uMLgHwhqc
O39vsu7Sxme/a486nR2R7hHToE+BjryuuIrnqSdHs4eL3HtlvGVw+k43C5ZUPBchCuaIKKThN5F5
bXVdARQAUh+5aITNLFeqhrXWlBN699/x2CtA8IpFmjkbmypDeNaVoN8F6buRCfcwCkSxduTOzvGW
8LRr7G7zYYwsDfeV85XRPOnFsmqM40Y7OjQcseLYrjeTpMhnac61Ku480rbLH5iGffP//DoO9vP4
lTciNPjpXUlTgivl8OXn6u+0KFCs0AT53HaGa3wwyq5ivCFuBlQNxrcilOAwPY7LfFFGUQrM3zAB
cIHEs7i1mC7eHLbgP8HHf6uVt+6E3LariZDELvBqscqrFs70+FJ6ex6xEcYI5uAPK6+2A+wGtGEl
vJM35bYADfpOicfqWxoGcoCY6btiGSWKbUbDp6tBk03iO8sxxZzjtfE3GfOxmp9mfarW66T/8LfT
RXo2XWpP6wLHEQZw7x13NzazTFtQ04WJ0x+xxYR++e6i30QRqg+7a089kLzd+y2yS4akzuYJKlgp
BF7kzEF4JvCtxfoWJ9gDCnXtLql+wrZ14vIPB2/HlJSVrrysVI6Fwly0I59zqJ9lEqawjOeXlCiM
xzVLij3TQnZnOXLnQhWV9QTt/vOLIHZvcMCK2qjbJMEIU4D63uLrNecILkFEi3MDD0RHM5/c++C0
1kiDiHR7HcQ2/NbqL7Iz0FMeAG6YpQSYBpouIORJidqXGL2MZvVTn+D+IGyChW71K+dCWtA0ZZc4
IjR0eVdZQWSsTm2kLo/YwYbzn/lEBsd/zDUgNeIwgoRY9iX+XQworT4ndIKKRAASwUmVDMT7zoXN
k6GWmOyVGMnqcFaRTdcr36Xs3cvL1XlzYZ6z3Cuzue4LuoVbMgNeuPWpKY8bHJlLH71Q0sz2tWKx
0J9jD3l63TLNiV6TLBsm+lpLO3OLzkJmhuP2xLwSexYIRcRQlXrV87y/iMbmbfkVR6j+bl61Jsh7
VLM1CrEVoTKtfwbEU9QaZoPpSYMEH+putsKVdTCJyt0+IpX34RHr2ZNJmYAVHA+QmUs1h86cXjw4
UGM+EhIV4lFoll7lspLnrf62lB0lkCddBMYyh4Q5ZH2ZdOBt2UAhLLF13tOxyuftis91flUkyvax
DIMkBSdVNvdPr/jhGPnbvjkED3xNFR83MQXuLoHB7wgE7J9L3RkO/ViKzvKO5wbcGFNI9xrYBtU1
kNplQz+D6V7zo0KcyAgNNuYuRzgcGLN++TMLdNJ9f8VhTnsKIazddjrxTTC2i+O9MeFG+VGsweI6
qC6nX+Vc3CIYEkGtrvbXERMJ2udr55by8K4HVXm/6SieTpSRs1sN+uXMhknGJ2gI1gQYhKF2mjF6
WBWuUANq1GEeVQvJLCKzSBraJ/YV7MY4vrWStzSjdBMswbeKUxPLP2kL8hqR6IwOuigAVkRbvGhy
AnY53tV6tvEOd9w3vicGKCEWpTOa7PA6MBe2MJKRxdfoSdiecI5jcUOPNhCQn05eONo8eSKjBbhZ
L8bX+P1187rOKG1aWJ2xNyx3uRfs5ks6YPF4K17A2BqGU9OpFzoFy1R90se+4uWT+nZCz1qF/xqp
cf3hTS+HDxi2Nneq77TfB2wphO/YmJlSgj1mxtN8ODmQ9s9YQ2t1+gxvC3vdMG0FZXFpwjtriRbP
RUBxygPk1ky+tYvV1PlzQ6yXdXKoyhhcV5W5kEa9IdzMxxMEdDFuQZhdJPeNE9DTNEApbNI1r1Rj
1RWLnvtS5Z6vWY7SmH1HeTIgo3abXHj3Bc7H+ffE7jtsRtPA0BeyTErtdMRdFgHj0O1Pt3KMJBKj
A+TcmMkq9IkK+aLPY6qo4aPQY1E4WB1I053FaNpDIsygpnsq8fbeIRTfANS95zGB08Drl8FeccQM
rbwpa93Sk5pGvH/44DxwfYo03k6BrxrWVxZ9MCOCyGboNMyAsW79tRUKU4GtlUyq8I4j5Me43G6f
q/ck/Iw6Ix0EeATNM/2jAj7bW4XoA5va1oPwiRVP3KglPbcgqsIeyIbsrZm4YPpoV8UoqqdW/Kkf
W/3+pB0fctol+qJ5hLKlTQjtU0ZdX12bZjLrl9KF4jUsSPQ+9xPONk4wfHC69C9+j+wMLCBDNZ93
yABcX2gJ5RqY61rblBufdhsEPjVSq8VyatYSDIOwhRVm7C7PU5DHKwDJqN9TX9i2uLXoz2t7GrfU
jf+A7pYNI0dIQ2cvcWbG1s0IKqqZItPzorYB/odNb0Sq6vB+giTVQehkDFsmFtxQKwt+jOl1VJFA
B6FcHrZbW7eOusYBXnl0teW3OJ49isFm0RMWvP9upvhgp1XeF3QL0/sB+Gb3uYCMaHwM1KvVwSBx
0nCmbg6oT0Df2P2yHYcgTqex1JDnO2TSx5kw+yA28ZLuAJUNHXDF+2xWmWDId4NkIjp0BODbDhU0
NZrG81r3Hnuzl9Uwk656wb9x1CCSZOCd17c0R+P0YAKpmCroAS7CEBp++BXGplgwk5Z1WoFw8tmG
wE1BXs/XUVFs3RduGCJIDReiAoEdx3emyRd0UBk5lQICUmmaxl2VGdZBlTDrPsw9Mhs63JhFmKTM
vNpzD/1ZsAm9RKL+q9N2ZV3RnklzY1xYY+v7Lx75h88Naj7P28OdsPdSxdJy9XQxaA+D8tf7Hf07
r5cOoQFfhcanYr9u2Ec6cFrOYgiyIhRrQZmjotU0YHylyoPkm+vnSSCQdfzxZLSsbJ9NxDzqdsIN
qq/52cJ/Cel8fZ+GaAC+Ue2ShBeqGCrbfM3+0WXe39z0TTAkwF14P5pAutHqdRuXl0npRoMhmkzQ
9et7+TYW7nb2r2lEXx3BFuJeQQnQai0XCFwg/HfaSsy8Z5bPAuKQw3KSF4aiz/1TJMQAVHuQyTeQ
1+wXLzu8vR6xznzBCuFGp0orA/inm0g9j4CTr+k4Xfzp64OohD1X/Btrxlmh6oHLO6fRTfl51hc6
Bl+wI0GI1NrraRXsdOFakWZvqqq6fPxA/pi4ywH1feEtXfCOLv6W1cBHCTOB39A3vrSISwpKxefS
0ugHS7t8E/Ls4TW3jPDZskVPxWf9WUf3AoP+uisLMWGrOXL2dTuJlJGWk8rSuatNiT0/bn0Bhc99
WvcGxnh4RNtIKI1h2dEAJKQt+rifx/45CKTPqZGQvU4f3kq8vU4t1PVqePq0qdNSf6KdqfVN5OEX
KvuS3/H6tT8nnIC3YRs7mFCcoSi7UYw6mxZF9Lvha4L8NZnpz0giFDtsR7MxVx9XQYFRkB/mzHi4
KWPcyF6/wwhqvL8fvDZ1FsmUYeWquwpNO2cwXMgYtCJbGnIeBONGN+KFRj5GSTKJ2SrtrN6beAT3
PnfAuzj47l6zMtmcz8bIg5TSTKoWFl1C4P7cUBdIutm06XWusCrTb60rCHguLHAf7onf++460zaf
va6DAEnHbt4GlFNeazJtMNkPWGXYL5C4QEG/igfbKP+ZIzOQxKxyZaK6+fyDnCwHOIjS2TmNFkKL
EG+1Mr+3xWYbYLl9+BCDOillpSqkCsjObYGG9xZ2Z1EvvLLPPMhQI+Je60Dq4kXNa90PshUhLinN
io5dUiNhr4FoqaDRvN8S7T43HH4QsZ9HS1i3lWgEfgaRvzB64DfSoDIxjcBW9wSt29tlk+abO9W5
EQqW2a7dJJ0eicY08H83WpBhFwQSMFgKeAZmWLEdSNfMQTfx9HucLlUTfHW2ecMjJ2ir0Kk11J0d
FfrV9HH6nc0pgg87WJpXi8OaOX+sFRhMQwyevN8HRzlGvbF+G2Av1uOnLCebNs/Z8qfLy0UEOeUw
NjDVW+w1fYEp6WB5OCXclzqA0yQO9Euf0UpGKf3c79keca+hIvD/sU/qogBmJk/FbmpY9MNCbvPW
hPwDyKxpFUAUBrzAeBInJtF4fNB98E8qoWxc8zwYMCqj2DfQu/040IYrBT8kJ0FuHzj7pgg4/lXm
b40ph29/p/t6uqkS/zMCnheMBHq4+9tsPebDBGoIpqtfM85rN+U5sSuZio5zdHuYOh5YHfqeGgde
s5qOY2H7QPWJpBSjACv4dWIk9jRk0rPzJvFCDsx0xo5pFXz9pBYoPBdu1OW/8aFka5oiMA+nWgoc
rl3ocWnkBKH0UGgvKiI45F5OIz+rKRUEVvYZPjKqe7u3pZo1c4pconSQR9U4vF1oJsgLJWOXcC83
OtcBUbC4Jo4CyXs/2tCv9oexjBLQbJrsCoift21EjBczHpJ729m6ThKQSap6P0RmGGvE4p2FHCIt
cffMQO2nR010BozAbtVqmqSA/bJ2DHJorwIbzoI4HiZTOjl3WfiWeCYFrS4GF1JYwUKlbm0bvXKi
aJCYAiOzM3RaS4V4v0ruZfPG6Pe+IAz/Gn/AAmjmcU1tKVkKsQ5G8aHIoixZ4ggwXWAaAS1zY38K
9/yPdyb0M0wMv6TJ9ev+EfgvzE+zNUGHNyH43m7Xs1m+frFPXzcToDezPrdxcRMML0YfvAgyKSsf
kEOvnTU1NAGtVjPtKZrZ6okpwigC9BTxNJEUqas4h0lGnyfXrQcJfXww7MPPzhvNjg8dFe0SIsl2
3yoekaNhRv4LMXSgNyVR8cads7YwdlzxMk6Jwik9WvHxolz1dDbZxt2iTf/l7m56i/Gz5fQ/eX9X
LDH9wng77oW7+nDTkDnzIFbnSg0b9JYWvswkagx5Tu+sYPbfdyZtqQQRwWPje+LkIJkzTXlZiccF
klfNW8OFdzfahk/VHwrHGujCBbem5Eut+MAcdUY2JN0dysd/6QyY6TMwK6GbClGK2w2Wk4Ka7U7g
vqE30iRRYXaXouSPMdKO6+sR3kVnRpEw6GxAIJ+G4mjNviripXxT/yRybbrEXLw2R4MIFpTaWmo0
v8Ez55991KAV4BGwAJSRSorKEykqhihS9Za6Fl6VjYTl5coCqYfvzd945RWTNztHScWyAYD2yvIA
BeGTu1aPLObuMbDtSrhdnZQudKBf6YRrN3j6/aWia8WhSrve7FDlsY5w9ATUVTEb3nsUromUWaCr
kKfCi+Xy4fxRkzbdU+OqJHFOMAkzAJcQyoZf1mNg8c3polZ1hwDurmYNI69Yi+H92jqi2pho9iyn
q2bH7mRpGQqq0fyZ57pCn7fbKY3IiRmE1b/CcRHdzReHTyTWmACHHODBWJp9z0Rh1HSz5frj0om7
XSSeCmvfytMBFk+wLEjn/iZ5s0B9rabIamwFnq9x6SBvxxrQSTsPRKmoSAg1takiLLT8mrLr+pm4
qeB3tW32RBGVVd4p2zmlhMOVI7yWITDh3I858jxxJwoA1KZjUVuAwIeAWTbuEM4ObjaPm0t3HROV
FxERjyH2zL42tjDDrx9ywp7iGHhQILiO9Rb6jV+ZqfeU52wfKe0MmS8C+GjwuVvj1ghNK5wdWuyp
IUimrAUIJul3TOqFwTUpBHiyFOmGJWk4uDbzSQolVc3tu1CFDYAeUW/ZApManMEH09tv2ml3qTzM
xbD3keoQDEzPUvMn5cubmaS1gU0McLA+qalstpEL7ILBBzcbDl7r6HE0WbL8eGsU9llIO5d9rnOX
WYMIAuoL1R49hvlykKQVP83yniqYFvBm/gDfwCWV9tZpsAbFZz7xLFjyn4up9ySIS9TzkRzekBSM
JBCMCY4ddOqQBVyo8Nxw3loiw2vNgb71xIVluTxECtbUziryMDRYSFpSP/A6zgIJn4QI74UenyI1
WG8HdC4mtXl8UJHOEfo3P/geELsWdfuQPjMrMc+HJf8EwNkJx9vH8Z71b22robJkQ/CKCJ5Eczce
DGk15SIQaUbkO1gknqX/4giTYRorzn82lDRGJ3vFoWvK6AEj42BsgdZ/ijnItUMRdGZkL3TpiEw+
n89EwvLWfJ64/M5cd6KJ4YuZs+ljm5oAhBCt3w7K/13cXNnYWbOH6oIgN3cQYyD3xQns32/2/zVL
GaVtYPskNmBThx+jFY9c3e7mKYpFNK8y7l8zbfBvy3go0RtIhxyEcp3S4sQ3x/MRYMP8Or4VDZcG
Qb+OcZgGvPIh0k1SYylsSwgp285+EBsrDRoRpvron0a29vigZ83Heh20SgKWUYNV95MnPJ5DTbn2
c+jKL4jbggDxAbVfD/M11WHC9Up90q/4P0CshidAK/cuS7JRyNvPjLl0meQXGEn7Cip4mrujcRlf
gOO7rS2JMM3a6p9behVBGJ1EriCxcncdS3qWWPVueqoKRGb9yPITlosLyFLC5AF0z0Otmb4VdJmt
UlsrJc4HF9zkh9Zi/XDj2zGmhJdmJ819Ece8BwaWJPxDHEWh28CWtKMUw2C2d6ZYPvYwemvRtDtT
Thb96vc2Nq4GvGqhy76GMYnL1eVkOz58MIN5AaujByd7711MbTD9kJshuBJ6v7+zjW8hEn4+Cvwq
7r5yBirnDqSXMCVQnlLnlFYEEAEQLK9NqBj/TWcftttn+ul4wN79l/twmM64J4fLGwy/V/DLlfrF
0OUaissdlREWnKNhj3EmGN0Vbk51HRfRGzfjeAqmllRHPMoll4TB+BCYthq5a+7HvLQLKD2ZxSI4
ZNBB/JoLs+bMitBfKvYba/A1RQnniEz4JTAh6xluiTreyKyGtJaYIqmPEDSfoadtta8JpVdVTjmq
e5SLiRYTnCsW0Wwk3u9ThPVYlJ+rYLWd2CYkkTnpP/kfgdJ9pSowdF8mzIsb6awFQnNS6E/eQMz6
Kl5SDBBeN948Lqiu1eS2y4ZSAjmJ7neh2B+vQ5C4FiFkp/pB+R0CtdZO71RCkbKvC/YhZ/Pdwjeu
79puS9hW6qO/s29VioC3H6gc/WPpfJS4RMCkrUU9Ulw2BvTFzya+scF3pkw6lnooZ9P8P0wuuPdT
XxmhUb3BXtRMx8GqW+H7H4C53/3xUniPdAxJtHAvpVTrv5ZQ981rwhRKOC/AYcxg1bsluY2S8QL/
VbNPuiyrfeZ1FGW2j4D5qT/hUvnLydDUC0K2Zi+6Bvxc98eofoorolxW+nVSrc/S/CXE8lQDVCyo
Z6xrS9r0L35Y4r4WAkjBsS4F97ZphAv7eIQIoCxWRDOz9PSi4QLzyMRYqM7HUaJZvvL28Zx4pcUw
XyM1x6RqG5OYWx2Qy0cHCVuzM93sSZGKJXaSlxB1wC02abRnqCVQRrgCYVpSi4iXdw4e285gnQAF
hQmnsS/xTOz6U/ASbImNGPUVNyDH4D91dF+aibDjUOALCaOVjOW/SCeoJlnOOxnkGzDNGCn2IX9J
Qmlv47MpLiSbYiF2bKfH+fzbifuNoHttWcPXZMXQJZzycbDW5W+ei0OGdemRDglmL/juACufFzgu
nHMHkZ/QIqtat3qOrCsqniUvgLejor01Y6uyNPglnz8CmKvfnOk9fNMCZTG+cJ2jYVbSbfpm8D1U
2AfqaXnKFMg6yt587xJAahkcyV07KKe2WmrRN6DCyphvc8Bk+CDZrjBTNYqf0wwJ1jOdSvg/P6LO
ljGMirpOROYVT8zaiqC7MH/s+5G1hS/rf5MdPsrFlwSvIj3m7wHKHsxGUfrh9wYSGerWYkYKXyM/
iUr2p0jwBnxQHX+e5Xc3dp1qoaV5TJN0ltXtNIJlCnGLnoxi9mLJiR8LAaHkGYNodklkzVWhrb9n
ZmI+yDyNtdXLsja6utHvWXszi2UyQzC1F9RtBcmMXuQsQitPPmHV/bIc1RJGSdOMTYJpCmncFC3x
0DIlZyHy1YkV9Msff/B49ASfbiqtf36awaBW69iRWWyY/AFB+lGQPuZq2cO38b8S3OnGvhXU9EJq
UT6Zqr5QksqTRY0Gw62hYOpiEsdSrNUYctEKwDTSSTWIPwAeW58TDd/3oo8Sar5W9EExvgi8Vo7a
nai2aGgIOFeGKvnSkMod00GpE6yeRO6xSTZkZPdOuYGmpNsnxZcJ6PC1JQiV0wfpoYPI0CXoyB3k
rNTf3Wwo+2C7fmhVFKzk/fa4lrPgeQ2HAVcqmrPs//1XnrGrtSl218Mj0jLdHb1/okuPJUJzOMzX
i61OZuD/uiWw0kwMzsdfIm5k3QYZFZdqybO27VxE2qJJJ36qSQNEaBxellVsFBhlGqRKyhiDbmKZ
aBEfBAHVoGFhWOI23QkLZMrvIkyRXtdRFeHbxTGNemx98QJ285dH0c4kg5ocyjTIdqs3hYlUaCCI
+0RrZRZDbrU1ijUU1Pv/P7g4u2YoXfIsJHXnoSfQBD44E3Fk1BHCrSlw5/5H0PG6EwLpsLO3Zynr
k9PWxFxjCl4FC2Ly/TkQOC21f4jXpH+liSXDej+35e1L2ieFlOn1ZpkePmnJueABAc0sJp69+V+q
7C8oX2GPhcQY7VsL+DUvAO0zKT+4w1vnMFNymbLyeaZEgY61Ygk790R9d3tPJtcoiM4DnA6SjSod
eQPB/W7NwgKb5AZd+bxZfPWAL1a8V7v6AWR8f3WMY1Lkez6m42C8gKH+XY9mlfHOhDDHzZSTAru4
4PUQpRXRFtgROjNnue/znPcdBxHPOuuDdWaI8rN3VIdOza0WuqjFAosBI7UAZJmXySa0lwDKseel
oqqFllG6bqx2hKHYszFIQAXuPte1BlD0DLR9lS3TK7SxJLau7rhRytDaI3NgYakh4NNI0e6gxuCv
8JTrVxe8/Zom0r6DeLsPbxN+K1uPaYfd6+ItDSc89MAglbLI7oaYdFkaZysU5CbcDY1bS9QLRdns
iOIfcdP1wx4QA5AmLNq6qldXoBMVEo0lLQI77Fv2v3h2la9bGw+5gJYXWZSn9t21oUA7RwOKkNCv
soRCtP2pvREnVhxEu2S+mGWqFVNepiNn1KwQMFUauspo8kgImIH/fOSlrkEKLrD7HtWshOzIvKUL
ipbwDn+FnVzNxMV83YAyb3sNBegcpy2DAQ+2dWQBOIhs/xjyI8yzOAu3zP5CG1Q8JiQgKkm+sN/Q
ak8Fzfek3j6xlsl28AA15OK2sfBx6ycRCHEGq/WGgyMvX9cG3O0Xlp9Ku83pQTdjACbqYdNLCZz3
s94MvHjGZ3c9LDaNA6aP+y/P3BeSVrrPhur9avKRJjJ567dzmdbPZ7bqr06eTrvpuT2kcfs7/2LK
i46C7EaFxStsNVS4Od1Bbr7358YzVnMm1BOE+rH+B64b2Vv68wnhzsRTL4TZPjnWhhC6gP/163nh
25aR2X5WhGGjSO4/kXJgaHFMOpsf++2qQRalASvsGAKD5mcrSVBJAEt+ffn5dJshmNFXUtkUD95y
fWvetU0wR6FdcdAotfF4bmnI+ZBaNfzxv7luxsz3FQPYslpq/9jACkBtZ1QiwwF0G896bmhb+hyR
2IZpAwOFdxeRRzbT9fxtjqHSkKr09Ik7pElRDjiKsU4WJdXu32ydI/i5UPr+ipdI8GRYxM7LH8ho
tnEhBQy+yuacrCyVI7UD7mlKvIP2dGiund+OO86qGJzCTQ/SHDVAkrp34IrmZgpBQRX5gYl8jg0k
sjoycoOt/MSAwjstYpnCCcxCVBCSxNJOi/XmVSS1u1yvVxRYaab23fZVAU1IzA0DCo3yVREdMfm5
/b6HOkOsOQ2SLBCQCvyGyFNY4ZqsGvwI63LfGTzzw0ccUTP3loLZiY9dvpKnR9+bKbw03mpmO2r6
aXf7Mklv7YTzo9jdjzR8CMKn7h2k9a2bPw1rdy6U6a5xAXD8Xeom2d2XrtrREUoVFHEiV2Caiw5O
EkElmFYc1uYGkslN3yeBlf0RIk0gdjSe+QpB/ODp6ZqeIl1UiLZJ0+CaQ3Tj4zQ2WhSR0x6A1spH
Nfnqjf5GdNfdt6M1mHKEUM72dlym6JM9XS7jE5x4jsaV3CbEX83UPVUeLhsEYLrQi7daQvWV7z0/
YDLZcGv8ERchJw7Z3IE5rNIG5w0MNuZ0TLG6u8LSys7yrGRDCtMAyjeYPTcYIwrt5RYSWOlSo7JU
gN5gAUVQoXrIULbkRnyfauASo3b6MZ1E+0F4bshFgg59Ne2RnAn8ChYRcRAq6MmgNZyK5VhAbU9F
MyabbubwCP+pJiYBP/UTFwA8zCCYl8Sywa/NoIYPYMb3U2vwwJl6uMBhbePPKcFgzzkHKLFadf4C
O0EuX+1AjhefyMUxFTCfLHvLkLZziHbD6tQvN7u1T6M5AQIqAC+CddN94fM6xrPuNAbWwb0Gwuej
Ph9WY/3uhYIL+P4BvIuCs4dAUqsgFqaPriwKWzTmpQWLvaf0mJTh4Ol7OaJuwvqemhQs3NuNv/T8
eH/yn0+uCFUDB4YpVQzye61vWo26s70MgpQcWe7gJ6+kA0kMZ4G6BqOoVYOV97GUMSWpEJSlXwUc
h5o2pyqKA6iOn8ihPmJ8JxnhkFpFLrZV7fbBMt3xnc8H2Ktefo/tqFv3KsRe+NeeG/ACBQSnmMGm
MZWEnQhTNy78n1AE+wKsnm4a5H7x+YnvxF7svVkR4aQK9ykUv+Fn806w3yllMWDLtXoN+MSfB6G/
3SHpTsYsz7VTVplGStS6GpLsAUcgvl7XOu5UJbFG3b89hed/m3tJMBf+/T5tYiVuicTmIRtKvKRE
CLhMBO9Mp6HPu/H3mo88oCtVT9AFwYzRii80dXdAWSXpHc+QJi3iZtEb7vA3kJSr7hZtaArWI7Bk
6ka7dyMWFNISI8xjM9RGMduOlCfuCISkkWwtoJkNmxQUTKuhcQbKbHeooGj721u4g9mOs21w3Uk9
C8js0OZ3AczdnTbd8LHJ+oes41jsyuQN+O7oQ6JwjG5Efs79qhuOhIWjj2OIU40iP4jnbXPboDWL
63jGuHrQkOIZh/baAQ4VChoV6bSBhUs7leL8+GbRJPmRX1ZtnSGSD/kRbZjRX5BefyFV+9G7CyX3
1l/e1LP6Ujk7tL+GwpuJPwtQN1cEZ+C1q2mSm6cXqmcjziaTRjb9jv3QGBmItQQi2o0Q2MO66wrP
Ok/F3QiQcNdZB3YXnbDvAiI4uLWVZxMEV1b7WW4nQHQKxnCAQ9SGb4lp4Q++/H4IKDKWFPwPYIo2
g02JCZerP7DKEJhoXuSLilEa+bWyltH+V+ogBiIGdZUg5WSVsYrtc6nio56pChjQy6+n3DKpHgYc
TDhEb97MUYgkHWeQkWaxosJOV4nRSAl2BfyKORhVwEbi4+kaB7XTfTfHMfNaDT3tBvlhwKwz27O8
5rhcOV4KIZwA6TtPUEXpQytykr8VFLoLN1rD1X1+oPZW/0634McZ+wr37p33sJg/NnrtiFz37YNk
mtWTeRXvVyJUGHoMQx1PltTSENdhxl04EHFzkhyk4CaFZUeHouCHwrrACEzBujIEJbIuto/B4jfC
v3FnAF9fvQjOAFBhSWWY/ow1Rz3Zesx7srI5eVFNsU/sz9xxp/tGE1GLN2H6TIu72UULyDZcPCbI
gDiALXTY/cTr+qVEnELjFB8599S6cjtksUKQFK0p4+y6mXEBiLroH+dtjEnEqsEQ307KSn4n4zll
PlBd+2lAeBx0SYdXMHOiOM6OJDwJdS4X8yCwG35HL7WCG7r3udjzu1LVgZ4Du8sPblj00jfosnUp
XbId7MpBn8Ceor0K/QIzuFylNUQYDe8wJdh9NxztEvSWo76dviasMmjPbP/TaaRnzj/dwwb9naj+
VXo04lqi7ov1QhzFVoHSbVGMAhm5aGqFlz2c315/6REgP5EqQOHxxB4u1Qe8+t+p97P2xEotkg9P
1WEgAjAi2ERR0WKYEM0WjhA3vZ7WHppf95g6DTFOtbuM3t4SfxCu5i33VRpER7SWVAjaK2Q9A7F+
/WGfK9IvU66W2LliKUQJtKEfCzdRNlIdOgMqw4tnRuUwxyz1trKVDSrSxn2H2j+53+DAQ98CYSKD
Eyi3Cr/qFU8i2FX/nrLwLPCpdT8zmt+Md0yisAkR+bLBWnabJLgUtYDuPMai5CUlmoLE6TWFHf6F
Qf0teoy/jiKC36EqhZ+S2omtMnrrdiMxfjtetLFqdecus1iRapkq2LgM7Af2BWm2Jj4tLER6C0sP
azzL+jn6Gi/OHhBh9edluGNV9MyY5w9hnJ0iPKfdb5mvqaaoPS4v3dO8CATtnFmqKuDvKi2GuPVO
80XxigFk0oCLRZ6fh8ABXR/xb0GoR4RPwvZMVBqyD8JbF7ahRafxU45DfWdJ8Nff7KQAMX16Zkc5
T7MCjxnGO4Z0JR41Odl92TiA0MQWGzyQrLlr7zEcmx8zNzgXnjKTVXN0LuckveILh8TjmVHNVjC/
WNHLUPh9xp0FWjE2C3K9DpEKZARh8SG3AHWYFdXHPBArPQJkWQax+uyHcYQ/xu8P3yvVZ/VhB3WT
Py7RqaamNXJYIO+tFwBAX8AMOKTZhAlr529IEpIGU3LAC16Z3klDmxFHpG4QLJL/B6Wix+DphwSY
gRf1evstFSitxKeixSGHL9bcx2q6UwAnkvxzc3STG6o7xJtrB/I5/POLSHFv3RKlc6MXX5aSojWV
PKynbJAuT8bOxHL/OD/vQUUuFv9J+jYpymousbYOOf/leGrkvULUPUQiZrQG9PF63n4oyHNwEd0N
CXvj1Xwa5I+TVKFLwCSxE92Hn+jPVWjwvxWwdcfrKEbA65wvgaU4bjDIXXXeakXYgbAj2fFJ5g8S
6kZTKFs8Laa+3NC1P1W9ezKjhRsbbq09tVN3LkAVpg1w9kaY3M+O9P6ZSIFEZwGaSXSYed9Pk+1d
Fc5SwIqCFWnFY6p/Wpw5q6K3z2CwGlCLjWi+tJ+5j6RwEEjAo06KUvVrlJnr+LOUhjwMyYLZPW0a
54OKpvmC4OazBLDmFACzhNTecWVIzp4ZYCEVl4dT7B/ele4MK6agBfCW6/AEmQVnkFeZk08FSLap
gQBXPAXlQ0MdK3UmrRZQs0hQPiO6k/Y0ONeZMUKGCOeiUovxG8qCSPbJyipY621/Ua8GqJPewrBS
zMP/SVmzswnH6zwjsKkdI4TfnN5ulmrloKwoGhrnnMVzH7DZ/rs+TS8JGxL0dJ2BHv8Rf2BafrfS
zWkpQ2tm8F6T6vARzTsU+xegSan8Yorik3ttsdHalSbLnStP1IUrEn4eIrE2yznlHsTo72ftCoJe
uYcIopZHrsB9j1THfhPxVX1g9oRT/XgwNh+24FFhLeJIZw9YGTAFDXvZa9bWjBcCzy4PJVdRl4Zo
s66ow7F08U5xfc6xbaz4lZFOOduKh4TFzavE1NxuNshqYVKfDKqFu0s5+OAxDstvvIaDEf0lO4Pj
G5AK75Xx7zcoxIM9Lc7IiSUDp0gop8/H89IfZiRVnqNWQqIjsE7hEuJ2z+iY+jC8hudfZJfLJA/W
8B9VKg5KMhusdLpVfdNmC9DTOaoWQrkgLoYdaa7gcSFOmRGmI9xutzX8BHVtox88JU0IW6l//adX
DxvsyQY98Zqf/vI1cnhE+Na/QGh6BCY0oEN3c197OlmPH+QbsOrXquBklsVIvyI9dWY2LstaEy5P
ofcHNRD2SAxof2irW23ETjjd5z9sM2CfqCIoQPwobXraiR8nM5hAI3yR52LUl/FEQq+hsW+A4Ek0
06Uglv13o4meDQBucbr4KvnagtGX+sSpEtKjmX7Ip02PGit0Ad/jNi5jMzgb6BGlpD44RiHrughl
XXnb1ABAHiXxdo3R7rekyl8a+M1iVxYrgN6pbm9nUPRB/+MDt/29uAsU0rs6Mjc5WMdw12FaZcFg
6GYMp/Eqz+0e2yN0dGbavuMG9Uq3l3A5TkIWXIkmlP+6DV5aJ3fXEefkGOHKl8PwQjnCZU1fmpFn
hXuP1H0laIR6iGrmQPRxtfihhpVrpvglgcvgM/V9DSKXNCs3fumWs5XgkwLurU2QcDevlyZr2KBb
ipKEdfy1woIeaawwccpBoWT7G7x1KnueUdO1Wb7VQGAdz0N/YVmx1Lo4I8R3K98E+qatO94vJpvi
yhyJcf76HjLeF0fBKTVf2GPEq+qRT8SaJIT69P9/kk0XmWR0qETzImIyGG8XNkhJr/MytPF/jNNQ
7zWu/CTInw1pYA1ahRiOWg8OQxUpFW2wRJqPekiiOyxvWWTIC6QwFJiRMtsSGwnZn1qLFZhkQayr
SfcB+bZaPIXJdV5DDb/Ava8YkNneKP6GzIC/2DY7FZI0D0EYEMUcRX5+s91BUGX9K/j1DhYHzb5j
dd5sPsD3ISpDRz8PY5EKNqknDxk0kC5GFxGGusDU0bCT5cmnNWkU9L6sEH7mfCVtlnHQvbpfZXdO
0MJj8k3ckeidWRU3KNAJylXSvv8ERWPGZx+Hf9xPVhrU9ijnTdqMEHR2XvEsinHnihA1slQphPtf
jrFtyMnoJOkfl6rRwhB6CMlToNAOGR5lTZ9yDFevbZz0h8ACoF/0uj4Sbcmv2FWiohNm6qBXXwNd
VZK//8649F7MkayEOwTdUHFRUKvGDb40PLd5TQcXBJOQBijiBLY5cXwgI295GJW9rupVFgJdYwtP
f3qbM3XP7IfonIxhIKV6laTz0PFcPm3jYTw/47Tcqyr/WttqnCyENNiPerYm7AzxbWB+0MI3itGH
CEF7EIRbQIZ3R6Lrewzs9N8KekVuzsoBC5q0YaHVOeyEvTSsYfCsEefLvs/iWkNt1BdJJmf+Kipq
KeBnte0/+eJiEQ7YiC3OIwD9G8ZzfvUtwyqX+IeqoJVUz3iX9UkppR8GkJvD2SeBbUhjzQT8EbDt
PL2pw80Ybc/2LaT2AHD6dEmqjtLDwiiSyRwIWO2vdUVWnXYh/opvX+gnOlbRcpVyL5+5E7aDLYDV
gtXsZyH4zVUS61v4wTXmIct+B2c3w3QUVBxnk7IV2PJubHshPfOW99R3WxKg6tDSFNrNm6wdjR0X
8M69U0/qdzN6E+fyM1HHOK44SAO+81aF2iFogjdYcLiG5cbnav07e38rZ5gcNDb0vpakRqZwtn0B
dS4alKRljA9+Medt/G3bZgMysNGzn8Xbpk9PvLrmaeP3HQpWJTbuVK5KwefSy1Yv0OCPKKECWQWv
t+P4mYdivGQbQqMy7IWPcioW5jiAtj1jXX+TCtoNXR0W6Ht5jCw65AzwbtNyJ2QCvP3JjwyReW87
xo9iXEVzF5pFa+FdqzvZ5W6wV3DE4az6R5moUYcZjIX8y5uxO1caRx/CrNbMblatO/DExvBLDwMR
aJuViaxCi1GX8uoENpD9qjyFHiSt2oauHFRFygo4lvsetl1qWLpFU7XttRhViLxeKScwDGoAsBao
y4FWx9VZjzpHepE+re3v2kyJPxRan3b0KxWmX1nSqso4CDbO0xtribsgVK1AWMcMVj5SWj4k+tNj
x2DZdRW6nHMEOdrClpmBkjxsalXRAfFfChTrTmbZWA+aaMxgUH5z8gNY5f/Cy9ebTney2VBdQ3fz
Af6QYK7Qh1Y0KUjZVw7m1IP+S3VBBb6qXD/9o70Xo6oLWY+et52+UEKh/44FnNMm2f/3QG2q0zTH
vYaY1nAhJs+vk0CX9Otes2/3ekqPireDZWBKvZbd8jo5ZIRDtyF51/t6/5KIP1H941fmos/80vwt
APJYAuyy8FU09tsz6Wc3hL9kbKAZFUKmE0S2IOCGYSvyj7TkXS4bYOHOyNyyYnn3KV3T1P1aVsB9
3TPZhUCAgpOEamiL8c6uMASlY3OvxGiaFgCjE7wklbeCsecspvRCXRfQ58SHGUQL//8cZ6jLCTuk
Uxq8p2Fs38DJYzefENlabHwNzef75w5/EoQrpXzm/9eAqaZNhwRUB89cGGsIeHFc9Vx7u5pAKfrL
Nw3H9fYQxJTxRaAyeygcceKvwFlfYlEe+f7AOlXdzPfztFeEdDoaCW2Z33iwhw+d0KeF4Y+ESWWc
HRHJPFSALIPMNd4mjEzFu+mawWMFOBU8r0BNAei0x2UthVMJrPjTwvYbselU6ngQJviLsb2pVoyr
Xioh1nsgHFBR3K6yk7M9LrrO/OPqvdQr8kRiZrX8YKJDsRr5AVU1x3b7k5FgWvEjGpFt2ik4S/4L
YfO+fb8ipgh1rP8picmfxuukSUIbsbHQNtY6V2Kv0/3XpDd7V6vH1R8Syb2f8y8v6xnlou+RS+cZ
wcl80tVny12GFdi+Ll+RdeuK9xQKCIFABpZILP4dlbEQGZfXgd1bmyDf1Hx02d8+R0v1WsAP6xn6
nJDJ2KSpK+xEdLQcra6MBamVPaRbhxWqXFb2mtiRkEtRlNk+lqW7PLLvMB6KNJKfGAaMjYyUwRoe
NwGB/yIrrZJuuOv7pvqjOOQEFCZ5KXtxOPJ+btVXkRu+n+n+Gg6QjCG9EfN0+MQimmu4Wg03GfNM
OW6yrO8/6k8Mu13aR1vJgLvgy92xGF9pD9xxSwxZlZH7QqFlulR3skMkwtg8lceeBLBjanS7jc5+
fjRqKkgrx3Khc4+yvhGHktcOdHfIc7Hnjv4EmiVHZxlY7utzXYQSfSEhWYw6RjcxnVi/nP4NAfDp
HT+MNBwRdF3d+6l/LbJWb1oO66eZ0973+mILDl/ipm9HCmn4zmD9cnacbAAovtgKCcrV1fjv5wA0
Vv2otOcEjYsnB7LYJTeQsSCX+k3x1ZwXiCcT5bOBYROCMNVXUXBGL9IHssksKpDtELyjGyEaHDS2
j4452dZvwQR3loaKk2KT9RJnWs3Fn+Pao7iQKGdn/t1FJ1V4jKKlaVaumZa+PfnukvW+v2buvgdv
9hOTZBAkK3Cu4OzoYc2sn86tTWE7ccP8cvqXgajRC+p46lqyqBaLSKCpaDOki2SCz4ezTLrgkNZ5
jMUm6QnX8FzAYqSo6pWfkagGNhpuolpLpzcPn+CqiL0OLo2N/zoimeUxuIIXC1udNk3ewi9YRKhE
1dXL3lSVBk3zV88VVWUoJMVXurKVRTYUxyFYPkabgX5RR4+G9eLDyXz3/+Nbsp6g/qWYBL1iFC+9
U2P++xqpwI8/QTDnV0FYj79Wav40u3eZ2CulAopheZxR5SbpxXjYZpAJZkZR0/kzQfvw9eK7ggBE
z2PBFhtOoad7T+oBi9QifcQHdqeZHZ5SbuBSb7PtPrHFQ9HJzhaYwXk8GivvptDtvKk5K9l7uOaS
2QrI1J6HtV838KcA15e6c0EWy6OuQWQWj9j7ndrcKfrixEmPWJsF6OMXyNBlRLraMgXXnJp8CgXg
JTKSJcCStNDSov4wEUfIj5+jTRQ+hXs0DB7tLbLibbk6XQnZMcPYRE8V3KPkeWnTLLaNNJcoON2I
y8cT+ubL6Ck+eY1S8atEN3jdlVsy+QHDZlBpZ1uGdaAydgfWOeUl9H2uy0rVII/+di9i9XaJBD5x
sndRMzydbWxrVYr9+QgZA1FOuAv+xrKNkVc7ZGEbkxQ7iXvqKm277Xv401N1epBg5u+ZRR04ERiM
SpcPdg1sRPWT4H7KsM2WHQvlD8zTccBGdRuWx+4S5+TBjEm/fH+jMmTgT/K5WajG2nmt9aCVcXnb
CX+LE0gf4/9VWSrmOqhykQF2nYcXIpl7TRlmPRTG3Qhh4IzcDqezURauHHQBp1iyhcL98OWPqH16
nHYw6sGOQsZG6SMEyrgk9aTKMv1F1EdIKQoGgvdFakHhnFUJFkoxeHDrloKY526ffZWZHpZFWNDo
EKb9tNjZON943hdOhRN0vqrgcxpL6sN3R02yZp3gbHrUTTj3PyoafC5rJ1IcICR3GP2/Q4L8inzt
DOJA6TPaaowVSUrZr50sH62SU8wRcYX/VsZrD7UxgnDpjXXdfHe6njcO2gTm70zEeX+atVSXqZ+v
pZeqC6bkH55gqixf0W95CJVrG4rig6U0AjsLjXpvHMIsUpdEtW+zOXk7zdk9khSiPbijZDnMZ+n3
XAKOgLFneNWSVnu9eX3S2M5XTa/dCd1p2PQ0fEUWUfTB+z/0BVrrM6AAQjwN2ZoF5AwmhIZyDV6Q
1hJciHrtuG3MsgEkepsf1h54SJhYQKxIhxfAhQqm+XgZjc5LZ7zKGai7W7hMqW3qWTnG7+qWNsOg
yKLk0WHigeCAI4FcWjpSD6ol9jLE5Yz9jsAsmMOFmeQdUSKBJNcIc7oiVdy7J+ueAArtzUW0eKLu
EwHVttI0Axf07H1LT7TAeeyUHch/r8elPpT7e4tear5KWDXqZD+XzzjKE95DDndxlUiIJYlJTDb+
bP3aQiOCYRIHLdsI6rLx4+P6+MUBTjrvGwuWqBiTDDMnZJPsCBW/f0Gv8BbBCNLYkwgMyHh0u9fi
ca5D2h63LwFWLvUN9vtkXiNr6EyvzZHMgA+6fEaL06XKiAeRdnsLywjxKEq9b0GYtUC8gFgnltQw
/k045jmNsLl7E4TYMDQ5QjYP7WsW1bIYQbWuMK5rs6ZaLBc3fTHcN1E6dDcsUBiKv9o4/oYDv5fo
7634WfYKztYT3I8Jxeo0/7bagPoN7KL6JABfbVjKSrPj/KtuQWhwQpjAvPF1mOrs2UZAl5LZL5MX
dSsXyKpO1XyKH/nb1fQG2g7zqchJ+pogb7P+LHLehmhSIGcO2n9igKhNYbh3ECCZriSUqfndCG7T
LGKZUtcVIj/J06zaPeGHc/9Iwt3/ArKS8nMcTKCNJ4PTMM2wM0fzAsnnzmMbrDxGZTDqCVZS66Gy
x9f0TMcUX0tGBplEtaedgo82En2dGBkTaG3C/INrfHXQfoEKz7ewEhnYpD+u1d+7csEWziQevptx
bc+O/y/hNvEvspeIc+NzMAWVL3paPSjjkNR/9AKuRpd5XSNpleFDxLyjP8k2Mhl5oIiDicvZl8Zs
+03I821P4DvbpTY2E5Fhw7akSW0e+mw3o82gP8ZnJ8+6QVFTQiBRnSA18ZlNkWYK84/jseIg3ybx
WkTwVorSFatu0Qf8o7+fXinO0VekqX+mffFsV91YYi8j/kKXXKsltEUflnKQCYwiTJia3Numv9ru
wle6sIF/TKQtKxdNNWBhzSoIii8pAM81Rn9I0T7GSEmlqT45RFpA4EP/HSOgj3QsghjzX78tl6O4
VdYMZTkF+8tYp/ru/7w8FBSvfkmLA1dy65yN91mb3wmXP1zc04e5/5qw8H0yxgeGYVVGijn5m2/X
O8WSYbr1AKDJnw38yUrLB1hTOZeI8gzMXCLX0Eo/MTEZar1FdO53CVTtF+kGKuS+IzYyJHP8Tbd7
nosHBe0i7I5ueOr5ttItNivXamIxpLweS8Sm/HGEQ0f+Pbt9IgW4JNgNM798DYVslSiYMihHNqs2
FtarwaqQK7JQxoHi36MMHiKtJ1OuTZwwgJrscYpyImUfKOW9ZwW6YZ0sjf2ZZVyUqyjvxPHuByjg
w5JC47+tvCGQkxsHTn038JNWdrJ5NfDwdkJn9I60cnqW9FZ6DjRSG7mSHUsEUt5hJDNNU/Hx3lF5
umRRlO32CVTtHDvwQB4SiKaeYcmwFoHwjkRfbFhBDgo9X6jlYsjPIwGJJKhtT1EE7Qmv2fbvzOvt
U1GsGd/vczeVy9+0wnDIRAu5EKqJDxqrnpDE74Qem9VC3FmZ9aTl7B2ljXue2K8D8nILrQzCyaLe
zw3M5qfaLCJTAR63rUS1zzBlDOhysc1eycDFZPyd6msmJfqkwz5u5rkgDUgp2LJaUO/f87yXzYFO
wXwhTuOX+8AAOthiYx7gRJFfbGI6sPR6UklLR6iMktCJx4yektwQQWVke3U+TdW/0obvQ4//Fbik
68Y9aGziHzFOISdDOy1Zx+sKQHIq1zE9l2Yc3+oaJ6XYDOauRaz8w6knYIDmAufH7+vpC7BmFDhq
usbsyx/218rYcPgFGVZKnREaVOWWDuui3/ppn8c1fjgsl9K+hor8AlOlqdKQTfax2gQHWdLQGPNY
V68kRdAEtFGK/C8XTI3nYKAlTWCbImE+RnUXOGmTSIooDxspRxXP9iV69qHwD1yyfeTdjdtrtxgA
QPQpDefwWTLz+1LpBtglhIfTd+oeOmUkkJAgBxVGV+s/4RlfIvhWoHJLe8sDhtB70W0aKghuILj+
iIMZQTG1pCHF4CZXTmlNaAtU+RgGuTkh9QUb0lU+XuBQzMyrh3bfCBHqeGoenUc27cDhBHq8L11D
10CNYOQZESUEXoGCn4dJjsjl1IDUX/ckK8LGRqzCFMzLKyvVDRSTKdPD8LYzY4iWxCVoLRiUBX/I
iLjO+w7dyq3lXswdAZ2VBS1JUjFGvufga/0FpDhom4zeVgSWvuileVg+tqobiZLSZhFS0pYQenpl
qrYhdTL8jVoQNq5FZ845javfB3JQqnDIzQDMohHX5f5Ej5EkYEENWPgoz74K/kxw6YUn1y7rwjaH
3jWqmosOrw/k3ml7xHzkBNM+RSLEqtScfbZa5k52OJLoH6Yy4pe8k2QcX4hoWcbPE9EkMeVsA1aO
MvbsREvy3x8upodmdyX9/sphAVIN33QmFdAA4PY53kyE6tfdnlZ4wenS4h0y6T5gWmTbhB16sU5h
yrsFFh4tNyy+9qR9ArhzPECJuMpZPaPbFFwqeJZGegMCEpKLiBrtSglPhuv8rxq/Leo8avK8yaxo
TxIADxVI54Rr3l6JVRhV9xt3vNej2eOVOUr9nMkVL43rNMnLUk19JIBJ2IMpkzQnc2AsDbSfjaNm
KTNCjdGqtFMCfqETaLJITYLwWwo1lqRON6aeHjcQ1H90CNLpV9Qt/JH1CR0z5TiK4+F9iZlu6tYH
VP1uX3Fv9iegMFVJuirdYa9TeqMHMWGixq7XbVeGMGJwo5YAC6zgjYgnheE8mt7Qr2sRUFzoKP8r
fk1MkJlrOKM0+SU0PEsZkunwo7mHW3N3RKlQplYDjZhgrFuYSXS51RlxEilApDaM1rSdBx2u2ZU+
heha4F/QV58Wm89ptAcR0+UaStWe5NaeopPSLmbCVPGGf+hgEJHHDcVY3CvuIBySvslie1ydxCwF
xt75pDwU0fC1GESSzf5KQrP1lDsYEMSB+ADCNCu57/RqcMYKXF4qgY42OVa0TvlBr5xc0/peHOtK
XegOm/mFIhu3ZmvpbMt6NrAun4HfII7KSfiRxEFDtD8+dbJUEFw+Yra/JMvKn5tYuNb8xKtsx+jR
LFf2N+y+jRO9Jd4mvI5xZ0TiUJ6gBC9aP+ghpdOvpz0y8xThmpMjeqr3UL+MuxG68H+Mt6duO2dq
yB1xLUItRVuX+2NCV0gbmc/o/JPCPgCL1hv4YRv0N5MIFw9DJIKelRlN/yznVEHHbErGGE2nvx7n
9/bRZt2eFiuqQmg3aLPDkZsgdMYMP5PXDFZvZ9cTlVur6gTuA3pJjzbh4naiVHk5MAda6RCaUePK
IzT/+rO9HkROP068titDSzAD/0FeQ0dgg22zjFjMQaPqflGTD4WxDwJG+NBQYW8Odq6laoKx8lt2
KJU2KO6YI8F1X5rgecINLAykNZflF6s366U2Q8B+EH4L7LzUXp9tveUN16QPEox5no8L17JtSfWX
7vpVkvqK+sOdrT5hf+Bs8PjxxFDVP6eROUuHHCwEruL+DQLf6T4wiNlYZPeq6oXuc91KaRq7DXFU
HcHG3YiEdGHTfzJfC3RECuCz4ENPuKN29QsyTSieB3rP7ejYxd7olCZdU0UUvbqy/KEAo6uw3Fzr
3Lgp7Q7yIaLnsk2jQ2OTlJEUMykWdxVxsZB26ksQ65YNGqtxFKO7Pdb+1p7V46nb7QH5+HWXFxEL
Xf6ZBoXaBmENBboRu5BmdeggxanPCHD3AQoH5zXpcRapZTlspGEfvjPHdTWkcyfOugOWc6d5McWg
vtfcj8i6vXYJWOmz9PNIEydkXIWYCLuXYxITStMTwT2z3vI9UF7v8fDZMd8YL8wAB4B84cLkexad
i6nokDW/QBu/Gz99MxPU0j0FcXQlmqtm4MgVyuSEK8vrJhgAjvyJ2kCrzduo3r04EOwKH8t1Z4cj
YtaVe7Pr/QwcirS9cSfrdfVA1bYreFuy8AQ9eFda00GRA2aSiojbGDE+all2wIXPfScIYxzDerRw
Jtq7j+NaNz0tKfUnbuQyKovxxPty4o5cZwRIEwmjVpA35QvmFdGeHCoPFqjAdtxHwviyuSxfwrVx
WkJ6bh/5ta8+090GZy9kWeN1Ay8ux2kL+73yPwDV0lW3yuH3tLKwANAegswXFORNKSKxbJFOyMII
ygouWNekETYE1Ug/FtdqK3qlyRPCio0XB92oMED8LE8lkD/AT57FIFQXK1cZeXY1KQ8Ed12Kwu3y
cGw2OLoqOq/BN2ElSW1W33f8Nxfhp22Vugbw+1vwjzs+f4CsXWeuOV1ADbSIra9B/SLm783aNG9H
fO6Ob34BB/tzKIpMib79YppNH1errKCzsUbldR8N14oIAWr5xqkHp2LAOC+6HTSfLrAIVADoo/Rq
VlgbdbFMz3LcBlhORHAjBqcrbV97ff1BZCroBPxWdxwZ2fbqXvjsNe6SMMYp8Ns2z2D8CuMbVqIl
+YwTueLbqZ/FbA+k16BtsP36RH48yIWVyw/bzgEvh8irNCxDtCylc7Jp16iLkCYMo98ZnGCCdoOU
ljvKw8coWXeoJUdwKzzR0Zzgr9kWKviLz+pw0uBqmXRMnOYASDpMJXZcyXMExsxacyDuzkPz7I8I
ftinushZOYqddzeOaYqJgDn0l3U88tZqRY9FCmMJaIIb2ywjzVlCp3/xhy+HENUjYZiDOLffkBT/
AkjsGxHRvkNucOTxUCCQQ/fPwOsP8XgRURIMj4d4u0ozxKED3Ah9YIJLynVQK0bzRty4inb5Led0
G+uyg8SF9c3kTgSajgNEtqfN+CmVXfrtEw7VeiTPHJpJs2Ahft17THKW8wk/F8xjGlWnmSgyG9H2
UcZ5uG7y4FMWXvcqVmaZ/mHSckLmj0Shimqjcwr6JmAQVx8xljt9U83C9WSWnmt8+2qt5efNNIXO
UsWv6NBzqHenLh3R7sCDMXkkeN0vX8UTICg/YPSlbG7yL/rbSAmmNYQimC7VYUBgb1LbI+eC92aP
tNZIuL06r138uKpC5MwpOOHXcwZONH65F5lW8TPxDcfwpD0g7Q1H4d22Q4exdLcFvwJ1l/dQtu8H
Ni9kxQn384JWgxxVfEhnN8b4TmTT0dTkNTbd8UF9GueI2G4GzXzAlacM0692A8JUXc/GFY95sf4q
5JU7z0atzZilIpJhMFeM5kB5MfjfeTI1x7Qw/3A48efwALfM2avS9NGUQus0S7YZSp1DG5AnvZAs
2kW0Wtly8gWvDtQBxGIaURdLAq8bUAVg2rAtLQXpSWHwjte4Z+XBSJeB+Glo0vdiojzHFWj1s8UV
xYH8mlubP8OfohQqW0FHDOHVaMbgptwnM91UFSeVdDrbBuhE5KXQrdWoYLnila8k/49/AENe/cU+
6xC7OfVPGRws/VicTf3TV4mP9buz12gMFCkuWV9wYGceeBe5FPFVE3uYGNr3AB+PtVsmM5en2Y3Y
D1Y1jFK0yTHzR85MYp7ELDnt8Vo8jo9ttKzUMLLwNxiRN5cOoEzaREwbp+x2rZmzcrtEtp8bth83
x+bGGrmRSUDFGcsJ/e/Wp/Jfhmrnwq8aj5PO62++2lfrYGrZUHx1owoso6lWe41aBRbpUifgdctS
E/NegDLr86Nef/LeU+uytpKAD61JVcmTfb6MNPgFxpIHmyBQTY4X2wjS8fdkydBtvj01vXZ2NzLr
5NgS0rVcJJlaVlC2DEhUJ/CMb04EkKUgXpcwz24fV9+PAB/ilw4EEKqOLoCbLiXOCp8n8keGMP2j
QsksryJ3clmJIkpjC1SRvuHpWmfAFfILEKFAhsjddIdgymWWb1miZzl21ixku58PtFoNLIZz01fX
hjjNaFp0GTyEINn8840a70PEfJo63+xoRN3BWi7stNBSa54LVocS1pi2KK8MhEwjZlsaZyE98rnb
S8aaQgsN2aN9U6z6Hzi5GvpqJ+Qw2IN/HAkW9c9g8z21firG11NxGr/uFIvYBsd6kM41bRo4mexy
WeAmgA6HP2dcy2m/wzX7J1xWPLXNGWEA/kpWayfMD0y/XEa7OPNmYKCSQP/pncTbPTFBDO3ACu1k
JF0vvZ8EHrkLKNmLStXp+ooromDKhDwTjlrKO+z4LWx5f2Y0WS7oK94WRzpr8Vw/u49glJ0qRhdQ
51CrJ7y74a/EApwufKvKyEvFC5HqbjxWmkySsPZx2ah2Y+CrGF4Bo5lmaoR5+oQPAKcPFeqUhIxT
ereY+MaakOuL0YzGrC2uaeiNHx60XZQ+8m4eR1U1NHvoXdlxswVrBknscUXBJDzQHKTUert1cMsF
bYrm0CyORwx0Fn3/CO4J+UfqvB2TQpvNx3MWmmAcL1AogdnDoDcEQgR6rTlwgdvquN35DyvrfJVF
QUdeLZ/Fe+D0SxuY3SiZ05YeJ408HKEnap4aEbwUWfu4aXKVL0QzCb9+B9SINLbB0bdMV3hAQTSO
mOrBG4f0/VnidiQy8zc48hnCYZ4WTDc4v7g62y+riv82wZx3k4pZ7LgLJa7kiIh7Uw7nRz4yK7uP
zRdSlK94tJqE7rJ+oXeRPqLrUU2d4a+64HWcBqcaWng2espBckalxS5ZpYb1CM4Dzgf1ZHOkYVSY
eQ+09ZwMaoJqILS8Vb3kmHzdvdE4SS1CMFDNM4ZscBHjPMmyqcyMrn0dsXDxC+df69aGoSP/yMWq
C5/2AOr1huePn2wnObBLFA8dWNmES7FLpjJAwTcgMmD/IjaDuZ27fjYp2XkGBpjWKQyhlN7Z/rJd
+AL/bqftCpLTJRAZ8szWKDg8z5eKafp2z7+4Dh7088rkbCWVx3pj1voS1n7CiWvCTPz/HnnOGyoR
/a54VOhtk2m05hKuMF+YcghzYKGSYYyZmXbmI1i56RehcoEI552YC1eUZjwuT5xapBP2nTR/cBaG
r90IQjTkHPkWtPTCyNCZSe7+VYGi+q2NhKar4kl1Ojun6omv4R28GrdF+egq+8eIV5wmplzBBA07
CTMCZps6R88xMHp8eqYNK0wj6daohcH/fB7akTMpuRjNbZPIyruu0B1CGfeVkk9f8lqMaoEYQGdE
Vo4YcMAaa98dPfKM/Jm5Ccra4lMxfAlOo9DpSTj//VVPqM06pCez47KYz+v5s4tmBcaDP788kIgS
Qz/1YaU7a9qZ6Y8RFkKBHk8CDJRMwoV6VXtt4tNeJY4DjYGib7FXtVEmQS8tp7vf4Jwc4oiGjZ3k
ZqExBQKs4Ay8qvxgx4Yogw7XfaSG0cI4fxowdvcNWVj04vDJvMdF965Y6Bu23tGiT2kQK9i5UIyV
CoM+sokehoV0pd2eCLZEsl6Tm1Bg5iIOaTszsieAFCJUPCbUvB3Sz5pC4gydTfOYwFoErZKkC69w
YWLRfQ1qYfp5/uiCH6w+rgdhHD2j45S2noarCkdgQtGldNoqWSSpmHPRt3yTo+Smx+KIH0o4q5Fk
6GhcXeCa7z/OPcFdBrNU7sTwhRQ8k7J6VwAHaDLSGv9ZcDpzPAxLzQ+6DXauJ085m5gsM4kQ/+wQ
Bugy4HMiBTFXXQpEKJUctS5lkdlYXdCqKwH+OCD5ua7Ow4zX47r2MH/ARetktq9DZNKYvcyLnp99
cOR4tJdWEOsUtvi6EVDyaJZ0QjJEkoXK5xlYJMqyFN7hYWK4oh4PKcUQNPbJgwUB9I/HJzmnvM/A
zFm2z1+70xm1BLS8fg4pk+i7D8ptqbQ1r0CeH643xXVVL1adohkuyVWgEz5Dy497cCBBcCCofsfx
12bIx7xJQyVqX0cJkrYSxanKlYp6+L5JnL2rZbJAVw0Xn9Xx6hBW5Fyg4Plzy7fXeeojrtVIN9tR
awKd6m4XknSrrAEHiiK1F/oExGvBoCFgI9ClnknTk+uP0CGFH/oPS1HD2kQOm/morCMSqc4ZxqPz
xwSNQ1qRoPcqFD/miAvwJwoLz6ZNsFSogvsSj/zHKef3zCj+WemHxx3Q53NjbCwyWsBXJT99EGaR
oqgOf1ZuP8m3bEaSCzVwFyLcL2rB5zVFOWEQPodzEoMDyp1CooIShoNSrHWsViFhbtdLQtmMmW3v
z7B34mvwbeZzVM3yYDB2FukSb6BYu56su77mBvC94ULFiJRx5dlyB+owu9VtzriCdylR3KssNuuD
nFPV4Vtjdql6tThZN1/I6wyY1pl905FWLpP6oOkRajHCekD42FpwGK5mrX7BpOwdzG2e4YMhlSN7
3D+BpMNUML+Un6RBwg5D6u1wz+m09YQ8zsQGJyuqImsQhraPEBCR4GJbNieRnWfRrzXMTGL65rgV
deIK1mQk7LmfV0/DIqjOlzHfGT4hnMFf7uKcYqjf8TftThxcLv2erfsDo5ZtoBrcGrlJ00OW9aic
ZH7lcLd2ilbGTQu+AiJ71mkdkMEGCAQObxGe9yR/98G7LKjI37qBzHj6kyswLH9lEZHgihnpqrmm
Bs0L0tbPXeDyBa5rCGECZuWOhfQjDo3R92Anl+4f7b/HVvxpaQ7vK45H/qDBMG+Lw4TGRpUmi0Vx
dWQdzGPAucrW6JGZ29y4mCOw7zMM/ZZMY+v1pGxoSH18cPF0YAt2ppUibGpvg+JpESYrM6AXYo14
zf1kZdV0OikYArJ8tcuhFVged6ZPSsHFwcLY7GdIFrdvLCcxnfyiHU0oXIbJnYyT2sqJK372e3/+
74Zi4Zv11mn8xIgXpziMALqrMUQLd7j5CTr0ZOUqXsT/P+nEBS3UM+YJT+dX+ZGPh0BQMYrtTn7e
uZE1CES+ScmnHy88mbUHCE3wZ4W3OBnEF2quFfQYTjztw7nLI9uE+ploblxHwX4BuJ+7PYM0OwP2
lqVGHuMeMVmFoeqTTiRvKxMDt+PUYUPaUwuIxSAL+wOxU0DxenQNeMrTJDVepeeF3bh9q8EvNIDK
VbOp81e9WwTskyTCo4+fNMCoR7AmSYmi/8Huiefc/jKEebXwmRr8lm/a+lqnHHli/BXLrsl1FC1c
1t1PQK7KJQd9iFgymZ/IK9dvhItyfcCVM5rfr+/ddqC84Wtn8AfioeuQKZBcbDhx1vY3ixoPX08n
NjiPNgbZdOWvDdviaZzxMn9YmAZyRHtRu/FE4FLmwjCOvau3jdXXpvKp2KeDQ1GXXB0Kky/nr9Eh
arV8UWnHUKbRxRD9pYnBAMFIMHXER0070WqlVMCZDwpJ6l1zdktXF4mTcPNNjVHgBrkOLxc/6t+s
GxfohMmQZ+3PGCUZq36Fy0gw9XdTo6X2zs/q1LIOaqZI2n2kc4zUm5oHeddq6S/irnE7TUUAnJM2
gPfQw/4Ckh0JqwydAtVaCK70uydPeXOvZJjDTGfM9vla1Pg2WNlWr+qPA2ih4nAMLz2EemIyvqql
xeCBTxgbNYYN1zlPmG+t2S7fhf32HHNdGVXPxF4HqbQZwwm3pbBhqc1wbsw+odQl3fErFS9kfS+j
PF0JMfQOrBmbh9/nQvLgvGOBsejQg/Z/ztT5HG3JEkc4Hp6zGnam2WjZ7X1gagLGgnsjBriKO9gz
073UXBfyZINlSat4EXFrA0wnN+zHTEW2wblaK9h1W5soIwJJeNHQ963K0KVkiAJA8VqvQh2ulBfa
qsPgKUYNURlxHwGUIbw+sRGd9ajQpfu5UIhAk87Akbz3pnd5w4USLjQcyQUL1VjObyfAjz4Firdn
l9sfCAKz8QAOiKems0dgtWKsUmuo1iidD/iN3BPU8xE8cKNeDIBdN61LauyRuJdzLy5pvPOxVlgg
xaWojii6Kj9163s6MfxRvlUtV2LuHcqcTPniFnKkK9fidVAytNIrY8VU5L6/MUUJxlJ2vTvMred7
5I9P5IFzIHWCertcT0Tzm9pjTRbnC6w/KCQG8Bz9bJxiJB5k79AKEkEdpq4cT0O5LJTjTDO6bksk
4QgpgtDz6g/Po6Bz4G//TKsHLQIZeLM95gqgPiIvkwZx2SQulINdX14B5ZmwVITeL8b8n0Dn44UI
WE17Bd/0p6e//YxRJ1lK7Ms8l3YQ2XdQ1+IPBKug5C8JJeVN+qHJJ5BFORpw1x8y9EapG62192x0
4m6g5ygzOCw14rXaJrlApe+7wSYDBXzNPCwtrclI1wJETZV5FuMkk7StoYke8cXoc6mfUDs8XFbm
Uswjs/GelvZI4aMkAgytZ4fyNm4oxGc/u1Ktklb3WlzzndQe7P9p1u0aenU6mATV8Jq2K8blV1qm
E3HLOdhoYd3Rrt/RgVe4jYwgYbRe682VfiyUKgaf1gOC0dBt/vjVElWN6NW03MU48ORfUz3iw6hq
hFr0iuGquYct0c7u6FlwXDTBbNzxx8JW8tyYlMOejATzm4C9i2rjc1634rBk/bIaVnQRtv9Wo4KU
knD49u34SWjEFBIbcrCcrVQZF785ITVPwegm175i6lw3wUTT26qdRaahR9+UnV2A69B9aRsjSYGR
FBdGICx78gA8B/R2LqEZcxxaRV7AVVKS7zF1Jpt3eLwarlbJhQ9hCQ3A5hwE7TS6aeST0ECMUS87
CAiNxIQ7Skm+dQSRmi+YhoR3DWk7iyaX05nwKvUxEWuWknu2HBCef2G2AXVk5S5cMLmdTMmgeA85
pAyjYkmGOuNThPWExNeSyFY6TgbOzXyjzhFsqfyniSSbJG153SuGy+798zJ3B0+asBry2tP1NA0n
ZRldc59J/y9r0DCtnZ/pF3uztXYX6LWPcfv8M1oEtIjF++wTwHbJ6sDoMLyVsKOD1QxIXKrsYMCD
GZghnd4w9IpiQWAjbUyJk6v5XEyCzIZo7OfTfWdA4lKbk/Ac0Tl50tGKd0zAzFIUpi9gF31ye95y
L/F8O8fOm9vZQmLjPuanX+d+Drg5M4mjzcTTRWwYNNsZL6eE7Vt7tXt3mZqjfXVUbWtlvsKUpfYP
xZdr/kwvbpzj4x1kbP4OYfBCj/kX1HaQVuKJ07QShjFFVeIbrTE/zTaS08nGgAlwo2sTs7y2bh84
tYRaoX8IsbDrD1OEHuTe7QVMJpwDQ2Qqt0/bPKcoF9vFhtkWSkWReFogXtHkmMS4aAT1E1SXn5cB
6duTPc5acHiaApszHx6jDt+yb2ZaiLKllWwrHxYe6hmcMfQefIXceIzoEVyBjROC3KNIIscAM9hM
99vaOTBBTBCX1m5g5LbsHDupRt5n87SejAKFCw6ESJOZ8P6H/40nT5ZGnsGc6MST4zYU9iTN5abP
4TCIZRVGTkViBynQWiqcVdi6PdvE5xrUq3R4NTmz8aJ7+DU2Nsv81/82ba5K9aaZN67DhMRh3/7m
/jwRaz0HfJlCGopCtjpp1yog2qObTBLlRRfuPMLgWMyWGQJl6cV5pkQfMaFExhy1ha5rp4CiO6IF
WbrzBvfzN2dMq74gqOynB9G54PpbZZSyZ1odXke7OOhQllNfa9SxwdJMDDGsVzrxpwacEmWZL23Y
KjvidfYmgQ4MOlQMdUwhFqCwh2ULyJAP6mgLA3JVceCqidBOTbPPAmtIAeBoYGCaK0h2D0EmHtSD
bHyi8KEl8B6pQUG6a/86qvl816FK9v2ha7LPK5aQ+52rwRYFixRmK24ikeqqjtp6zlBiWr45mTfM
TRPq1ayOe4cYEYFB3Nfkogtxko5LabjoQgj0vWibWUjFTCmS0TK/b2JctFRHdqRgKDeNzAu8PIcx
sLBUrmZUbHJyqKEsgFWg/DjoMrbN+a0CvidCmtrEC4vZPRmMjr0lORFyZPS4ygZxufj5a5iGbVZR
U777xVNoByKbN5puOd3JW22Cpkf5Z/6IM2gRz/NXzkcam6tnfKt3451kQxIzOE6pRGvaccpi9Bz8
l/ABZyiIz9oPsxfHASvOCpiHiZddaZaS4DrgZLubdGo5SlFSeF20vNhbztdBBt7zPEhWMu5xzjYg
bfpZWm9xTIkqFPH/CM0cMeHdU+7IwRK/xQuR/3UF+6hnbrqsI8DWIVOuzj3G9EaM0CYHBI3hASTW
cmmg6IhJJPF9LudwpAtiP1BsWjBZslyKncpubo+a64KaSbPvucBVcS4AFbvrhQe1bdY4qdhkcMfF
4zh4Wyex2FV7mJqL/Hmmo72MV8vl/P5ORV/oxPLyYavmhjiQeEgh6e+j17yEOIf4VLiTOxIQ2Xph
ogke3h8zXsm1jX/ciK0kgvW1Dq0xOlLqNZm7Gxm55Y59OWjOXBDVrF7TADaXtRVJMhsOmwPYk7tP
hxPWDH5Ut4ZTNNy6jdfGmVjwcuUZyB2HHaSj8wtGgeYgZq9waa5G8DW/LL2JCY5LLOgUW2DKG7Py
W1mcCE0tT3j+59Miz+A/TVNY4YHRz2L4TwXiZ0s93l7fr83zw+iie2hmz9a8ddO0ePzIVthdt4/M
qRlXCxQ/eZziwRcuTgcNcjiODqOMj+c3MttLev3CrCVpPkpMUZ6Wn4ohVcNh4YKna8Wu+CxQdlBp
nQCM50BxajU7oy6W+WUvKs8GwcrmNk4xMX/yqdVmZon6Pe0F9FcgtThFDNcMaD8NBDZTJnc7UGbW
JiXsUmGj/op8Ns5Amd643jjxEP9Cvh8ObVE97U8xqwYZW9dWBaAONnjDbMd9aqfFcsqnJxu8wvvB
yn+5MMG7zOuJyjcUsaVlG1qfY8OJtJ8CiD6ekjl7XZNu9Vbg0w+v69iV9HZarizck1VLY0zbcvTF
zY1MKmUiLnFo5+ESGqUF3zerMUcNmGjVFk4K7IT/fX7HV2QnAXPNS2GrFF8d96o6HVu7eUF9+vzW
sY+MaJbWClbaN3AOksMdKigfXYVP/QZ6cEUHahymXPcXqHZ+ggVT7xSWjDJbK+BMAEK4Tms4q9Dm
Kg9xZu0qdUheTN1WvG5cTt6oQkdOkh2MEhBGu1dCTjF0XKdRMIauTBPDsDcHEeyz3vlZMezUm7Ns
cw5CP6+Ywjz19D7vQKWor4TDdeBREdzDl5El+LWh6oaKcb2bS6E79io+j/+ni5d/ATouUMHTfuff
zqA875YWwljy1vRV7lhzbEjRsQex5oFMVZKp0DgctO+sape95LD9UWdIV7UOq0OT16NS6GqSMoCi
inOMjM/pwAhfatnbtpvoAxy7utlKKdFhcgvTAUWBcXLjLZTmt94DDgoemNwX8dhMnDCViJ+X4IHT
uAQwmSt4/OTqCqUxJNmWvfYFM+RFGH+SC1/e6yZUImG9pe2F1JIQnKncjIWWKCzOuutkF8XyHWnt
0LvgcTkUaFtkPCm84CU7rCZEeT3xHZM0Qtd5GuxyGQ8Uaw3ScMQg0T097M7Ma/7DOYIDausHChRi
gvlRjFbx55Dkk1QfCqpQvVK5JwAutQfc9N0rucCms39os/Rx2hHZONpnXBuZBbD19iA6HNch5/wB
JX3PrkeO6VfxKQZ38Gp/4jmvmvyqKZEAUI96YtaIr8JvB15a831hfzMaNQIo/1vjFH2wHaeyjGwu
iWVr/wDwZD1TUH+kwFVfJ3p45co5u1kD3BazXeBRZGsWDrdSYnM/xHttzvWPXKhtNSm2LHt00+Vs
drhpTC3VtO19lhhXcL0n2zmBwXZ35J6p3RoCkYjGjmASgk43hGthcu2HP9CXleqVlRcB3ldhzNKa
5rzXEivG979/XEI9M7wJzVTvP7WDpZRaG9FxMtVOVvCufMonqAKqMcqcUn56svtFxWtO8C54DPvx
NQLcqM1LWPHqUZmooNe/HM+0HvsrpQYJAdHcLiyYed7+4OKaCmsvkpJJfogYwaGn336M1b2dcgd0
U5QSmiA745nSib80jYvkGzZOf3doWFABxRtaY97Jb2xlWahBnkVUnFphtH67m7/zkAbqwVQQ67zB
whsyXZyoCt6MfwFxfPsGir4AFqA31DOGguwm5NNiPRPLFVTMGbiZ4qwX4mBOZrm815uFb1NjWWwg
8FO+Myvka7gIBWEwfkPAWgR0ERU/b6IHWKkP5AqFYj55GHlWFnZoVoRfjdK10vU9wsfIwHB2Iij6
mVqBRNP3vMro11sx5llfjunFqdO/1f6lekG36ckdUtHmcNj+JRk6M33XnUe0KEOmGfTQroIr0KmB
YMzRtVQMMrXdKuKyAQJHtBwNrg9Ej8+O51exFpriIBQul8app/DY2CiDRBPJGUiGv+o3mfKRaGbD
e/z5XG0lcRTeL743EuD03KWUdfuB0q4vx2Nj8vYGvz5y7PRABeLNilwGdsZWGlyhCxbMsfQnYTHq
Zo4p+YE+AQiByws9IYF7pp+/F0QMPqAsopbUpU7zpg24kzsJOP+bM9liBuYOXMQDr3MqKHvvYeqo
lquTJnQeSKc+8jmHwBdJnWuBD4T0GxyK+00wgd5L4x1PcpOQPyeJ9QCWnTEY4QzgT21kcUn615X5
fFRZji09h8Vn7IiKrB0jf7+sp3G3xx5mK5XoRMUs3SOKSsWrbV/fHHytgJpRXtvH7gkxGoqu8ruu
AoISQeMT7LizIKFv8D/QC1jX0qavnL1ZMSOAAehYQ2qViQ/EFAD8L/WZy47cJwH9VYQloZrzPp61
dHxrzv6xvQbyJGCmCL9NIRFzevVhajQgBpuYsmJLZKzU2TSy3jmwOwNsWKzvp1dDMRtsev1OOyEz
OgFnKQ6HfCGmk0zKF6LJvEoKwXj3tefKGPuFFt8L+rJRdMwMLNaEmvIDvKuhQ1JtIDKvCUf8I2yF
hr/Vc2GxXB9LKDZ4H4gIebzDpN+ciAhgh6UkZL35zOqlOIBUjnyYNPsjnNQIgod9F4QHnffDKyoG
M+D/BA4D7oqOlZOxva6RKI1jigYh2qw0O+wgyMEUy2RcTXkfX0S6DdQtBKAhH72PkDJY7h3GBPEs
dvQqi8VRDSlCf76xQp/u8cW1Rq5WcEGP5SxtR26r5xzMGUiuwU5TEJ6AP2YCVuMuKuy2JPrkW+MV
gOKmqY3SyAXp7Hjye+J/YL3zUx3eTMOHstVLDJhcMROMgfdf/dSBCOMPiWNNoEmHjd0vAAAeHj3z
zbStyyHoQwdgpWeI/T4C+tJ5FggCE8/K6l809scLZtBlkLdtqauVJM4pK9dwOv+FTJXlna3zxewg
ngcUV2CiSx1+ySJYZzMhezF39v/XX6CCooP3G94s32tMOvj3E9itwTXE4KWgDIxUmNusVvC7Tege
bunmmSe/vQL7c5IDqmxmdcAiEV4FAbxjtpwi72F1O86Sd0FlsWgwM4TPLDZ7MJlHZS9xahaE7+99
lxMtZc/dz8JOI3hL7ksE9kkhZ2umpJ/JrpF/eZCnbETcoqtzVm1j7iuQwrBP0/G7BMMXfQgq9f/3
pr3ms/BcIbfr/atr/OIJhnf+kZwmsM/IsbZu7BmskxqBdj3GyusalMmafk7P8MvUFdGiuoI2/koG
67TZ2p1ZRj+YW5YNCZp+MKWQ40iadBPVjM7Ca2H7AWiwCg4bA5/9iOwHCqzAbr4kd9jcLO3jrLEX
7m/HFPDOlewMNhVrAzZaUoufDsS1IMg/JHqNEEjV4SHgsenx5AayfGGEokhtNuWQIEGrRzogl31/
Pqjs9QRPok5Hjg9B4O2n+S6dfDtWQVTOLKEhMLHHHRatPzI1E5jfz+q7abtseIaA0BEZCGIu3SxW
YF2UXo2nJfhtUAMbaCLjkwPwOFch0023gzXg33bVc8IH/3YT0VRpWdif8J1eBaRwfMclYDf+n5CB
OP67mbW2Hwb4UzYwrhfABay01putY4VplVO0I0himZBV1z1hTIC20nZGhXRgR89ftHqL7vkdlN4G
oc9bzMKfwt3g00r16gfEzxYYRwXd5h6FpWsOQkJlJ1sFBmHJRteuh6i3VXxbdpOitas87JNcLRFe
zgFbbioy5AK7gqhTXjY+RmQZ0PaMJDjw/oDOZ8U0dv6hMzQKhBNIX9J+mBjjxLh5b5Nne0bxu61l
PgOKvl2k5E+bY1VHliyp53OA8XTCHT0AfnleWivKDtkJ0WiwCh0OiQPAtwy9hC4+mfen7IY6TGQX
7Z/8kf0qRir3LLez0Z0pNjymtJetEmcPoRQJ8ZrZjqrqaOsICs6elZARVQhMYDS2HYudUhTxu6q5
0gZWRN4Of9iBZzULNoFdJbJRuzY8vSx4yEJLGXeS0tm/yUBumJSBip7Y1dqYUPTH1MxrZ+2/+8nP
BMRsBmOv+PntNVIwDGpWpkSvgyJkizNEPXNA1X0euqPu2dkxEu2XXNs3rIjgbp3P7ZVlkPHuAQQj
lEwZkq+C4woSZNQyjqSFAR80gP6ahoOew825q6C2pOhbSYc9M2SGlsjN7L0YksxcOk9hQY+4WpJN
eTjWwRLsGkxE9npGi7NebZu7tlYEAl++1Fjl7M54T2bYbkxXIMDsAwO7vQYqhu7A8i5kkUJdJHva
laNrMXeCFt0FZedNTTq4at82hN4P4cQQULlDar4lVCdSfBqG0DeWuBcMl3T42rTgWlnwve085WvB
JWLuYEO63s6Y2xLQagPtr3m8mglL4t87TrrGpl6WAekhFVWpg2AjayC8lQn0/2fL/LQscBXEpqt0
tdj0nhrS1tIi0pZk9p6JZRzorGZReAuZszALfpo4h+JnZMqC7+dmw3mZNM4iauaBy5ISPqgBRmu+
SNNEomQF8tvdkR5Ztm7j4u2DvGPux/+193hepg4yWKr3hq8g/lMCkfJmiJKZ8tQMcdv3djJzuh/O
sycvtdgJvVCRoeUnr99/tOErsz48kvs/+lf2ItlH5XEo2gCOVwnEy8jG+HQe8ZgP7IUmPuKHAy8b
BuJmQrzbg8CUDNfY/NQof3cY+DqLBY/YvB8tm/ZdzP6eeAIqrhpUiT05Cz/7eeDLxS9slETXudAF
VmSsy9MElk49Zq731OU4uepBkPUG1NchYD+oWCZ2qxQYCDlM9tffK2ZHSLXLHCNTAt14QpjgvBLv
mTe1I3GjyAKkidOv60MuNGEw5PCf2qdsrOFgOQ82NY62KIjqgOKDRo4wXlO+fMBSp7uI+j4AP/eE
awfWOtim868yOu055OGtJU4APvChqlbpDmBwoL8Gu1Ppqy+won9oH/lLqqHyZJU8eWsgFt4yKHkQ
JxeNScMP0qiYbggv+p0cMOZoC2qTM5cEfR0r3mN/EekFiBQNilUfohXIYAHkGvqtTf8GhuJC1u7Z
I2Mdqq+XvhLWwfVT3lNpbf7k0Efq9hGxexQP4DWG6SCXzx5a7jbeCztXaFxG0QfU+WuWu9xuWDDp
fGAsyAeIq53NoE/WRBY5WMhCFC4qlaC4LQiGwjMLvbJsVfk+ER8MS2gKdXNKLM/zi/4jf/X8Rj3r
ydwH0gBUuCW8EulbnBDVX7GnmbXeLv8Z9IVMqUqXs79g09txjAu3A3zwR+ZNY/VujkzPvbMPmYSj
2b3QtP/oqumbfsQBfxApaJUl7YDa3vh3RO8Sry8A/uPeJLMRmt5e8IkF25iHbRqk3JVsUqH723Ei
7cpeN6Zaj92nRQdFN+z3K8dpDEKlAOVHkZ8rxWasHZTlHBn40zmHhiyOnZlIQdDdlf9LvLqCVmBx
mfdse7R6vo3F4gFV/FhyM7l6yIS0cr9aazQcLPGlCFPrWsb2yGUjJZ93EtnY4xlbMhWuzIckCkxq
uY2ecUDsRh01QmJ59xcurCNAXsvUVBg3Lxg8xtfBfUViTXlGtVpk9El5M2KboRZ4+vp+H/hWH4Qy
UetR94Kmb8FdnJaHHoeBOH7LZdXdTfpn3t/bUztcDbXZuQx61ija5ans1ukTcESZw5Qc/OQA/swg
DsdIP73eAyi+ASHe6uaD8bhpvB1WelCOH9Wo6BlzrDgsen+JqY2xhiNGmCnRzUhouyiYjrqjQqeA
2c26SVVrqR8lH4ppw7KYSNtTXnrNVJ+PaZGUCtQr5CyRqB/er2/yVzwFYvKDKYVzJnXXB6PZREJF
+AMZv+ZkCjrV00AGxWV/VAEla49vtfCutLl5rQEcmZFrqilW+pgRZo2L13AfasLDWBqTODVkFgTO
fCkFn/q0k4lrNZEg1HV/hOhGAo+qO5Ch+IGFNUrBXGL1FugTtO2KW2aft2V1XNLpM+wgnkQq7v1J
vK8/wW5hM7xgBXw6MjQmtKR1is6JMTnr9ybvJvWXwi3gtS5Edp5yEn7hRycE6geuA73fFp7xhkbJ
7Ew8rKO3jRcoill8+746nJfY/l+jxQsbRJd8UmsEzEqrn4rQ9lynSHqU6AtnPUBsyeD2EohfWdP5
MxVPSJOUoqUs03WrBDkn+coKlG0Uk59zRjILvL6jvChAHrlpRmvl1XQ55KdTdJfQhlJw2y0Sl+O5
FPffDmE1+gxiydU2FeI/DShdPyuYBCIOjZNHibG3LIlhZbnkQVbFBamnBdGS142VtbKt/3o4xxHe
GL6LeDxciqNztht4nbFN+ntmIBjI/34ILDD8GFxEY9jAni0r6qxYhZvWBlJOf1AR/t05XdXxaiS7
AK/BHKXXzd+ZFtMQkqFLOVFNplndwvxwE+4U2mcuYXw9RIwAAGe5x/nS30TpA7XmbFKf7T83e3ln
YnF51zl8lHvfzzBpnvbLuf28My2iyptfb4t+M0byC2Nr3afYrPaKUkvZ/Vsn42ob+udma0WtKZcV
rqjRtmP9JCd5LKHcMBHWG7lpVOZyELHpq/SBx7WPoHg1WtpZoD0eUlRKL0+wotP4JeHTHs6K69bH
2IAxCZXISAnO/36W5CVQxDa+GwNql/Woo8vyucYaW0z9ZyEmH34LY5NKViNE7zUNkzAbeaPI9Lvw
TGgR+USrJS6kaMPxdK8KOkPkCPfsWnCE0RaKOdUDte8cKo97N67KTpuHJvIJl01DsWaQXC5A9ogD
SlqmK2W49JNgOC5EBL52ikrEGbOARglzJIO1Q8kaxpQGmE99F//9RFzyHQWWsmHeyNrsip4HZLHi
kycDokAerFDh0xz3JtcrzNuHVg9/27cQkSHM1SKM8B+cXLrV7aUkVjyEoXewEv6jrpWNorGD5ioI
fN/kNtAFCuJ7fEE9rQWIiRcPJFk9fwkp3ec87TPDtjqVd5nRN84Ir69HHuzZaYqmO4hxSnnpkAoC
pYYsKFFN0mU46tAw4dO6+AELkaeweVYUzsha0ff1IezrxPK/zmFkKvh047+wmSRBFLkH8w91j2SN
wEEgSZvBvu8MNREBznXO3lgpWPliQpC0+HH2est/s9byZfPqSP1+bPaW0CTIlcR/QGWysTcOBHNb
y9yXsFgE3LFrUmWHUGNZNRVmTrVxli5P44ABqRRCtc5YOZiFyWa7goMc5lIzxybTyizi3bOvLHPt
cKLEwkbjMMQxpu2CYE/AfZLBgUUsIOfAvoAJbDtwTHOVBoeiEV47RJU72U4rbYLmiKQRSIoEJBV4
pCxLCIA6P92OoWpgckCF9c0DXfcFChyESnj6Il0xiVIAuLQzwG9grIXAdtN/pCuR+0DTpAu2JAIF
XSbWOp29uzbt/4qrJnGo7v60Wnv+eK8K0BQjWT1ppL0aLf1tMfl73nxsjdXo0uwEAodnDuMW4yow
GaIywHRHc39KVRmrfii14C771ExCWNMSrctEQ38nyHkodYVB+jOduIYQP2qeu1QzXZDJiBuaJVmK
rK1NruWlurUQ3YV6mDanZnx5fFDE6Irz2OlCOA18cGUqJJ4NcNx2vKJ7JJqf/G4dX8ZZ/kIvlzUI
QY98olgBB3JZblQCguJd3SW8Wt7TR41FCSJVK+2ZBbzMHWdNMQ8BN5ra30PWteeEjr3EBF77wpmN
RgJxKEFrsfhd0q5CnYf3PVFSII2VR+NNxguhZUNc9IUNF5k5En++81ZGbPoYasQjzPf3DsQAfmJg
qEfPWEK6jxjhiElT3bx9biRcCBWNnTCJDjV39UzpRWFofPtWr8rZ9nJ5sc+RtBGstke3A94iukgT
VYcbKncIxEzO/QnsUxzY9VW3cZ2Bq5VNzSkZICijP/w6IhUeqRRxkL4Pp6QlXzsCClWWswgmXcQA
f4NIBtDZ2zrABIAZWNwm09o7KGKnMfMIuVeUVAig/pA6vzj3so37uzQtthuZdjismgrKNtYeXAsG
1W6xjo+orGNiYDJnJPAnl8KJotKk0tTuvQkDZ0e3n3nhDHEw24A+iUesV9yCytvj2a2EAr6M9GsI
xDUs2Lz59YS1sUveuoTWh2CzpQCzGnw9OxRqhvGt6maPKD4vuYZemxcYIB+bzVuVjGCsANy1trWR
UzyQj5Ps1hpLsMcxFXSjnyETwIYqRXgzesl9gM3LpfwGRdzk1ss8Gg2+xNh1nUa4/X4uVZt3U0t/
wUGhgqmrRTFbjvQX8yTW0iC/9sI3qrdVPgSzYbxryFexnuqmjhq14bkD1GuC17iafW23AI2PYvR5
IWkAL75rIY9P44AnIOaOMIawogQhYBAYUznvgCEHl96ct28aW/ayz5ryJdLuOfbYvKlE0pwgfBc3
b9UEBjatPq8jrq42ZEgHTn8uEh36QbEdTODuJoxvI8pmkTpwJcxLgceDx1zsWhurc4Deal5jifPj
vVL34sMbkLiUcr1wxWzGiTovNIh47iEQ2zehwpFJQi7grg2Fkc4FobEEIFPXCmFsmeFxbOZgrEeC
FuvtXzHYvfJoK51B3FCak3Q/itj5M5QKujkGap2fFj36Jm58jgjKMiI7nIJOxfZeLCNJyf8x/1UL
mNDa40REEy8VXa3tYn4mYWKLHTcBKA2CHT1i9P4Cr7xvw+ScWaHXbIF1STXLDYyEICmCPZEBSgaV
tYd93G7cwo2g5Pgyz7hnd+VebS+be0sNjtI9zguKQGnE/p8F6K7Fr4t22C3AsH7R/gs9yLlKQZbN
t9I/dD+PUtq9dwH1TYwDjDYgPDDlzJxBfZTlzMV4Wyp9057R/WPdoTKY3lzuoOvjqHZ97KOt14Ui
E6CLIE9bOsAo5G5NIynq650dMrrcyYGvr7zak+vNnwFy7JXEY2Z2gAram2F13u8bPYdZkodenUyh
OUjcSF6SfXs/Wby+j/Rrvv4RhGZWF7xFN820mHztE6LoyXYY80eLq2VIhHYOpdYBZT6pY5pOa6l8
ahR8lN5v1SE05bEd3HYLs4w/m2t1sLd+DIMpc8vYLOihZ2j6VdFaDkUjYCNjE6G/zfRUhyY9dHkj
AGltSKtc7fadL2iLfWYS6PF72tcpnGZFOXJChCMNy1ZdNI47BbUN8wHhI770Jm2Hb64UcJermGJl
R8GiHf0uUdNC+EaDBpf4AlDy/45FKuEi65MpNIr7m2S7SdSUfFXE7SrGzPJHTueh3GUgqqFcypN0
ex+92UbnwrNHf3OGCyuNVJErs5nPMxdV6r/X4wEzp2lHTi06RPHJugncVQ24mKuZ+YVl6qBrBmF2
y85BX3eiqJ/Q292VzLGRzq1Sj24FMpdS86+v+V3kDaffbOnCdjrQdErMdfV9PslO3xIjN0Hb0f52
wMV8yeOKd+Z2877h2Ngg/QjmhNT7/JqBjAtsh5JwDY3sszqJBYBgCtuI7W+ABAGDF1eZiidcRCFb
+0lIGSN7uX7NWSsifht/FobcOVWfY0wXWuOhC545UU6JIl0WedNgsC74t/bWWU/cWBpmFUX+lS6x
NrCJxrc3mRk/TSNnTKsZbgYrrKY9dGYuIlob2o9TKauN3nNg+J2inswH8gut+KsxeUSlu0pJ2lTs
C51iOmSRiSxs+K+fDLS3Wj+ZfiINvqhHJjEDY6EjdDn9+v4wZ8QjdTSLMTQhytVcZ8cbUEAIWK1L
sABeAJQVEas9ffM3aIbHzTNW9DCdH/X3fyiFxeu8rG66qBevD+eml+XVLYoe5SqlDscxt7CsC3pi
hV6xEEh/BPaFxhmL+0MgImzLUay4QCpTC9eCD+RoWhr1ONXzx2tQvWa98G5ffBMxq0dZkCIJE+x3
x3tOjRD6Hf3wLqjf7pIcKX3Hik5C9yCUdQ7TlLwG5D2H0P0ewlcXPKGefIMNNYn1iG913tsPSBvv
04svAIRK8EKN7gv2O6oOG/aDZqRl6iHqUycwcltHPwpaVDQ+P03GCBUKHAKg3rckqpNepCWwovei
qVPEqQwwnJhkYFXIoNhXNm6+z9TAFgCvh0e4fHOXlN1f4kuoPLsO410Z5qU6/y3HcquA6rhD8vSo
0iFXgsJGGJ40kJKuSTomDHjL/DdXq8ixAQ0oAc5dMaOzqbVaYJSiCu4Z32fg+pXWytzXklyG9A0u
GcBm8Ba3mIEUogwwAJByp7MQ4fMs9pTpLa48vRl2TYCizvhi6WW7hr3G6XcDJcTnrvIFX856Qo7v
B3CVR+YfroQ4Xktmj7QBxpPpQ/3x9C2d4I5HkUiB+HYO3WLHBeMXUMsYoSap+75evy6w+KJNk2+i
AcLLw7G8paV/haMDv6GE0x6R+nTui7XzFM00GPdkKOBHvIE5iwl/WFwucOVuBnz2KLmc0R6fsTlX
ISX5sd/BQtpHCgCX+ypL5kASCzf5FPE7J95gmZjBZpC3AL5Bu92EPld7BJpfq5HaYodUufvDYA+w
VE74/xA2TvlVFqlICkoGewSsMnfILs0J+NAglgv0wAYMmLrcgjtNW+dqJOuApZnpJ56Rg/knHwUl
yfhn/52btI/sKT3G2l2yLcHTeKdSTPFTGWcxRBvZ5mcGFlDiI7kkZL/Fi5eb38wpEvEmemLit+GQ
iGOY1QOXC+BCJnizsEwSWp9r9tQVvZ2a+X5Lhw8loW5nI/ipYnytlDlbI9gI1KndpBCRWYSkd73I
7s2Ng2XWUOIey1EoaVl9+aef7n82OM5R0Nq9a0HF8X687Tlq8TNsQOpoc3T3mFXyMtM12FKBYT0O
UNF2GQbORsPfhwJcZ5z9hA68YnUwVE60X/SNvgfrx2h6xLCr3vEyul5I66+RU8xG2ZK3c0lWhnqd
OR/rIWzzfiTR9SDYQIxDXYLAR63Vlc6n/qeSHGyeblU1Cg7vRQF6pw/OCyGQvh9QlxGMymCZFHxG
2wF7TOp8Mq5cHM82Lm1AI8HQtfMfs+Pee/BO0+2v06z+4hlHHdNkb9qyrv104pdfE91KAmuU1R9B
8oDvAprRNEyLf7pylalUtfzqCvE0kTBAtscYh2oleOHRRI2kuDAfnqpnM3CQyJrIlgSxqojVfxXc
aTaoc15kwRhRYcGkOGee2NIZ3xxh3y6rpuCwVJnxxtK7NwXQPbAL+X/17XlAbJ0Ok78tqa8Nl3+4
EnmSRXPvANEq+VHTFK+oMpX2EtRAVJn3HVNYx8P/xQ22c3QwPz3R0rJ8klJ2C94AnwcztQCF0uYZ
5cX7SfxrF8U7jCZaXFQYJck2uQ8DZkVfqtIFc1Coi1LqijKObBr6t+LnGmX0p5n9UayllZffH9Fu
PEBco5ohijwNboRu/EQaK63QQ4nrE+3zE7wCaOj8N/PYQ8If07FnsAml8Uoln3nhz96MhLMyRt0/
IjwTLlc8vCTmJll4l027kSX70b2kTv631YGvyjGf/6M0ggRrO/xVta++cSS+setiXl3fZ7oBNrqO
KS8zD5aVPdO+dFDhTpdvXxQ1WeExKuhdihdSn6t63SRG3gpoHXc8akZEo8zMLkQdMsPIR2UWhG+m
H2ZKmee1AqxFx7SWVnKX0gxsMuQjKW/KO01pmWXnff63gYOPxKc5COzk7HdA5zoMSJOQd7W2+o5L
Oq9VKK/9P6TT2H9y6Mp2e/C34rlvRvSItc7DfNKfTWvboLH58sNfQm+eq4w8g7cqUl+oekwZg3zX
GqZ9XFJL9M2t3KGtfOpkA/B197NE4jbUOkqh4b00s/X1Asy3xicpf5EarzeB8RghQhfLabzxIjd/
OvPetJYXX84H23f57Rt46MsmqWnxgmcpWy0glg19fDsHZO8onVGqUPS9a57JtWdXrpN8CNjw1PHI
fcm2wiAC107X7OZwOOk/3b/f4gcaKQiXWPgZzl/d3Rh40A0nCksLeiRVM1TcP1kXN3RvV39XhrA6
pYXjHNZPtsg2xq2UuoRP4jZSQWKflvUVnuc/CqUOOVI/rCFYfg2A6TK8dQHWHKaomsq7gcUxm+jw
Xf8x49tL1bHJJpVZw+a/X1IDISB7X23xr6INpuWkpXiVFxbu6bfBoRpTVEi/clK3oYJRb7je39UG
A5yGL5MRrgEE/M6hMUFq6L+90K8Nkfn+oY4L/sZ2kdXIthHWbtQ09nkKA58WcdcH4Xy4sG031MUc
sKPbXXlUg5jybLP4hHLMGxyMiVIFkcFl6iHN8X031+/BcG/T5hxA8PNvVMI2sGTytWQ1eazwQd0+
Ch5XUChvldYSsGRSCfjEkCtfkw050pTxUbRNv2dHum/hMMBeAL9n2kCG1eb7xJTEMr8nJH+32Kt3
qj01o1O83XnYMixIpKmUnkmY1falaRAFWuIW5XmL0jzz69hto80wyWYBcpHhuZItA76uABw6Jc7L
2EK416Hgj8k5dKC4++N5rpVfj/qb/h4A/Dg/5s0IgQ4xI1t+OnHO4MnzpoImk8vNTM6Vgb3s5PiE
aU6rvy8jIZJYq1pkl9KmFG898JnmgbBCmJLzpXVzs6J7BEpcnpwTkP4qMKzZPpM3xHOPbQDWkPFl
n0d4G4ea7FljON7Vtths/1lPg5qhGM+6f2tORXC9FnQwgi8HCHNnKDUAwM+ajv8InWQ3MymGeW7b
rg7ePODxZLmotErZmnvvYQQYC6aWo8dQ3/3NlJkBr54cnhh6CRTLkbRCm6I/C+OH9L6X8T4mR3sV
TbKT6O8SwY8vO1lPAAjvLs1gUuTHm4RmCbw5aMb0+xQPYoL6Doq7f0uNQ/88A4fzZa3tecyOIA5q
To52mcrOSa8OX9XcFgskwB6y7kT02VI1w9G6LgiMNBCDV0+UdVM0MQ8T71tG9kfjRreUZGfzYWQL
pyHgODNp61Duk1Vacho335U4uRro+W445LEp56P2SFYifDMJbLDXfk6oO8GRwYhAtTYihu3+Q+4P
dqooni4B8uodISkUFie6RhVY4iGl37k+YTbjccbbFr1/rl4yGLQxZ/oyjF5PaVoA4pTsPPrxeH2r
JvMy9TpYpfT1eY+zfp87xDvVJYiCLCAg/bpTnBAFulX16rLzDiiXFVcJ+en/DO8DAL+CHjLau0i5
9gbp7gIe9zNapS/AKN6sOAaJXroUeprZvGdrot7FXyJgeLTabgnBibH+2tIQe6gOXxUTID8ZsBjo
anbylKijHL8IIFlfeiN+c9bbqayigWHuJbRNZZgc1i1SjluCcfzruaf5s1hBBMaHoRn6S4i0EGTM
2980+kkVQteNknGovUMZb9er0OeAc/EoE8Sb82qV3/cDxFXZJDrgT+ba9E5nch2htOBDMNYv9LH0
RHezKvYuPTWf9GlP+PFfkV7e0t4u4NSyPBoeYHEWV5vy4OZw+US0dGUKtox8m2NAfksdHIL75maD
SCufK7nFk8Dp5wZKYe5UYVRnB1fhglaOgu+81VH4Qh+kkj+rdKVZHRVp4DG4JVYFv2YslSey0RHH
GsKin3AJY3ID+Fi13CC2qHodI3fLypG5R6dw+5qVqPathEN+r1RSdTwvVc3QESJPJ7runPfLxeT5
lBatx352ymQN+H56gtJR+RtU/oRW/tbVRS5AaNFMbI6q4GAL8uc3qcHfxZVLIDYDxyAAioduaZmq
ugTsEmLyL73ERmYx7VgdBR19hks+aoxTLdz5PiFXePPXEEhdooy/hLqkQHEVPHL54AVDn33c4BEu
3gN+UvOb6hM4hQEseP3om67jjao1C0ExHCS9iRzEEwXTJkLh2H8ypA3JDvLaU+rfRO+Jgq0k2ig6
kz9bF3OXSWQYmNfAUA24vSmKeT+R48AJyN9aPxsLDMPyDe7lsxdRhBWv3WQdgIWexyS+hRaXe55g
/HlKYKVLTmVaZPvyIelVd+YuFxWA/wHgrlM2j48m+xZhcrR9rTYIV/+C4IJVtmFRna6Q73U2fwhJ
R9VarTfQTMxVZC3U225LyQ1GZ0PNW3w7bNB//3RPoUlfzafUWNYILySsP9veGRblLr1arvJHOKtw
YE+M1WamltioJ7VMI58MHK+2QQOwsvBjoUvZUj7VjrPDRzwgKtLKBM1ikwOauXXCoI4+X5QdkPaf
RKvWTs1Wsl0xeRYRoslswZoBHo+VG/wXqsWqXWCyrf7+XW/czxvM5N0SbMNLyMNFwMxz+D/xY6UF
IP65zGhVw+RHgrzLmGZKTMIJHlTZyeFUlHBTQDkzJpMHdLFrrCtVJEZwaqMjny2pU2vgkTq11tzF
j6SaAET1DEL19SqRbhi2DH0XjSTAXCkGkJ1Q005IDAooI7sGYLMMqh4Ge0+WK3oXkotub1H+/8AA
TAhAQDFSLvKKvjAM06Lf+Z3x0Cq8Wl83/bHlPnHgaSsgsb/qAT7F3TJ+tkKRyYz7SmU5a6TWriO9
PYCIPfMa3Kcn/PFeb3RXQEvC6wBTaULRTmDIaxY6VMFB+U5DNJqBY7ZhT8lpUbeYi0zofgakQVwj
EYJDbVk05Fem3nYHxBbfZ1sQ92ZkTq+nAQXrOtY+hFJdqaPmqpaPYo5qiDQsHGaCnpQCNeiDK2U9
LXTb6++1XdtkizagWZsottcySQOdVETwht5gHbBrkXNFecmWC8mpObR8YsXLMXB8pCRvQePE37RI
yfk7rkDAIm15c92S6Mp15wYfjGWsLY4cg8KVOSATqNR1PJqUowNu2WDKMtxmhYixN3FsyN2wULM9
0TfoSTPOY3yzwxX8lx/1xDEIXfAqWp7G3Q7e9eFv2qMXiDGboDuJlXtgodof/hljBQ/wtKyqWALj
LW3dsBJ0d3/Ih+dXV3dQhhEV74GdcFIHz5PnyJwdzUyPQfKtwZhMI4Yil9WtOhbvlAgTK9Lnwsu8
FVXHfSLDNLn4bm0lsZ5T2TCmVoKIXCy2x0Tfu7XKDE1Sd6Y2y0UVAv8+R61hXbcjgN8J0644YUtV
pAi/ZcUhEg7MyeKvPLOzlRmFC3trza7j3kCzcgPm8KIqSolZmV/og4BCg/K2hJd4M4OaYl34Qh3+
gLtSq/NqhEr9vbZtKqF1Iegz6ucLF9hd88Qur5ukxUsEcZq9NHQh0q5MzTldm1XTNC1SqtIfWw7u
jtAuE+VOjB7DF72tuakMF+fvRzkxMK2d3z/EW3GXlraNUOCGFTobEqhMuKj2KRVuhQUtjH9/r5Bn
WdQwz81zIUh3caXoqYizDfG9YdobRRto/JIh0bDKd99YJ+RpWKt+PghGAcYfNhu7/Z9oCOfYejeb
Z2OlQ1bLFyUJ77MPzXLLOD99s2R42tKjNCOPA0syBfqgfTKhDUP+OdoWUobVxp+jn1SCjxVDZebc
UFauwxtz/EC/9oy1bjIQJVxfCfjFf7jv6aqALysrRpkKRznoLNJ6Li9iBW+0l7xqmm9YNdLC5EEM
2UcHDO+wZ2sobyLlAXYq5Ux5hIJbwiXsu8Y/AVyuvyRrHC7oZFzRhcEhtdkFwccCx4Su3TuBCmYQ
Z1NoTW+ShKkKlG+vAm/FfXRSfF25rxyUJpO8iPVIcjeXCVP/vV7RyN2KkSd4zL7lPAYwvQEBa8R/
RweZbDzB9nuX0T3qK0JkDQnkq3HWWM9E2kNOmMTzZAOWculoawV6nEOhMvEHN2G2p1gUQfJ3vmN+
NSbHIN6h/FWXQWGXFH5JQcTCh1pQ4dJapmDyeW+lySg3+enNhdTLL+GhA0ts/UOPOe+pAGunGPf6
GuPiTT2G+mDKpigKQ8B0BnFDQyxb5OmpW+Yh5Cwrch6cPyG0r2uM4Ph8s4/tWRqgrYuOUPeUS17S
dHqmJoaR3f01kDG9nyAfK2a0NECIJ8WGnQ0buuTkEHmPfFEwn0mo2zCK30iBNEw6rXAzLOwoQAWB
vZJRbM/AYa1XykXG2KPAD0BVHzv1NcI+QfgU0T/rLz8GjOsdTbnUIH/RSCfbFWmZExfIou5W30wn
q0qh0FUln+XKTjUV8E6KZGeSkQdSza+7BSbb9rcguj5/nyuNEn8OdHwOcND+DvmjGDo8KSGh0Nk1
kXvDNq2LOmdfklGmakrLen/3Gh2yVYsknX/x8pwot2jzdK7C231tH3LkiMLlNxg/MeWp9XG6zAKW
8NE3PImcISwBM2XFCOcZJRgEeA3vetbQkXOeR2HTJruWEk7Zrt9OaJiCpPbax8efJP/t3TIRMhVT
RphNqnHH2Oc9xTOwMFZ/DRu8EKEt8+WHhnVSiN3Zlpfak+HMhdG8EO28e19M6gKb3w34Qo03IgRd
bHDZW3ozE93LorzsK4LIFJZjd7Hpu9qXjZ6N0EVkg3nJd6lQ3FIFzwwq3dGc9VjBtixWOspIFteu
g/Og/+hzm2CyztW1UBfhZIXgMXBMZB0Spnpje3P4m7pnJOeW25DeBuIolNGagW6n8xKt+AE8DMSf
L9xFcB/Oib60XDOyPLdsnyBfDhLK7omui2xu6uRntD4R0A8dLYNtWy/RX/kEE6R4N/LS/HPG90KD
O2PAfPgtcQXs0qFj1plnajrh4zwLGOwyKhoU0NfkWA3fUALCgfWdR5DRwcBQ0i76z6yWWrYVwAat
cTEAohtHpehLUZrYtJuzGnN5VcYLsZ4O7gPqBKINaQpdqBZyDCNP4qkjZtF85meJ+VQeT2+R8fOj
oSGEQBXAdC755MJnoVGZGLSoK58terXr9XHIaa04UDKHfTA8j5MyHbMoxxmcKZU1F3ZwFeGhQ2Kp
bl5UpJeY1Z/SmvsMX2Ke5jQtaD+Sm/q5El61JSbBzl112G0BsPOIrUs++iF4d3vMG1yhx6zBiF3h
zjwcCVjmmKYwdssoPSDe42x2TVgb7KiIzIXZ9Q1265ckVgeGZzIocS7sAuObOIp8PeU5Dr3AQ4uT
TqFScRH5rWepLvXDjTqXTo2DJXD/UKjsI/9qxlo4meFZTj6ruCtF85OQZtzFfTf6AQ8j7McoILMx
6NXmOTD7Ch3gUgjdiYOO+8d25h4npflFPaH/tBrp8oJlz4ECIcNtSeCWSC4RJnFTt61eh3lKKx4o
FybICuRsP6RSytdR6r0mg3rIL/jjXSR1JO8A/qnBrqlmmQHAA5+7GJ3eG1ivvqRrZJsgLRNouB+U
h6vWkKlPXZdOI9xft7MGIqfZxfH5K4ow5YQYegC1d/8pS88kGkjiCt9vzSNSz6ibl4YqlPBzWHgF
yWoorjBULqlWmoby6xxwXV1ERlAALJjP3OumBAqbWYrfIR8Uw8ioneN3JqidC5jvCUD0FfQTT26D
qoz80aHOoZngoD4W5GNGyvusKUKw4/tlFaZpPjq9oB0NJh/+gFhbnHSEHd49WkfxM/Xrx+IA9hiW
Ol+9GLOUlo+HHVk8H8j/K1mDXHozPGX5AEERNrd8JGX2rHEthWRST1hhyhQcfG7IeBpr+OAa7qKq
+6BFQ37SDcvZYrjyPiN4JFFAdnnePt8ZRSBF4F0HFhcW4WKEShjyWxPxafRtMO3i2tGYKJuY9pdN
WJAGsV4Kez5V6GiM//xUQe5srYV+OCHuG491Zh+W5WTfedslW2RXIX+hw0DMrXEyXfo3gES8k2dw
tpUYx9okV9z6We6rBDCRsIAdXdOuICwLhLsjxRrUVehASF+8Gk8pcE6RBEBWuOGKuu0i1FSiOpU6
7ji4GtnCNVeJQPQIGr98aY+9kfSjVuAk6yZCHcCQrRj+uRpWlU1LUN6cAQ+v/vxpuu71ZFzWE+6i
FSbejdqldrIWwG4YPqqdiRvI4cSS3bjqzhHcHu2pNvdn0hOCWSFrDF92beQYzZRPqfT5Nkt/VTBr
dVDtPJ8gmqr9IHFQNy+SfZ/D1Pbm8dgSm57ggz2s5POVeAJNoeehN9B/fmUwUUA4jH5rG2GWNYhy
Tn2MLriK93OvakUj6iS0EAjgCtxNIkDm4eP9XGmk98eOoYCZMd+iznV+RtlPYU1SaHcY+c3grl3D
L/AWXKTdt+gLxChy2dZ7Kf3b84c6uuv0J5l3p6CfNMHiI1IpX5OFGnHd0sEFxwtIl9w2MNAbk8CB
Nd7TvIogVBu1947qRK/L9xTfXWcgWEVdqED17lC9Id9lmZNDugRgqpw5kQgtr3c6Zjql6dT4RWlS
xTMHg8mI7Axz6sNTZPVvNaKkp1v8Qt0bn47QiFHI/EGABdK8wqkdgttfGoq5OIC8WWgiW3c7LJtH
hbFypCSbttJrdKwPJbZdP8A2c/hjmNWp0ZFBSgJONnWoUiFI9vnJqeBdE9VOQPXnEKuFlXIwIBFB
O8+CIaC7tdJsAkSAGRVQYrY09QO5/xptRHPQ9ucXxHQ+E7q3BEfivhpTFgeXzkq7uL0jgS3hUoej
GEKREfK6GJ0mp4nvtvezFqJMf4780nvKT0iElMYzi+msfvrD24t8irasDU4HWwNk/F1LcSPql6p1
G8Qgmi6G5M7v+LceNEVvprUkmpK9dF4uAsofMFp4sFD825JJZpVEObUkzevQKSypLFz9BWXEsEPE
7gNShk9w47Tzs7HLmDRZBA9Rnf7pUQAQbIon5s5PWCoBy8O3t/ZJWh0EDaA+hhEqyA0HjQicJL91
ZtgaWQ+XQMN+6AaXpMQ7LiPXNYEib1deZx6o6Ys9KMjCIooLX584eZxNvsGW6KHTKWJvHgLyEKeY
O0eVvNDwtaJbvLtnPi+th2giuckITMk4kF64XbSKOjgNcNKowB8W2ZPlSTHrDdoEVJ7CqGjYqPQJ
lljywOoV0Y20sxj4xfsoEcGKpN12fNmlJCKloIA8JYVHJdcn6NfzMYmsmHaTtz/t7UL7AXgj9Yys
V5l8qHi5tw1IP9PsuWnjU/KLr3VRuV9uaU8/kHsI0cE0nRPbO+Vivllos5/GSxMs/vmD0ZusXjwN
2jB8n5vk2tb5u7PNlvZ0/1jDmLNuaAGSBSBMaYf/5Ac93t5qYtmPYTUOyA2CITOfk1AtfOZ3hmel
/BKZH57a2qdM9/Qu4VJPhw8OtIl3lYYfBv4LSJOg5rSSr+rL7dF16BcW/wK4JuV6WC2Z1z0xBgzs
JThzUBnyfL4Gn8uG+B/jwDHSFrRJgocRlx/lB/QNwp+mmpNYwj8wLUHY4kqwpOjhEq/0Tm3D+4Vj
CsUQMfz6yxcMYvpgU2KrEHqruB8JfZYc8dMq+LyFE1GqV2TQ33VbilpyX+ZIjUm5GkjaXuZeA23+
FiUmRDIzeBJejeymY532euHOVw20dluEpTui9tO1mNw/8PaP1vAjaQIpPNO7mI/0TlDIGu5uhfcl
J3DX10pObmJANeFTGEHNWSG+YT/TR6ELn0A6KUeQp3OE3FgBW0a66RlQbxQE4esH7lcPwxvxKTZl
lqYelh7Nxu6Zfypplj0uC/GgICRDJs5Ipd4XtJA90Hlvr50cdFbgbAkdCqK8WawrPA6BKu/CNDbD
4cR/fn4gIst+DOwrU5OXUrdQxzm/rv9jwqROiF33S73u16Kk/e0S04PE6nJzyTD5C34echc7IWhI
9TZs5rOnB3475REGppizpFTHzRzO6jSIb7botZ91B2Ah6pGENKDleg3eQu9xHfzHYFbrAOcYW01a
jjZ4Br8u14lPMx917cTxShy3Jsvd6IIN+srBusD3JnimWayrn8cFW3ip9aPFMt1OAdiC8IqWr91X
+3QjrADCQsMWFVOKCBRjzK7+llfK2PtSgG76hyWrJfAwz2zB5uZNjGENJJJU4CLt6mn+ei9mFJKZ
BoglJoX2YTqSDUku6OOcDaHoxlQJ8gvsm+JLlGKYoMs5gv/YVx7EL/LizLn46jctL4D1iQ7INh4u
+BB2vNbw0ixLCy7UwLwHnFUtwHScy1/7+aSWJ8wrH0OJ2IhyS8H+CeKIUC86QmnmnThJ5uZK4w0y
C06MrsvMqaMBiWJOyip/wdHLNkLQjpuxnENTvu8INO7yfsXQckWU5l0O9sWoio8ejDCo3ljDKNWF
Qk9H8lRNYD/CdUMKb/QSni88y98wpomYF6vabS7ZI4a8T/aRUSlQitMIClJw7FhtkpfqXn56fIRz
y9dlkq5VZQJcZvwRErNdyBEbqIXtcho2CiS1EWfC3y6H4t4O9YD/TCElt6LIGmd0Fd0JPqL72Hd1
kzrT6waqPX/imIUMLbv06ydn89fXXMQd6+dbvdQPDCkqtFJ+cqOrMs74iXZNgGbPRYPfeXvUQu6w
AvK86o+NXQYMUA1KqZ7zcX4cbfCtvNDdUKa8HmOI0yiRHsxcw9UAIb3s1yaloWMEoY4If/PJUGFb
IabNcl4kg8DkxRW2jKhWK7FkQJRB4ZKgej/yU8os5CgmUTJdWkUS2Cv9eHv6NQBBnvY7uYwTqS8Q
oNSsFqbtkRTB9qFVuvXsGYpWQoAbc7CSRiqW9MmV6wO+pMK1PKbd8jJZn437IUtkvcPzA5935DlS
z0MbIqX73k2OWvGohhVmx0wW6Dwrcp4+H0lz8xgoWgfuZQXprhEw0KxKz+5dC0VGorrdASfXAYq1
GB0Bb6sjZViuFne4qiZ1kEurYFqUzXWLqZjsS7a/pn2vB7qhifhH7ZCjqj2dDlMb0yhPbhrMe/sH
VAfiOgoURSH3LzEZMratwDb1r5uNETL4OVQVNl1QZkJzB6qqpUeMTtRSwgNFKLBdA7RsPpPn1qlg
Ci8q6xSwTsgOSAM3q7gba9HxMWH+wPpfNzk/w9Sg96DClxhb8s36ypg7FxvNgEVNpSBFAaLsdkiN
WO5NaQKdSySk7dZRGXkeNGVrxA5EnfEGEuVsAIMcz4uxyg9QrIek3klgYnmgkFwhP3kOMKvqay39
WyzmRUyXxF7Qz8kGkqOnfDJKCOm8mOIxFIeMz6xxC0LPQJ54TyJWR0YwHeSbPQl9m2iWtD3pXGRp
ehZ3Sun2JhLKB2thZjdtIqZ0QJUuMB6Lta39Omz5UG3BUulC+8WRzUwgIii2bspPidbm8ibqW2dw
uKDKFr1FVwv785vLMdNdBiYFYHGiOzpGTaZPhg3rCqDYqWGvSGhZ6KS4bUdnBczKl79Kxh7RlzpD
dvKHeT+2sKJkOEbhHWXQa/EA5t2K87hdfR4mi8jjg8xskZAECjehKCup7Z6+n7hRLiiezsEdjULN
beN8Xus3Ook=
`protect end_protected

