

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hYn4T1Tz8lmB8loeGYuHmgEJp5TdMkRKn5tdK0Pxo3wkkBR/aG2es4RXT0Kx9IkGgy2jVWVPoeKB
usRl+M6Pxw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZOTsELKZdXMGraSgAw9rgqxvSLbW0aT2lTeYBbmmRdIiILVX40Q3XF89sXvrmWq2q7dAJSXvpsX
1JIpxbCUMi40Nuru7hdg9WkNNMs1Q8UJCou9g/GNLxJnh56Wx2JqOiplBqlgeaLjd0T16sGmIYm4
kTNGsNPOASR/dWaldsE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o6ehD67QiTZFs1auOjL5nkbDEbn3neiXmbyTqqoQKK+v0TaPL6hSxGHE/Fz3NtmR3RIza9+Y9rVH
Je7RNuyq8vsgofAGK5Qpf28P/9kF6eDh0JgLJHOonk7lnG+gufS3pMHIfioCEe/2wyoIxzbwUPNl
TCIJtbzDvWpcCIKBgiQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cASOe3RHelXhU6s/jEEqAnadTjmj4ihjbMuYb8YjKT8lAROht6xaHEt/3WXUlUPXIpDwtJlexClV
csQVUSlNShzZmxBI5epxH/HJqLhQYwkRDFK2BUAagxn++cS1iWJGlow9Gha0EU+PfllVje3OWy4O
LbiqHgQlEG6sIGo0ZCj6KPC87SBAytHtAiVRpovpGAxLS/DLeXSJaavSSwOc7nmWFDaNEi9dJS9i
qixZxDI5QNaDp3uaBFLzKqo9oSPgNj1mYKRZp6XL0ganfqQCHh/snCyymi+o0DC5vSM/+RtCZHXA
A1u3UsiXv/IfegAneXJ/yU2Rpj4P9iaLKgmtjQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kAlIhoAHksCGo5mF85FXcP0dM1NExLuDn6ZkyfgoWH09b5qcw8bLJnQMlkLvdLRrczznUPKBLrRR
nUHSMi9UTzRZ0rrnazgGnHFEV1vyoRgDQDOpkZbrkgl/VynbkoMBhCQXYT59yyHhqjI6WeIYVipR
zyn+NdmUB+/GwlsSYygywX31rotvUxb4RZmCqg+UCemw+N0tS43QuIzJuG1JM+3+SVbU3LuVcClf
rOwWqAFHsOXBSrXNoPX6QeNlYUKy8gcjiaQqPSrbrSJWdgvqshdNnvLWuzkREOLY43TCoAFwM8p5
73h2VUHmwffIqzCELbp3Tee5sQXgMbvJ+Mbfpg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CFQ8408huN9E8h2/r246qkePkogHtf4rd5gf8GO4NiUzetOQ2my8cbvxYBjZy3yQSw0/LrN95Drj
cc3uAe9r+wOvBQ3aM7AKnKpRkAvmqyCRt8lkW5NRi37udLv8jQJ5gVByTJ76KIn8s2kfj/iHou8+
VyK641fcvp2Fk/dmC13HALsHzGvO1m9Kg3zHT1aJxtdh2FDGLhOy/TtcAEbSWUhNkclp4pw4r97T
urhhIiarPZZDEkAXG1Ezi9I9ebmvdHMRRa/e9P95Xg7vwS04EHfmVTpFKF7UHncoI46I8za8vjyZ
8MCKLS5zKbgCU1OCJ9lQ6mJX1roD79pJrnKYpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
dONCjLIZ5qnPblgXUqjwUSFZn7UKIoUsVojLyxJEfYr7T7cGXhclFxIhbjPpu/hL0iFJCzyd9OMA
S1sBXaUo89wBeRlZMDiqkxghl3EfHAUl/RD3FYcGOrOrRhy6CkykfMIlAUqUrnoU82Qqk0UoWzjy
HzQmlI/mcPJCius7vRClgLPu2rb+WrEuAiySAv9ZnspNFo3rTrwGofg3S5S6wzQQAU9xp3Opb8AW
JtKrAZqHXG4y/z7xX85PrhMf+lp39MNrCu+0GkrKP4ZwlaQz0Yx0Mk1k5XJeVR9pfSl/hBuIoone
poFVe3Iqi/BYArPch8UOLa+94rwXWS0CLMZgei5WlIX3cWYF+RQjGpQAhJ8O+MBHuFEjOfkUSLaN
UKCvY5rm8mraYWAz7LCGrvYqygX7BOMjYBU9/PI4nH+m42hlzZCps65IDpoFMVtCVfPH5+ilDMrr
LxljmNdqwNPluRElykBhUxMY8hYOg9VW+6TsJjuzlDVBKDBiWRJJFmIjWsybuqcANV1tjb5KcNm9
mTqgeT6cLP3QQZJY917n73SJHbcrzCrpQecLN26p7AHcRvk2yPzMbBltIWwInVooy5oHkhI8w9IO
SU9JC4DYX17R+VDFeycNq/+3R10oMbzMhqKQYjqBWTHBkaBaxmKi9u4evG4j2dvbyrPQYIaVT46K
K2kNEPJ8qT3YZYZcsh8bxC4nVTwoK5/TbeaVBkSXHevMGbAxAbsezPdphvixvwePt9WK9oitJOLy
ITTgeyqWbE4dKr1fWqUMNIqwWNFsuQ44R/+XcWW0AmKVRCvbXeZr6QJxph557TtJHjdq6CqIEtqW
ETQk8mMIBHDwIOQZ22hOX3F84w/jvHARP5cux5sw3VAtUIg9ojG7ayNgpk6bBx3yJ5gr3Hf01w4Y
ItE9l9PXOn8TOSxcrvwG40UC4odTsh9T4udZN2mnWxOli+SJJss0mMF56tHy2T2i3TWw1YN/NeIx
dh1RMR610K71LsjRFa4FwKQ4KL8twzcg1K6AIJAhGAKaOVMdkr9zvrZnGv2UWFk9Gjp3VQcwwDsS
rqKHdXAgN+HKlS0S0ioaBUlv8vihGHxMFYPF8Kcy7GaPz37UyD+HiCSMtFoQGNF5Bie2xJLl90OL
cGj7NOusGNk1pT/gaKZfEks6scOK7YhA3e/pebMrwnSsZdELaht0TC/jq3vGma4GYcm0uFGFMQFm
x0FiLgdKJYcZak/3RnyL2IWayW8vPZdLvzHQjj+hutnCcX5N1vANbWLgRLGK2wr/cKNqvBnOVxzJ
AS3NRG8ZqWeO3jLpTXYde8ldUjt/RlpHYFs5rJXr4sUW/e72wUFBTKMzl42xzYgm/3fMpIQeXk6n
QOFqsVF7Vfbnx91KegX3YhT/tm+fq/wWgcMxrdUBp5fbW/etN/w0j317+XxNWVYqzSi6yhVXlGes
/Jur64USZaS1diVWRUmoOpkhZrF7tZqOFWLKnKGKrFBqIX5T4fAOPfeFGPtwUSjld9Vj/PTUIPqX
1ab7TloK994DdgshpPY0XmsdLgulRsMFxdEJRklY8j0vvanPf4XojDPJygvJI6RpOQ8NGJY2dSt+
5QxKwo2V4rwCvepVFkEqAvQQM7zhLglV1pwdUfN1kTSgz9SPdN64eexegFoEwicDdS835llDUPxw
ShUbNm0lh9XAmQB2ZWBPBFdX9wmNrypg2UOBh0IMnY+ube7BfIVyU9IQ/UXFhktyI17fhNkIUIyV
aF+CunfdHeZVbCL0QpBiaSdL0O3Ak7yXrqn95ciMRKAHWjtFkNRnZX5/W1gWb1bXLxldyoKerMvT
7Trawte0y8f7xPJNF4cx5jTHejrSAFVwGVIuSOgSwDVOOJg9MvdJY9Sgd2+MWRnK2D+cGa4rgL9a
c/mxhP0J9j7Dp3i5hDoWxXuaNMAGodzxm8YveTxfYqKJVue6/55mBeAPAShXIRjsou8dbVJy2OOT
1Q1Metn1bnsv6Mt9enhuXeKfYvHP5QDPN1z7d0g+r1R+8ExbHNDdpVAYoEVcuOErtzwti6VQX37b
dBOkEt+d7z2k+3i8tZKn1NM53mTUVjgGQrP1Xlef02qw6AzUa+0A8zinEFM8a02FawKJBGgtQPGR
WnHgiUQxqsoZuvwYJaeor8qIsCtvQPWmaZL/HdetYGQ548KL4TlcgyvH0ipyv5Y4lQEN1qTigqfm
44Y5F7HwsaW+TpQU7mgiQVzVwJVvoTsezhrA2gUYo4ME1kD5+5KNWqWZVHBGLbweeGQQpUHRK1TA
EVanLGGmdjGX/Pg9GLZek66IK06/caJmXseroXaoqKN36kF+pQ6URhWuj/PIeOVttm+MpIfB+GjS
Y2hhfJNHhuG2ysZrPgJp3IM+PNcni02RxKDHjmk38YO8wi18sRC+hul+2zFmkbBqyFDYhMAZNs04
o0A5PhAKsS+hbK0tRnuSeYl9fvyHwe7BvB54Q2aw+PP+J18FaeMA3cWpANKcoaMKtLLOQ1Df41HG
p3UehdcSpYtstv/hLBoevk/RO8BsRSwRPPdUdqL+CkPr/Zcbox+giS9XGJaO5qfogAsGe+JH5E+3
P4KBIyXT65Ag3/Qwm5e0zCFwTI2w9ywdgpe+UnMl11c4QOAo2QoKS2HSvraMJa5z/tXz4BuPoejr
u6f8XVws8d97UfOx8Prc+wdDSzxn3Cr1BR8+P+aiMtdiX9zcV53GrtmB0oKaY1QfHlivRqIyyHFt
Y+ndf5IsZc/hWdwxnG/x1LSxnBXYQIbBF4hXDZ8jLAtmqMjppQeD3b/m8JXWXWUfNX1ZFz9DFN9x
z/+05ALYJW/BvPVccE/QJK29vYsKz4bX4qAQpBs7uWNseqfFQqpMhMpGDe2RA4L5SfixX3vlVxgn
psRpwMBFZ0ffR/M5dv87QurzyILswQ+eyMxuAfjRROyQAlGtxHwleGw6KkHA3Qxx1yYrqWL+BPqn
cy/UiN8n1gZ8Iy1dfghMtl4b50TjfxUFn4izDDSqYW8FaXbgg/dATtf5SA7LLI9AGvQfrz7I1UGp
Gk2ZalWOjgcwcFCP1Q5lQRlci/mRXHpgp1wE13LOFlSlooOfC3DTWkPm8GNb0lcddtV9Uk6vrLvZ
Z7cwD8ZIIXx7bFvUFs4F1f8ur+3LF92BQLngRBi3qXAOUsvN0kPR8Woz8F4rhGleDAHqkEJIov8A
Ov0d8nQZmdwCdMcKoJYFyeLiaIrYLJIKSPgIrtotfgD89YR6r4z5usjMrnvwuc0QorVN5W95t8Ck
q00Z1b71kwtR7T4CH37gpBGW4cpxeePD7ksaVXph/EDhKlxRVUKlEM/dGZlMpZIxDDd/693VVLQX
2tRXAL3KHVnTYI768H53mMl4bJ2XTOOH1BMrL+Nn0cPvpK8Y0gNPAqbZWzWkcS4D/AK9uYgdY+5e
KktM5smddTy4IPcoEKLrOQql5jH2Nt34SFKa077wD2s1XQ56Ja1J0p0+99+SdVRJkuOZcg7tOJ+Y
XSfjyA0HDXSGRxDb3zoOaxRmI2ZD46dwIkMF06OYjX9PJf2NPy69xHze6wfrOU2d5mPfEye6AT/a
7UAd3aZiQld5X7LuWAcCJMcLrPHzwM5eaQQKlFr71AviKCEbTa2fcfrnuDLcj5IkYteTBOPKSuj7
u+DQa1HWak9YrI7afdUBOOqNu/06YBbBMVcjkT3xjvlVNI8vYcsgynC8K97o5vrJouH2I42nkgkS
WdI71ds++kwQ1UWd3XVOxVImItZiABSO0bLGAMvV4NQ8Os5jwPb1Rrs7uMV+fqJ7LiXeyRV7obpo
eqa2Kb8DHpj+eGOWrEHxwkPmwG0IrWgAEEiDLCPl12cbLFZSY9F2Xjhki/5baA7JYgx2POA2fv5A
mBFv1BMsDIri25c6vqqclogThe6AqV18pxB8XovuzetqpXwDdZD9CJu0LLa0F4WOyokRiLgGFLyX
2fmkIjsGmNmSabo2kCcDRssN8HcE4AwDMFcsH7ySxPmvxeJT3Mq4tJ0z3eS+RLd35X8tyy+/ZHMV
nDJtCL/u8DcbIOxqMS0ymLhyEm4kJmCTs+oDA5ykBOF0K1I6/IidfOr7wYDSt1nh/IMQDzw/1bgW
SyOtho8mrgknyI+eaX38QQok8f2ozoCpSiQOawAqdGqtfhT2zCnNncbAogBgJ/HL0mMY+LKHLWnF
U/4YPvK7hMWC9hgEBG0WlKY+6CKLd4k/8ZjYGunHrvg7XAjPs1M9wWVBMwqsdttBCZUZbIflMLOT
0QtpY8sd+NaoaukdppNwmtrIhKqb1aDc+zr9SQ/UcZBN/UxBO5VSsVODQBNbHV7wWoi6DCNMWgoY
eHh1VXiDseF5K5VXORFVsL4lzBuf+o35TkXrtateSXuUPQse0783zs1UyB6XkCo0pFtz4YlXxDcn
2N6UUsK7KYi6dSrMSLaxu4/JQ3gTIblhKnICSZWm2qxGhXT9Wd/ObfHTu9lfqt6Nbkc5xs+c5v7a
Uif6zKmSZQo+euQh/pKoswXCFY1tGyczaaVasjmFDQbwATHVIKTwfM9ViGAskaHCSRtiRiKhMMui
MNlIQES+XqpUkO+gP7g12dTZaT2eo4+9leP3FhEE/giGmfBdYwlBlVCvzdq8jQqfYcJMXP+sBisb
FP25+rnwVNYr+ov9xKLtVbXcTyYBJmWZw/us0EG1a7ok3u4J+SEffJjNn6p8HClOueyOMFciX160
0oRQ8EcQT3gTDiY/0EiFr+VUod/77HBUlvXp3Syb3jSJh4rZqwSwUvtbmfAJxo6uNjZq5CdA864P
Ej/c1VEjIoHITseHUdlEod94UiXR5byjwjClN9cZyglf5PnTQ3hZRaYAjX7RSm5Rkb2spzFzYUM4
t5ZDPKYdAtRPGx/5BkihfDO9NT/IYE6SHwLn1dUFVHkJwiuThrLWnaMfKKKFA71Yxw1JpgdpcOzw
sBUmZG+fIoqdaCYkgJ+dcPMrU1hxb109GZLaZQc8LiUvLWA1viudkQMoB1KZbdEsQiu3MptVr9ZU
ZZHP1Z8cj/hzXGMT8upTofri58FuVXFv3Kc8g4d1MxxujuqNNuRMWq1qViG7+hwICYuwga2PcDXT
fSgg+Tu46OPX2uXlpvc9h0E3OScAT+Dz0M9l4YaUfTsOIKB+rUHMd79PIvLa8ysmQmbWK5lykzz+
Hkfa++7vciTPUQTCRwR6Iih1uxmqvgsMLoL4rKUmp27Xi7hatv0vLiT4DTGTwXus5Sjy+AOKf2DB
24imH5WIwg2QyZ8slT4UqvNgBAayMstDSh6Jsng516o+4gvqGb4/YBwYKakU5FUinP0fUMnht8IN
PXAVICB9hsejUXzL28d+qjp8Tbs1MrEPC/Ee112kai2qzzt7uitRRg4X6zcDCvaaN2ENDSgUghJl
yXlraWoph5m1sMDk8KL7UyQM0SY9wTyQEw7dLL6sNJ5F6aCST7lRnX9K+5S97CFM74yREZ8cAw/F
0U+wycMvnRhh9Wb//3MDgzMT7LGDO29hhhmYjINeOjm5gblnX46wM5Y/0ThgT2oNWz2rRB9bTvI2
gC5hJi9a0RtoEXqKw3XcKXI3fUfxw+rbErn/GX1bnwGJ1SeItXtoNHqxkYHDZtkdumecStWtGtWE
awQSF5D7fNVgm9iRAj6ntpoi+bX5Q58fin8E8xy85OYB8MWBR5MIV5ZQa5WbORa4cOBq4Sulo7F/
AOSogdZtAtawUgI1qJ0oQyPQdpX4TKKuhD+sXUhGpRgklTAGRXYtbqTDTxXvmqo2/7zJcPmL+Lk6
Qu/b6b2dGJWi/xauTZEE/S/VmiPeLuBoV2W7mUTM6gp9RaJYwWs908zJZJ7Gk9+5xINcqFSLIvrv
M2ioiNjyH1M17yC9w/evSVQMs0NpgO582H8qswyJARVfk0kiXIaTW6y2wtcy/7+Gh8FzkICTa4bx
oU7i+UfhVldgkAzcxha9plJCWyBfWO82Je9SyXhYUTMgOQJWspx9p+amWdsanWJkm9aQJBnwu9gu
optGGFZnC+Pdy8cd+ejGq8Mouf+IGZDYF3QuxiRKEj7Sk4TvCNMQryjaToesqpaQula83y2ZebHo
cdrPE9bkJd4HU+goM9z6WppprKSeWqqt4WYID6hqaIYqoy0exZiRJx6Uznw1oAY8hZAhq5AvgqaY
r3r0DnfWX0kPqlhgsCUcgL3PGYWMxAMihGRqZYMCXylv5vDYo4HUNGSZLvYyZY/zUTqwk+kY+vYF
vvf9POS3bum05hkELQj/2/rR+Z4yHKgkJb4i3x9rY0yAu4iQ9VFUBKXia1aN56kaLug8v5xRNtGu
/O36fcOyj8ZqNuwxa/hfsHFW/PIQQiW7jNmL5UfLLqIqV47X6d/BD9CnCvNvEBS0hf+KSrtBPYY4
NU6k1Z1rSUe1CX/gQ+fvJtO05nGgKHOIR20bNRD/oWjxjb6ERlZH/WOBPfqhzA+OK1hETSI1fS7j
QyAXr9ZGkxPIW0wgmN1BUjO+YxnOqL6U6gelrnDmSi8hgdgHMhqAdrELYVaLGnMEByL/oAyyAGUk
OGRACiQVM/7tWei6iPe/CkzjHE+8NVg+866b4CPpboVYCmNdKr4XQVc3NJ8vh0h3/geCGzZCQwCE
IF+ocgnh2fBxDc+7ydgcvLtS/Tz/Av+mTc6o5vYreWmmMO4chOID1UWG05gspudyFCjvlrcZxdld
kWDnkv4B8tCOZa8elgoUG7lsLAyfY4VWGINlDSH7xdJ44u2Gtf94piqfbSf9Z4onCbSsmvohuXyu
0W+H5uv3wPJo7ZdrGhAsH9sMuV5FRhLzA+2xRN/FmJGqzRDNY5cJYMjNrHHOXIB3O4F0TdGJNZCp
uVIuEVGeU9q4JLBejv8XQGduymmwihUINX396by5uJFJfLzxgUnsdvDXSYKithGnz84WhBO83zFV
e/qw+nIf85P55ROD6Ctx2lCbehLLL/u4L4f8yf5+r5LAKJ6ZeR3ZuCY20PZIzU1xeF9XxJh2PrUu
yG+Uboc44pLTgRYMaDvqZJ6aDEUbmuXi9U3bSWjSRpxeDhl4NiBuezdGLm9wvW2zJhsJiR20eN1R
OAzwGuNna5R0AkizfMKs/Db2aAhQ3EMzhvc0qI7ZTymKofUiyNeHaUNDflPBulTlBmeRYpkcJXSY
tB1Q20XiwCEJJ1fFfBiYr/Wg2yXtkmnC4pqOaY7NwDExWmLQSE+NFm6f3wkArNvk1Nic61MQHSaE
DR5Gl9EJeyVl5P+y2CGWb4gJTbcw98toxbX2g1OBuV2K5edOea5hrAzVv7cBq++3LK2zcNC8Fmao
Ag74c8zCnFXLkw82Xc3gQppLel6XryE2+2c2njPDKRF3GgA4YijYcF19S088URaSL5CExNtJavbX
+fQNV+eEARgi4av26MhL4k+H53xjmveaBkkpG1eeya/MQqREQTXPnIj1s+lT4PTnqKeF9L8JQgxz
tpulIrkhzpmxl5QhSy38t2ZJ039ZVYkYtGVDnQU20AWc34l4jPjmeSkRWGRqLXsFLbjaMnI7HOQY
zCitf9do4Nnzk+7gGvOKvzroBFDOpQti/EVyoY22YoPBTIGzbBe53vwIFf/ZcnxffdZTfy+HBirE
0qPueMsrR3BukJkRiXC+FZWQtznPRJV0Le/KYYb+SZmw7USEHiY1NxjkiTW6gUBTxIrT8s2cvpib
Cu7PmZ7VP+2Hj2y0A7fz6d+FaGs3uJ34kA/lDEhoI0MxA1jgUJ8ukO+EYnHMO7PABzbRp93YSBUC
baPf1jeH9Xn/ip+3yjRfgfJBiYD0fnTT+1xEp5YuADEglWW4Y3HSIAI8dGjtZ/hX1QC6+XiPkRrZ
qG4mJIXWIssEL+p5GozDYh4LdznMrQV75p/Dv01gECOJTPDib3dh2i35qLy0V2jyvveK33xtr9l5
9W70vnCRLZYqU8AAJGvv38kK3/0UIb35WGKUld968JV3qr6I/PecPLJpTAUJGbe5cSWi6ogGiLGq
Iu2NYOyfldfuV9TsDSgp8AcPTjG7nVojWrYvFLXqKMpNXB3UM6Kkn69GgE04fzm57SNXbto+TXN9
MFo/gZFbdrCbJO/eC4ttfCy8LIr8LLFaNAHA9OM4aw4+SDLuDuUJn+CjuO1QHwt91uc8Q8idKWZY
NSgT6d+VYwbVHnohAahqje5gThmW7JXQPGJDrmF6SMbIrph7xYJvQb8iiZwTBgNsz/oZdP5CcvKb
z4llSKBp3nq2Tb3Uq9bFP0P1xkV+NtDAYXXz/SCqP5C+rCs9sEHXh4u1BY22Q6s4Z3KAg7bp0bEd
wwcij4sHi6YBnoYCjocu387qFrMhA96KWiyt+24NSNHPxtMiuk2RJ4BWGebtrtd5l4PME2NfvePw
Mg259szooW0T+F6JD5s4v03/aZWaFZnuM8bSvhBodWRfQneiLFyTM77PGlqaJDnvPPmNuUYSIkB0
sjXlEsZUgvvHCrqxOi0igCj5xl5jQB6dmfFVjKSsdrEzJRVd1qEiK1l8+ZhQriXn1M3fymWVOCDW
fkCiVGCbwSdRrImlgr8pOYNW64F2eXKg8z0FFbkvq7u/rXh6iEjSYMdj/NjRnz4BiUTugOWFWaHV
JmWZcd1+g9kSjCC883jaj2W0VPNC7SS592i6lVDo0uY7pXhW9p9lHAf3G2zgy98K995HQ9fSOXxJ
c/yOsjV07oqWVYFGZoz3wpza6iwQauIJkFdTjYQ31dfeUgEx9ejroOo0S3I5zDA7ESw/yzniIEFQ
DzvTax7RUGmCNRetrj4fw7r0N9oCPFbMZbW8uO7Ru6lmtE0mk2tFMdf2pI40vlLnPNnWpmDMKfgY
roCKJgLakuB0Ygn8NtlTePKSF4ZuIsK6BIm9JOFLHAYtDQSgMaWLzuIJox8+63otHLcwpyAL79SS
zXT5aHqVUtJkPCB9lQq82DvAkLA5b2+vRyEibJTjruSvId+km9uBrpXgI+h92Ary4KOw43j4dQSc
FMbF7Qmc/UDOGKveEejoVh2tCzC6mNzXFHY1ed+CVlDOfWmmTiDxIRvDXa+9bbogme4LQhK1rmrR
vb4Iqh+P6raQ87pG0RSrq6IUS2aykAS9n6tkU9ZR7xlXYM1CR94bzXUHPyz6TDs65+PVaYM9azPS
oep5EKnFzOVCAhP/ZuZWMDDi8hLcOZLyUrSjRDtr/t/XYW7DARFKa0PX06njcvhZwfyBhHHO2V90
jVyP4LMWuFFGau7yxC/zoRbAo6PYIwu9yWMnB56ynXP0o2KJZn9RaPss9pBpnQSgKXcaA9+uTOiw
Hg/sJThnAjAX3vx5LOIx43PrqEP0lrWLB8tm07N69L09x6OmSpoZNclfCy2euGk2dVjUZKvunPEL
wy6Q4jJoc0T2vIWda94xkDwx3qeBuTpWiPAKCPAPSETHEKNcRobFelhvUeWUFIqjKrhKr86Qwfbm
An/58W634Ya4QE/D4p7fwqMLjZM/kpJZVjXVoOGM4citUqQjcfP6NThKLoNkt0V3aZXEwxM48UJd
nnM8rmmqbk83PX7hoSxZB/MuIYtVg2hQx0z9931q6zOdO2r7TzdjA22PHd9Q6u+YDuDyJh0Wnv4e
+0C16rhKxN/8ZjrVTzFve+6Yjy5F61iF9Ji8AJxVZxBLSdEHxY3CI6FoXkM9gz6Fuvr7yptCICwN
cZAx3TSlnmpiUydW49vH4iT1w15hZocvSFydjsLk4v85ThnZiNDLaPSRktNHmmqs/YMJXP9TZ1Tf
NGMIRj/1Jixn6qSzizbOyx7/K8OSTv9CeK4njkaEqzD/uWipVoLdIX/6jjPzU8mu00gzvrLoggC2
LcY8qgwX42QwJ/SoGk/MppO1d4F5xQdlJRgf4Hb2UlsbGryhdnVu8jUS7TyGV/7wOVF92cbvBj9g
NLWPZLAw91zhFzsvWCUVmNUTA6Ze8GxQvUv/fQXdxFcCwBJr8ILhrWvy/HVLjbBncsBeCD34xOwx
HbDnL/rE5RMNIW7jqZlFYS7wgP4xn6wynJ91B5VDduFq4imHdJHoUv59j7pimUU7HH/jWQjVGpxe
fdPDl+yMkNktT4XZWgr3JrChQIm2DIRdRuf8257xy0R8F1YzKJlb79TKgEGOeVrwpIsnyLndl5aa
wM7w3OTQ50FsU++1Iq37YL4WQUnx9HZnMAr2mW8W4FbbHotkQJC3yPPhPGwcetRCKzDMVQKlR6Ck
hRRz3+3YVIDW4RCCKai90PdHWnlQJ03H90LFaCZ83HhukKiwe9wYM4OV2SN6r74h7zNLOWathr6S
H2+alZACAQNsoPLLEEnd7B0HOtBEVZliE0jbQb4QEfBP4IhC8Jw5PwPq+LkTalETpVgs5Qz20/zx
T3sUGcjaW2VAXxTc4lw0T7Jyhz9//Obh1uBLH42r2Ab/fwzdaRGGn050gbMkuN776pC9Ioy5M6Wb
tmA7MV4o6In4BJLcTui0PZzxJWQiZUrSmKOA/HI455S68BseJbXdMHaEYBzB6Xbo3x+vzdeztb0l
XCYFvUFN3dKJf4++27tnPuNGYGxMGzYFwR9VKCiVPrR/5VmYxKtzs+R/osDfVJf2Sk8LKrWZAcNS
w+Zsl3MxLHPczu7luznuDixHNAeVE/aR3Sz+9SuTXKo4o4XZ7wGKPwQt0k5ZeYRNKqRKCpg0DFMX
mCVqvnmKxgqFuJK4hnBmU4YYu0nHemd7u1VxubC8z31hWssupxpbehywcqdRGpnkPQF7cnntCgIC
zAibnTuggnBIM7V78ByOkGKJnaDvlBG1OpTUJQnwNH8hTWyu8rqB50n8V6tnrWaH415YAWt+bMHG
IMO2q9Z2R7gZbTnI1fxsXlycZmRgt0P/JDvbRtZCvmWaS5mysZ2Jl9f7vLEKeLV3qwnmf+YtwQux
Yq+gvXt4QeuWVyCt5lrU8UoYyoQMSy+DcJRLr1FMatV9q5q48r34pOL6sxnIV7aWlZxEckws5J4b
CPFeIL4UAtjWlkHY/H1LJeiBQGivT9lhiN/87QHIZ8vpu/0QVHADSMxshruXWBZvzsst64dZjjAS
nRHNYxSiNpIvsz25sdh7fdLFxJX8J7Bh/9s0lf2eh9foVNbSa3tthy9ZYGcHsnx1gva31vIvI7ze
QUgOpok4teWh/To4FElGrdNaA4U3QRnNuST5ylqNBBFDpbRsyBvlVzKVpnI+4xMz4rSQsp+X6ntj
25lLryeqPiwmTSHXofQui8qbJP60vApI+2DjKD+JhM4HD6SUTGJZX+WPb+wjmSf6u/irWN4pRJHb
rIyBIGLY3hPRI9Qlx/v1HaN+LChGHs4M9wCh8U7tV5kj3p8rGDbxpzJtUMS5TPPUfUYHyaCcdzjl
yFWZcLbCvA5UpWvz5QarRYuDlrAqI3e7OT9l5OHkf12SxpWAxb8YODAuJPcYvXSc39DgcA+ytifa
Z9gUfhAu1eTPUDpMlQ+pvbedeojkagFBbCBcJrzh51sYMCNVjKXYHfxP6S/6XuOP+5aryz7TU0kC
XvRfO+JBfZOSTFTtDjjlUZ65cjY+CudqXaG7AM+oFRaAnCwzzIJEqbaQkRGPXKd+ep7nix/XwdRG
E9DWbByuIIb7ZMRalNcukdaUlOrE3BEbvwxiwkyRuce6vIS1bbzMYrhUUIu8RV3UWQfCH4Q2NA9h
oH0LIFijGUBiDejOd/W1NMNuFCyxGo7+FYz/s3QxY8WcvA8TEI8KnZPWZV8Cbnb0aI3SShUXajTx
Yyc4QNHt1LDiCHf8GhOBMFhhC0XgBmDvfx70ImBJnOHCw/wS8m1Fg2gYRXGu2wbRPyesfOB2ui1u
XrKU+2Rp/YMLcE1XXhcLIK3auhyAq71F1+L4PE4Z+2KuNArvo8608Re+1C9wDxSTT6cJ3OD95C22
abEabrt19bAZIEfcvMcN9vd/oSDJTTD4nQKszsaEzJTUanVDta6pE0mYJwqR6EQ9emJAo5P5J2cD
zv/6VeBtkTXg2r4limaEUD/6qSqn41DTgwt9/C42G9symrHi1M0jnLFbuJQQ4K1PNfSdGIzx8koF
qv/qKFxduLcyJfmt65HdOpEmVJb+/M+FjDL+hksp69AD61dma13iwVw4U2Xssgx/OmIIyUdvNTdt
g6W9tPmpRs0et5w24eaxXWWX3x898yFPT1nwntvxmndwsPysm88MZivUlRsq2wfkuAqWunMWWHNw
QoRT1RnG/TAF6zZu2flKUjS8GZZm/U3BxAFxSd/RraeBu17xAiVuqJzmfizyOyrXRuH+GVRkHFyU
Grw2qYt6z0j/9/aCl9o1eC6QtH2b6YUrn+RK6u52GTlWVfseKcHNwoKW/zH3vE1GvZjzvgJNBDWy
1hiLH63bhf9mTfR2mSGOFNntFYF2cid0e9JjnPgOrj6KdiZnGN5zH+qBEqJ9MicKwchU57VI9P4e
PiVeWzHbFg6hPVvbysIDVjQklGInX70xzC6rFwnrDSJlICm4gNCz+HO7+z0/Ej60hPw9wjny8N29
SVLf3kufVuqrV4+ldIlhwsoFJ4AISklf/7vhaRWIDXbVnZNiE1BI2+D68NGAp5qWzNz4P/Ak0xJb
i630BkVqLPAhLfclA6jcCRo03ZK9CeKCROmYRp4XFYN7Xy4Mi58VEQXfIHTMDm1YhLKvgBDBZFQ1
WPPppT/fnX6wJKolQr0h3fcv7QIvy0LqO5OFKC1YGrmSK9nJsv9i0B92LjnGxyxyHaCRP6BKlGvO
P5Oydrv9t5VefnhW+84ykK6F+kc7ax59vc6Bu8g0b/lPW5uP9yc18PJ0mff81QmF4QLdBVpUzSSD
PswwlELgigHtdb5jvMp5FqLVT4/rRQdkHD/YfpItIm5hfkLLHPAE/XBniuI5oMDtP6YJobF+yc9e
MM+G7pwf2E2cTR8JWee0K0RCp3WspxbLZc/Anu/3PXpsxi5MxFcF3cueAkYfTVjX7CoIgQ3jNEHf
FeYDJB6JJh4W5hGS8FjNcDKLYKy2Yej0XXmjrMUtUb1zej17D9II9v6/BDcAtAx5CyzgceBW+rGW
1cu2f5rK/blwl69/kEliNGG/dQzAPIkLmVkn5ySh0FgaNUzZtTSBl1IxuixN1pWfLePU41oXBC4B
nQU3q9AaDJT+R5aOtrHjOhXwYx/EvoWURPC3jm5bO8/87q/qfebmvLufdE8DdakFrrpnmzubnTzm
ERg1mrDQUAmteIqLIV0oRYDnnRC9HuMuSmHimxrfNItqwLUOKWKEYrAJThtX2s78Ed/4pJe+4cPy
h+rKTTDfTRRkC6IzUL2WPHPXVNCNzy55DlGVbQiRJJOZfHeZRvkr4Qzo3G5gIu7akRcUv+afxsX1
GKSPtuHhXQPOBbRtPMSUNopmNgH5E5yPzo6jJhotL+/dRBZJtW6D8zWVuXcIOqaaw5YqTlnP5b9R
hJYbkpHt9WklVOc11FIp/VtQGLRHTAvw3kG23S1UCWYxOByzwj8PYIv3btjkO2TXiiBcFhMhvFe+
68m2JsCTWcz8/+tawz1afTrV0lrUFs2bxU+c3oYdowEDuO6V094yVHiG9Rmcij3x9av/np/y1stU
gAygA9YLqRAlTaxzenbYsaJePePGI7nauC18rFC0I5TTzcS+OBTBBchK9A0c9/WYqBKlvybp3VBf
x0j8UA6zlQyiCVNVIxM08C7sIPd0Xb7Garn+AKeihUi/IEHi1b+/JOR175UccZHmElpUiGQN62dr
SSELIdrrKUSJuJ8V5sJUAegtaVNar5BbMlCm0JwJfiDGpNvPLO2C66bIch12Y1K1KdmngSEc7StF
AhmUFMFQyrYTnH86DXlTT0+fLFu+XuXIcGlTfmcg3BWJ/iE01QCCJUXRWJTolODnplOWCpnl/v2g
a1nkGE3eHKw4K3NV5pJkHlAIk2uZOD96cEqJSoNJ/XGgxkEvP66ChJx492MCf3+jhgYTA+SUr+Px
z4NAYwKpNpa8WwhiLKoNWlYryufF8ACT2GHpUnt+tCgLU3gyQCRnVpZ+gkypd1XJGgmGnmSgogAX
9QyYncymbyu0F8QOTkW+joSZiejWE+5XpA7hePcA3Qe4hiODKKdarcCFIcyNtYfnsiX/XOzajZs9
/dwOmU2AoWPlSUfhF2zKQDYLIAUNkc4TkmcDBLQqXpo4fwyLA3OlllchyYMiUjSx53eWKxCVYt/O
h1PtldFARAFYDInjVZmz0m4hS09IR5td3G9Pea19ozKoqO+PQ6LUSXL3D5xKAfOpws+soWEJupG6
uW1Cbdkjlhcq64A15kagnFmUloEWO8h3pMNiPn2rTH8DA32/hskz8K6l3wsA2revBaQKhEk+8BFX
HW1ZGb3zT5ODpKseZzVD+PKHU8ke/AfwP+74g+DBUxFSGZZk2KDxxcACM1GqM/yXQ37EX+opK8I2
IvXy7uJK/dxZwnvrP09mmAwTAD+N8ukaeex90tBOwsK9Rxze+YsPR9rh9gzmVAZYE+PG+PuJv66b
3NTWVgOzt7MqWOo5IpGvvin9uwGNrZRMv82LKJn0MwUaClXe5WsdPuj0kdTUszSrXpt/d4ipi7t1
5B937KGLf5dW5N43YRt5coBjs753uXlKzxusJwNeksfIYqk7ufI6SBGazDvGhp/MKgjVb4k3KEjO
b5lpRFZkqp/b3h1GactInaO9a7SEKOgTNfLihkqa9TavVVU7F38D50zgQkoZ10lgd7NwpornFNen
6csraPd+MDlG+I8pCVlSDZ9axBkYaGV8VG2wBRQBZZeINKoLJuor08GeZ3Te9yZgGl3Tf1vZha3+
37NjH6V4zaMtRz7cM837EOA4wCjCEqqspdny2wifldadfCv8xY2wORi1IBoVJmyAoaa7OSjeSR0C
LZQ4mHcJ69q/ww3JraZiOmu/7Jik8Vuq/Hqdsr5w0PIkCJr2xBEh6pCy61192skzIHNovX23vzAT
kBUMO/dfi+I1p1qy7J9dbzHoAxDflOWT9Ql8sL38p45sYln4loaAavLr3JJY4JzahTYi2Z0ZDGpV
m6qAYQdJljhP9JDOs9FkIAYbU72P7VHN7HYnwUQZViyqE9sShutdHUPc0EZX3lMTH8w9f2ymCtM9
y998aX+6io3r3YllP1IAxMh5C77cg8cPozgKFTG0v+eBhDp4uAhmT1TvVyyNNN7Ul4P0lyUEPmRY
4rVjmNIKRtv7WWNtk+vaIYTKk740nOHH7u7mntDlsnHaqsKeJcBVpCKL/6bqa4w3Kc+Q9x73pAqz
ibbLybeqt+id7xfMBkJbcoEYXe2H58s1Y0DofwKAj3f78q3hkuJOBXakRS6uRAtRGNl52XZbCjA+
ITIR2pl3H1GlZcRQxPZBsZgkUygu9ChgFWJCK5xJTos8+eoMuDx5Hd8k/HjmxSusvN8nGX8Prflg
ZtqcxUuVnm9kH/ugn8A9l8+fonCVrnCCEsSCRs5IS5dw1VYHvWx2//B/83KewZOqsckRRzS7DjTN
88AW1PWfjRVpkNJg2w/mVr8ytPOol7lSBUu8/QCBtDUzP7I9Z7oek+d1j1nXBvsHRySjNmqrw7C7
Ksl1Tg9ZzD7Q9c53NzXXcWeGDxtZUDThwj+JhDjGNBpSNEQ3fW54RSHkN+QqR4wL6lDdkVoO4isr
5M+cCOC4iIRVh6+89esp4EW5TjVvHfWDthBV7+bqmc2J0kXsg6qzMoRuyU5t3+imsqz9E3zf8dwB
Z1uJ+ielyCrwezwA3X00K2uqBFMCGFZenWhn5U/xpFudKUPTYk1kJmx/G7rXBXwobOa4C5boKVY9
B0g1UJs1OZsCbp+jTr7JoTOrLi5XIii1+bub6WRV9er+WkgdPcj8a8hAKL+hNUi9ztBI9CrhBtaT
RQYyrYDeO7sueNOBav4gXstFZ3daicUOtjzB5m/w7fW/KlpkrnWbyg2sRGJSGtkrbVlUlK0IKph/
IATHjUBmaR5NH/SStQNtcPXgIFLSb8B30UAOSmHeV80AI8CiWzwCAXqer0doTJL44K5x5Erw2vlB
xDc3gkL0oDNtmbqFK5mYF/zJCt5rqcO0YMuOMkOxg+9wVreggB2Wdt6fKnJjYdRiymocdl90yB6m
0eEc76qMD3x3BuA6hzu99KB9wpxne32QLwHMtUX9Jg2r/w0Q6wn+CahZy9AKo8OJC2Ml9PLBC7KO
4G2qdUVvJBYMSHryW2RZMQpP6oj8zZC/XoRFPs9BHhWESWDx3PvpHOKzEmenoRRN1AO9vMW32gnt
FFkkrpq/l4rFZzwl/G7FnxJEyOxF3W2oV89VGHdJ4VH8SiDPKZnpvZys1xvCPxe78oscrAsm1BxK
nfX0TnoDkgim55sJ+vHt84lae/a6IJIrhIj9za/cNL69fcw+CDLX1sWG7dLbNwN9vxwnnEAUkyYd
uvgtp2JvesqPDusHGrHy9XH7KzhBoR6pBAUhHfw/G/7CxOwzpHyN+pMlKH8VIXnqJ9OTi2Crsj+K
Nadml6PF52JqqGlqz4K4ZFn99FI+amfGh0VjyXEPgZKZ8ZxRfwm96zAAVoTOq001nHUZQXQelcJM
fgA8aK5nccS0H6hDUemaHrPcGET6INpQNgLmcZqXJFG1/ixi79GfekIJB1t8Z3Qxt8HP4id4aGDj
6jPzTdI6U99fcT3dpJ78grnSb0ita9qNTLG7wWkFiFaGLgID3iJiK+LetXyGtFzNmAcdXj6mzMoR
uIChAg+u6zYJzuU8bNxQEio23O2J4k7vQQl0ehLrIQXC3LJo7FLX1uUIT7dIEU6Z401/hFTIP6/j
SCZQ2bz1zdIz9gnlWutr/hwSquQqx2bY3Q6TWuJ/7h2+d1dv10nHR84zwawqACeK8YQcRWQ3AOgG
DAdgqVf7DOWdWm0oHcIT23a/6wKrSbLrAC99OMlyK2NVdQLQg/80DK2tES7K0/XdzqocVqA/8oUu
kwcP2iAk8PG4vAerv9mdAmW0LdNRq8epGd7N1uS7n5rubTvXZaLphifS9V2w7fWUeXp9zW2LBmO6
8qanzzjVvuaTeVz4gS8D4YGZ6IYV28QzPSsMhBdXPOeFqSoxkSnAi0R427PDzCB6SY0FXoxW6YbE
7JpR+MKCiy+IW10JAkHAjMfC1vGhEVNcsMsLgDoajGxh3pugeVQLGzvPrcDi+n9gOhudTJ6GOiZV
jNLydc/+mfiigDHnP7SfsUocSPQU2VsV73R5LrRkZ4Rbr28MSyLrsISuQ58P5MzE5LBFxU7OJrEQ
enJMog+9+d4nw9xzCPoP9J8orgvjXg7WvE3qNnLnY2wOgXYcGJFxyo/a/FP3FeFYCML2UMlAKOn6
cb0v6i+WjxxpcOjeGJ3lEh991su+94qXyvEtKkZJuwHSVnSkZ6rTtOLYSNwWExAmS4AkTSjVf/pd
loW4bUvXv8RAYc0U79TawSfQwxQ38wGdlBIgB9bQFMehY+js2b06Mq0+aYZarotuk5lxIR5Ke8LZ
0Pv6uXMRcZNzWxLEAdsvPKGiYSn7gMhjP1HZ/VVnXGlNnMLCQKEncH/kpJi6ahPQLWHNM1q9OpeI
ysLi8mQG28iWfvYGOl6aNCZFSBeKCnvpAWoE220fY9i1eHsjMLvC8TIzhZKLfxrfE+AvxkJpZPVz
7yYKOXJzSWTGfHC90wR36tkvz1IOXrXJtHP3hZbNMDEWhPcvfROxScF6rnK1k8guCrS9DmLqKShM
cho6SxAfEi/xpisrbECr+xEdFuW3FhMxCEDE3m5WM/xNoliQudNdgFSdB+u3Ou5cSAvbga4ONGDj
OGd3TkepwjY+nCFjpqU3322hZXjI78SmqcG4kRQUKTbZLcLOPqqj7V7sq9hTqtmVK4UgWKYsXr/Y
Rspy0HK7qzej3g1rMSM6ksPDpg7NkOiriPnhDLRWgHJarp7jlc+4j3+rnf3p8a9tecTahip3zTbE
ZBXz8ninSHnl4G3ti3UJ/kISDRrEUWhya4ihc8kt5Yx3aUw56ze1KUbOvxEqX54WHUC+xog2vvqq
RqefT/NxJcqEodAvXrC4VGpPnqVGo0TYGoIlOqE/Zoo1u81cciC39poYOMK2dPUH88dmslcckWP7
O41HtF2CggSYwJi7wgjeA73S6lBRZwup3IGXhux8xdUs23nX5vpHm6ml0gE+fbZuuxdRvY9Q0/i+
uHqlwnVNoNkJ1OQ+r3rKlDe+wn3xefhAoCVhaU2IeVLR5WwC4hGjeWBi7IbAKPk4AXE8dHxb4BP3
i7jNtOM0MmozZKi/mDKn38wOh6k9KYe58Flj0+4z6KAr4+ZyMCBW0srobQYBpEPaStrh6UvdA43Z
IK5WQLZ/OpKwZgnLQG/D9zwYHCJNnfucGHV+w/SUt/WLC0RgzFzCiQWcHaVgyYHu/0KO59YRuL34
uxOpxowml9cFDjHR0/Ltueo0nLrlOJO6l5vd4cUJI+UKd4mnNX7yKuKhIuNzqSy3RYqU81EyV7Pr
8Sm2G1XV+p4BuxWKYt+d2piqPNQZqktfAYnqu/xAp5E1PHQ44WaL4UBVehClKkWaPU86NO0VYWVt
0xSJixLjBBDJIFn6Oj8SJGbvw5LQ0Aqv4kyfdIZzMqjlMBpfySvvpA4s4Qnu82oIJsrMIcz/SvMy
r0dP0ujCzAZ50mDeNh4c6n5nut/r7q7R4/LaAQFWwrRSaC6b//+riqF/fajE03Mlq+HSx5UJcqkN
8EgG+LkaSykJ3YbGhr478mN9BG42XR1TyPVEp5lYJIvbiq1xIaGBsVmY7fJwcDbn6b57zd1KkGzC
bvdBa21EIxwSEl+5ySxtMGnetBkxQ5/woLlo/sun/rGfwS2R4n07lU5nvMEfoBxThLmYqojLkmug
/ewML3YqxU6r5cYt27rkjKH6PtmgxUhoRmD7FwtgPvPggfAm9wp9Nq0kAqQNPxHRnXHdU68QGv1Y
Ag1ey2MG5VT777So9e5RZfIbBhR1UmMs+yPZoKqsJ9+Msv/R5Xk+myukpHS6dBk2mRNs96EepNdn
3sKu66JXkFLkIjvZHoEfOWElzZrrdBOuTt9uCZFu/OunnWrOl4OfSt0gIl/U6zolYIGEePKIALcc
R2JLmdjAprQ0Ujj/XekzAdgXDECdMRIH7Sbv5bdBkcimU4Jx47fJvkKsqiy+/5Sgo2ad434UO57+
7Mfu8dCzktaEYEi9m4YZdleek8pDdjflYLRzcy91M0bHdhmquQnu4YHY3zmw9mTSIxX4E8dxsMc1
uMaGl77R0o0+/fb0JAoNjLrngrPnFN3AX9P7SESYAw+4sY9IL5cDB2wltLSmhkPCPK9aVptugqg2
Chdn4dV4LL1z0ANJmgnjeYr0PVI7ECt7HO1Kb/I7rOpEprFP86qEDPNtn512ORLwbu09rLuzvGc6
z7hu6EYJ9dLMOoFNkpKxIsoymsxKaQqV3HpjMplek/yF0g4obAPaLUpCFY1S3yeDZ6K/Z57p7cLu
UQpI9rg90WDu31wlrmDQZGXgD819AF6V06dFeP3sHeqPsm4G+qdT85Zn8VQq7OJFaH5Lvj9iWY0L
Zj1Z87Eld7ypuMnJaOaxs14q9d0A2f8AaEhqtTF+8rrsh0d7NU8XX/5n0EFe60WS8gnHC41jtRKZ
gD0sZ722eEM5NJpXI/1S+V335LXZV1rbsiV6QQPj7gnnhKQzo6MI39TDDF55NkWe8j1TpNL9MxOO
lkr5FUhcsbutn6CSqb7Y5t7v0AgHfXDOXc2yr2DSQAoqdv+5wiOju/dcAvNo4jWsfUR1wltN7Z/4
g3XQxjTA+r2YCLyrKWCcXbbh+ykdnHmegbAKynSl3+OyFNl9oBY/bkzCXHizKyUWOITbv2zAFome
dHStdJca7vgmFmfTcq8ylwCrnysoVa6IXgGC27UcYP6KCTBotZddMxfGsjrlWXnfCCiovBHnGIly
o3yMihjpX6IDmlkElIhlK5IdqXQhkTtlR9W8d5jE+IqdeU0iJ301w5DQc1H1sTPRN3eUWO3Y5y0g
x9GFaH6AihmsWh9JraFrxBSI1dkojXkKLP9MbSvLnMsYXzprgr/mGGH2o/+MQENtT6I6YkKw3TC6
oNj4c3Bwf5cJVM2yMK17Qk8HKsaIsaOA84N40qVmo01oRnDvhfWGUuG91uroD1Si0T2AioVcdvHM
/gLte7ojnQSstoEfwaZ5w/qGITOKljRae9fIT84BriGsf2azIo6YSRYF11zhje9JWVddSBUXd5iu
Qzjk5c85SYuNbcujC/niVboBJNs/oTuqA+8pArlRJDR8dnVePIf/f53bmsZB+M0zpa/E2kgrA5Sy
ipiC3eJGDDS5RPBZDd/g+BFzC1U7aulyLTgagGxpEtRn6khnSXbHh1U0xfoqpzC0PoaDpDsTZi+b
/pYxazIK371tSbY/nvdWqx+AZG4vl/2ZsV8HO85mcRo7ULUr3QeHlNoXpqLoX8y1xsM48ISbnVxj
tCzmoKf2oPQ0l0qPcSV9YfZVZKnOlCDXYnRoUdBfk9D9sNAwqn2/TiR0c7lIWUIasIcg2bYGVH2Z
iC/1vI9GlLYT3MvK19nX8DQt/SprA5ucykdToQ5Jc6JHVt3aI4hu5BGncKsVLChPExPF3lTVx6+h
vGwFoOQbKmCsuBEKSp89z51I1Yu45cTY4pSgYRvHzhkQ1l4gGWl7byZ8O360kMXWovJhS6LtcVH0
MGULqnwnGll5eS+sAm2WX2eRkS+xljPLy9a7BhkjycVtErmHf/pKP+msd+FPJ2Ew7w183qxkchLf
FOgBHnz06nxndPwIlnDaJxEwclc2plRGf1xUSmFL0FHQ7CyMfY92hm1Sq9lVYr8rSwFHTv98oDqY
zbiVX6QDUhioeQoEPTvfi4ZNdGiKkr0dF/8ROb/PBwyDO6uPZxd6xJ8K2qhQLWhw0trqLbnz2FyW
A9mMUZ+yjyQ2Cu1OwEjcmD+sihP7sm4wGR/6Imm6htz9wEJ0ZPGugef4QAwWdWXWu4B7niDpxG3o
B2n9ne/t8xGU+TmjXQVwUQEqznnfLKLBkBo1RkKC4AhENPuHG34xJTJBIMCcYmvvdXLEJce7FkNj
uBwpKni8DCaHN+n9Rg7tzLcGngmgULdbPpJeTA8OpjWFoGsKslGUD/wxebI803XdrfS6mWIt7wES
fSz8nzqU71x/kgYgfhu8NS6Aratiw3SK9hYrv3K2OW+lmKpUpSgJnwjiRBVwn2+sJhCM+IzH9gAJ
oduo6ci1CPvVdZqReTBRPftHIk3gGR0gg5kB5FIXtzLFJQWT0OkaY6mrt9aN3TFoZv0LPIiH8xmb
YGwKLN8MsObqiPiwO6rETUYCFeZ4QYP9htgxBHev+JlBZ6Jn4l9nLx4b/tWSRJH0zq9Qg7YINrS2
q2hErq3LvZfXN4a24qd8zK/jG5epDRitBc8ib3ZhWpjoKYI0fLUZQI79a6JcCYAkSn9HxZq51nhs
gj2eeqyN7EWHTKvDUBA+1TnFeoktakbOo1HN9zsT5YItG/SUgSGgWMprYcPtOrrbvJBuADvp5XW2
1ROv4AFFIP31HZVsZHqfzZYwdga5M1BD6gwmnTkFQXsx5C/6jmQ4kd+QE1WBpf+7D4CjTrU/BX0H
GOSOxOowek7BeRV0JCtHiQwpQE7Rkft3vanxRjbjKvoXS66JjpmGc7S2XllX/xtbB7rJ0gCRQpOc
07z7/zD6XqQb6sG7TecV5lfPip/cjWx0ErmW6BCYSvfyC+mS33CLabDg8kHwPHN2Uhf/cHHjoujr
K6YXuIcf6wZhYKTDOQ0R+LHzCrBm9Akt5Z+loxsW/WrKi7t7YNY5EjNUTneh3D3n/n8XLSWiyBOu
v3NHNFtPEuNGXeKDIWVvApSB/EI3N7ZzhTSjuzU6AnZiskM+FO4Zjvj2q3fnR/IApTvnxIiGnxgX
GqB4+nUcryZuH7nZZW/b6WEz3dokxcgommCqLj2VPjXn7d8NzfHwxC7dfUjkIZKYLHT51T/rT//T
N9CI5Xys2tc92+5bn++JDMlVo9Ov01SM7NVRTQulFh+h/EjApkXswPs1JaUYdfb5WdWF5Bauz2Y9
KwXX948a9f4wShJtjZ7MZWNS23Oh0A9xUm5XjZbUrpeGiZb+UoMq7Up7r9BXDhnNwWan8cNZyWFR
5vokdrTD1A6i3v3ahIVJQJfdAL/Fvj5RQy3Ynz8jQcS+dmm0vS7HbYmbXU9IAJCzIbdgNBLowhDK
+bDcI0m7s922V1/VqROEyUT40wPsdv9aUQYrNY5/os2pq1wuSr6vK0bvafExfzz8ZxlHWKGr2OVT
pwlt4XCorrVy9M1+fv00N/eOEvxHF6X2chJ9/AreIUaUGuYLb7VDBPwJXiXe1zyVQGtlf36/Suds
HNxz6ecLcWry+GbzYqSvyTZqcpnUCTlc513cYpGDUTX90UDQWnQyZZxOLEm5D5ks+g+yrOuMZG8v
K6OcnRBiXnYbs6YYmxq+/AxU+iyevYVGRwK8ELWKENoHAHGZw+0OQU3gm1gJmxSXaj1aeCBQrfd1
K3nmaZeZBijziy9WmpTyqW/rlwlKIYuqQpB+BUGJuhS1BJ9LOChCgE247dwyVFzqhR6ptj1ebYId
w9bUo2cbVSwJoRn1mGKIZ053j9Wa0DlyP4MCRqpNbBSQnuikzveKeVllgTTXcn4AxfORcieg+w42
8JhBILhaOL53MdLiWzHzAEcY/TT1T/UFBHOvra+KP0QdWzNHC4PSHqPKKGSfhvxI6jc4pEoq6RyM
KUActoXbAPT4c2ghQZZzobsWQ3uFT/Wyb7RSzMb1CwSK/pX6KQQkaO4N9BojvcC30dZ17UB92vHg
jS9rxkfKNiy7U6ekBRMPY2bsCu9cFOxMHFGlxODqujRjSrsSvE9md/nq+5B78AX5HzvT1TdTuerY
dzCTljaDw6SDoTJAvFsv5UFnGvV185LJeYgs9xL9DsesqCQVaAAbqYOzbZwfrUzXFwVhpNOJDbTW
8OO0+nf1KXjfsCmpmrcA687fN0cAGwoTG05z2ZuYXwliAUcRwLijYTpviFE8ZXvI65lvN2qydK+S
uY+G4zQlHDm6MfO79cQM+M03gpi5onMIlhThyKC0W+UnP8dRZVauOa2BJvwDs2k6kC0DRf1CwdAS
urRy7FFxJUbTnR9Q7vWG3lLcJrUbJ9tFb+dQmVSlS+u1O7IJfP/VXvchaC9oPyFcs/aN2Zuzg3+c
ja/WmJFNuEddMWqUWCkvfb8CxKQpx5QbjYr1NljqUcugaRWzwcfsAyFs3+FqgGN/QGkN1VU52mee
ZHwzcuUiaMBwuXIVHR1l3LXhZmZjB0vismzaAbg86N+knoCZQ+CHCrzi+EVZHQdIOkGTWLUD6WjF
w0ugzroM3p4TizqjIfCEoxi9681scBWegikJjfXvqHeLlH3W2TfSwQIY2T1aCGgdm3GhLD/uVsr5
SmAfo6sAuHa4PqQqRwUvPzb+aj0XGrdDtLnJ3bt3uUEOMOYUUhS//Qk6yR8dtHPqHjBGh4mDo1Z7
oD34HDtCF+dJPm9K6fmuEUbXza+npyuqxD+erW97g1a1/5QwNQzKmnea4ErOOjDxUl+legKZVONp
iuyE3rf57T8TyOpYSh8v6ereSRWQao2ctXSpskcFpy4gEUyPatpO1Qs+h+XVJAOAPTJTyVzlAY7X
ycp6AJ6+RP8ub1wRJSmDjo4Mq/2QayP2XbynYH/K2+Rg1vZ7pSF32KxLEVnQb9VjNlHJBCEu+w8V
bCJ80gc3e6VbYwHcUsDyeCdkOyfWzWScymfJKU7LJTs2Z2vBuwU3NLBTQYv2c/Sk3kCz9jIN7ue2
j0SvTIwFJSxWwdDThxJpIZeowkNVZbcjPWiHvigRnpTzJlEDAWLE0IsW6M0fTWIr4hODzBCJJFnN
6opwFf8hgfh2g6gNn3DPPEkLmUh4rTyNZwR5jN2LhcWR3Ouz+tI7IWTVEmUR+P9z21blJhXAqxSI
HSbOBfJAhdeFrq4ixU/sBxNKN98BANuKdEzviHc0g2joizQka7WBQifxC0UXpISNoVLBR260v+AA
2TG8eOD0U3SYxStlki689DkI6ijz3D9Osd3P+6o+RFrQy/UMszX1bVuyAKx8MD8uzRQfwcxglEtb
zNEy1rIQ1pQbvAoHGObaZEdaEx/zn+5hBoDgWpnO41B2CzFmD90OQzLuyH6yfvoeVn0Qrq3fbrJL
XxMdrKW3uxkiva2wCCNM+8xAAAC9snnDSfi+Dal8c3XaABqroXILGBY86J6RWRU9mQ9dq20rnG6o
zDFIpj2XIkElPgcMk2Xe+DgSTwfcpZEIl8Q/U7WDgw8bZ0vCdaFHt5RACZO/6Wg28Lz5r2mpsXui
dMKjCFah+HQrUik+kQEz0JxCpSjYZxUakE0Xa6os/uqirvE42wUtA9gb8CguRgmYhNe+tdlked7T
i78XO+S6mjcb48XL5yNknhdjlB7SHPNsDXOBeMaZNdcYqCMIUSvSVrqNInYyasytUQsNiKLnucuM
R9euqQCCrL2FcxbA+ExpoNSvyi5x+7ycRXq2cav2DyuaIU7qY2/lTrhjnrpOopaE4NGdd6pc1L8T
xLfjJxywtA+WWLyWjSqGmWqakk5SPhP6uwCN2ybcgSKkUNoEZgbw2SR1aKvsdPCI21U9/II8Sw0f
EYxNYcG1Yab+8YQe5Txm5Z6Mf800xjtO+Sj9jtLuQvUj8CSYZzyov4HDfwEkpRIi52CQ3XGG4QDV
5+BM4rEGikniZ6fXrPt1Lb1qogpGMhQJm70SZuk7Fcneek3UUfmt1XNDMd3MhhufKNAXcZDz1F5Q
Ie4JIUbU3bc757YRk3L5t2F/RvyFBq/Hcw/Sd0OnH6eK9kzVVqeyvcF5CwbUuCAXmgdy5MiWj70N
eEBb8wDwgRPPLpnzX7gpstQorYmcdQRRDLUqHGVFgW3SO5bnA2zkZZjyvodBg0CivIRcot37Li0+
2qX6AqpGXYKXV7W0x3VzhVw0heg5YUCpBS/8+8Rqc3YYVpd9Gzv44tdA7a3U0B1EREcfU1l4Q/rD
zU/gfDCNeliP+x5g7zy5oErHS532RbNBlw6rWDR5e1VOEtUzaPG6IgHqvesuod4XmZFgX4oaIkfS
uZgOC5iFbFeHTHXCvoRNTG4VUPnJiYjQKl86sWYcFuEDYrLBB62lDhJaFjdNxi9Ur5fPMSZLVhns
LBA2fnN1qhFdBWZnM07ECqmvLKR83zwQw9ZSFzg7JIssurgBIAuey6E2X8L/0uCsvTF3WqXHhuPK
50PNcrbZhrUNP27CiZLv/GlyHuTlMOq/3oWTCXvGc9IXIsQYXq6JPvV0uYyHsA6cGW0q8pHUhEFs
1KjaBuEmAmEvVWVV6gBaRxDICpVknUvW1pEM1ajaAzB7r65fTycEWH3oZuAsbKxSIWVIltCB0clw
SeezyQUBXkaYGrjE/+hEqmoI4P1+u7XatUzpKG8fa8lYjT2cIx9PY3P7Cugm5V+1cZ/5ZcmhBBhd
aXy9KBlHryutfdMBONMLR8+GIHfI8EluCI7kg3IswYunli7Ru7P9jeDdHmIqh+0TKLBpC8QXTJiz
PaZEul8Dtmh8Snd214tcI1BY9hV0Wms+WJdpNahalDKS9OnupkSWgU1+veduUCA8jukl/DmK+mae
iVYK/TWkzNhMEGisMYi7GMJrXNf5/r3Rufw0IArZfJOv43S98hTdkJKOehonQuzlq90hDz44yLm5
lLM4+BsHGSWsJQRauy8MHD/Jlg6wDmgKiZgCVB31TtRxpc1PFZUsAA1ZuwBGhmzFG/+jMQM3VQ/1
YE3fwUt1GJmJ818mlqpaby7VGFl+GoOP+D+xb2SLNFKOY5aLPLJs0PvaJZDZ/nn4DJBIHZCJuxD/
KTEW0uoTuisGdQQ1GGjrvoieTrE+8ztfdEt0L+j/9eUiF9y0xLbpTECt8iTMp3PP3FwHqVtRBqMP
+Xzxme20yVtuTJUTMh+JKbFKKRY35SHyN/q5IkHR0VLXjOKxuSYTSMmTYNOrfr/4tASQof36q4+Q
3ABEV7b7Zho3scAXMyaBxXlm8fYdO/+VM8qQh2xRuzBHw6e8sWoOIZUMp5q+t/xYQIfcq7D0wtfd
/54LvPLsgF1kBWkJpGwWffeweSqDpB80odJuaPdMq0vCeu3fSV7v2w/nIBMUR/Kti5K2wDTkA/HP
JMdqya6pKZyfKGYRX+i2KmtYjCo+IlNdfDr61G7BBZ61PXRIOUhHXvtziYHP4JZi5xlLDRIeIUAr
cV/hyzbjiVpBRusv+LGhVZ66rAMbHjNBTqyQUmEp0oQdYh/9Nv1/Bv4r+KEvavEKEs0TxRynXr3d
n2klv3s4MmemOV7xJT5wXWnEurk8pBXk7lgwzPxN//E2VgZqRf5QCMGNXw0NtqB3O9D+5adxAEmg
/lUqKXJGIb4+FyQW5fibWkUPrwxZVb/885UOuJLPmI3asijtqoe5wSd8QfPGgvFb9jJpZqStbx0v
kPCs7THVVwgUtBWIhgGnCOB7tlOGD2UDSMWo7g6vcbzxCg4UuQIDSL/UZxw1KXqNW8ZwfbQAE7Ps
7kHb2ozSLeBYzWIKdG01d4PDUJDkDiD7u+epsoqcmuY3AH9TPzXzBwZ8H9Ni3xxHz7zN6JpIymUF
voT2WKtLCRFJPwSgExVi/SY/SchVDdxTAa43zR5xseu9S9z3nI31hC16FUPtqoM7wkBB45MXI1CP
wk3357aJRSPa1UZhGqYGLChK15Pd+dRLe3ENTJo9UnWL2u9PK7O2MPKw8JnBOgTiqgwxYm/b8DE/
ITb8F9t+0krkxPN+Yay0drFR6Tv1Gq7bTJLwsUbndDynqZsaOTg3QKnV1hq9Z2PLPcgQduWFskTR
nIgHgSj8KKk46DaUwR80/4q8hOz7fcwHCzVtHlGE0nDnJQ29sLv2//KaKALA2lF92C9IVvsB2XRj
6aR7giZsiU1mhU2U4pWnteFwV56EegVPmjFUJOf0A1OzvKS1ZDPOWOMDYbbjO5PGPzUEQbhFEquj
+C0yZ+AneB9yhRsEV8AyJLpx+jtNgeSraSYRQKm6xQkcTjL9WW76Gl3GOTK/gnOfhqgu8m+3fBdv
YB7bUKh2gowT5qJaInk0POfKDUcpRGQwa3DxLlfZvD3hczBz0ZE88tqrXi19AXykOu06GDTU0obq
5HNni9zS2WipJy4SgpZG9vIv4rVIWnXzqZcc8GjVPqyoipliX3db+h1hsLjnju3FCufYoK/6cdeK
k95CskPXxUxXn1vp1qITEAPbmj6JhOrG1gifTwVeVKnveSJ8n63sxrVXMwgMFXwy0oo8wYRvJ2eD
jXr0LAJ21fcBjK7rcC4CiqJx98nson46dNFSWp8biaO/IskPJI5Tph/b7cT1CxDrv1IYqb+9dcaY
iwGdILqABk3PMHHYMt43R0UkMBrS7gpPOLxslEpVdrfiq+uoU8kuR6pKz7zennURFKhWaVEaekvz
+Elwi1G6g8jyv/0wYR/1WHdmLyW0K0GtKcGojwN6U+UhgcRZeKVYc4zfXhhfAZfHlpMjQjlrel6M
opCGxLAD3zwBezLmPFunrsTvui9UJfqa5PYTuVR8MV+Ck5uYgVvuUTebQaxtf5Fiir3mla0cD4Ps
ePyK5XE7tq+vKI2Ggt+Wz6JaqD4uex0Yd+XKCCQ02aPO3bdf7L0bS/bDjLK+w2fpO1Zli6B0i9Gs
mLS+GLbBp+LOVkFF/6qYG6Crm922dHvgBDCd7tHwwGfcsEumKgs/bsSLGyy+vhLZQB+k1/rH15Ho
/7+sB+0mB+ClhoubJ+bpR0VOArTT/rVerGomFmU8FQ/ESvcO83kCOXwlWxmSTARXpuCzkP5SIeXY
2e3Rq1YQtOWyXf9Xa1mxdXJksUOqBQFfSLz6HMfizuJ1FFsJt1jM9WF0VS5HYvTgNrLBsG+3sfhz
wirKBfs8P0oWX45wUwptbg1iXqIwL6yg2v9v3PTOT66gbRrO/3YNp/9J2yi55+HO3VCnoG7xrKif
PVZbS6zgMQUmiqqxNXUdnjmom5lcOPjvg222csSYCAEZGQijlsDZzSQ8WW86coypL5F37KI4mzs0
s+2c2ki8UtDzQdezYnusvlOOItgwc3ZW5jqTLo6oDBRbR9QwghP8Fc/7M3+nUFEIg5CwHJkFCpjo
TJcvlNATlWImvmJi+U/GU4LpVEYUm9Cj4P+7MhAuh9ZIIXC+SLdsNU3lCGHzk6y4vF4WQ0RrXlhE
URdLkfLQSel0QSWwC/ByvU32mkxq2WEWiB2PPD/FTLsp6Ir3xV5b3pv7SW/Ymcp7P8L3QW18gMsZ
VHpffAlka4bc6t/2vtALaqdUcnwI5E02FaYUoduDCZEepvd4zn9kPqNfnKGjO73i5oHdD6B8LDnj
CLj+VcxV51QBVOsXE0WfMclu5S2Vhh1swj+oQ3FSb+6btrL5738L26gpLqe3IF5uTHvge9J2ALuM
lzpc9iDvpCTnDVwztKksc+f207tRUG1gKyVtyhu7FXMbIQkpWDjWOCRel0NRQbSmFH+ENXlw52UU
l70VuaqS3T8qMJirSVh6D0lDSPU/u7MRbSP3ECm+9MBaQ8ez3YHvNKLvNme0r2+K/hwazleBbkSv
3SvYwwNVal7meIZ7TYIQvoSL/vfx+l4T0z2vlHZHiNl0P4ntZjGelRRtIFDTK8tOMpbdSoXmEIRn
xodjFUjAiIh0bM49l3cwATv83bRJYg93HRBM3uEaC0KspJcj87sGi27td7PoGb9TYe/6iAMTZhM8
4cVWy/4ayzWZXNYHoKrEnfGCQ2JqdVvSqI1qAcUpkRByxCDJTg5lc/t2K3EyrRk6j3NQdukXEIt1
mcl9x08+OFbjeR1MKpesp9eq07wr2BlYqB35tmUuYnrUg88DMgG+uys9dU0Kr/yTWBrpIIvo5RhO
GBy7jkZe+4OTZ6rWSTTR7X2DFk8eWSVIndVNqFkYandFPwti6WP37zo2Z9CXmwyqxfrZdFyjk8gl
Dj8Zg9SOh1aMs2wxdsDTKAzN0kCbdVdYIFTgi8VE8quwmhIBsVuxEjjtAvSjSa+XpiLb8tbeUZmL
AySmFXqi1Bcp1+WxfyL6Z15PM7DhddAShL2XtFBgZRqpWbg7hL+PWt8D19QMGVUXfZBKes1e6Fr9
+ZdnmVOXyuRFwvurXSAWZ9TOj3dKgw8ERdQRWWXi3lM2YJ/WXu+Zgjolwvj9C8nbVOdwguEnCrgo
7WpziTwM2aKaiuiw3Zs1amC6YXlqfayrPRlQyFhtQ3kEC5mDyIJjtJiDnO5OTEUJ7+ksm/L2mPCW
FqWGVKMsjW7kg4QGSyIelTo/U0M6/jRg+2g2icFxmmge2hKDbYCuLbOvnLeM3k0q3mOytbrBvkXU
0KgDoPMQdfAZCT0jfgwFoNmPt/fdiqXaGbn5vzJ3u82vJ/gJqjLFFQvXmL1AK5qrvn2RZptqLBx6
sfNTgtgpPHixVOtISM3B2bPdWnSzgf97esuPTiFKFZLyNMZP00c3Gf8Wm/OGd8+KLLbMPBxi87NU
D460zqdn8gsahyjT/2ssE+imRBEdEZV9lnFpuaenTNHQjSWfMCJrHaqu0SdCJcbqj+fQ74cv/6YM
d0VjxEfjjNAoP48yYdXRXB4ek87B5pZah2+h9jD9SVA65Zr5y3QK6EZcVtGL/DANbm3wWEylFAz6
F3zSdclFRs8ty+gZr94JAkHx2JlmbB2pcWa8NJTZ1j/bXWWcEJXcmd5XNdRNO5dNlHPMzi58quTM
LbaJCGOWR9j22+vEUDSRsEJ1iJOCs4dICapFhJBa7A3e9rGp2eke4o9HwdFR6YPn8R8BmIPsPcDC
1IuRz4aNCawSeY4UBQIQ0bSoMf1lbwKmILJCS6+BB5pBX9ddo82IDcZG3eqXX39RVOL1LYHUSe1q
Ks4syGPuInkuQ2A4/qB1/5bN80aH9Vlrdhr8bi/0XV/ZhDkOdvGYuj3tBf8jxtLB8KvWNPqSai76
GW6lmoRaHFAI6W2EJzxaRXbQj0DvAMk2lOLxLP8XhFa7fUN7TKB593zxz0INhA+ST46ZXXizDqS+
Z+/y3agPII2diEdimKH0OIR89aMF+8TnuZBwbUVImwLXtRLPOmhx0BtCUcFitUzr4NTXkjkZAtdo
I4lOWJ2RdBKOEUNvq9sXansuQiljzKcs6VLYm2BavHN5OY8FLOqpXEpXbfFcl7481XzdTibqj7lW
b6wF3gjxU8WwoV6NmP34+xkfr7PHpUW1Gl3Cy1I4vUWYBdsyXr+5RlMhu7eYgTLpyHR3A4qzlalU
jyVpRRsjM2PRIAl9hcuVB4HSWmFkdqBx329xgESOcV7yQ4KcykeyDjNejAtxPwy5khYE+rcBYtaA
Ourzcl19D4s2OBsbcojPJkhezQmfntzeT8He0pqTa/yAImBL8Kc2NtEegj343VflFw3Jtghl3gRi
yN44hR5PUDkRvnhAitYHL81O6N8b04yUR1hQ7d5mMl7ufHPBlcdrSchu1q/k+6w3WKSiN/VJPL+Y
F7mTzuPXqPe2cEB+WtVSfs5oxfJ7+IwAUSI76ryBWz4LKoS08iEM9/4JHjkyAXw1ObVUwIm+juF/
hBs3cL+vWGc+kLo2ysHXeZ2z3N4LJE9fljhyDorybFxd4h/IYubAUExvVOhW2bbBf28Vm8YiUHt6
RdtmUFb1Z5d7oI7TkjXxobrj9V7IyrRKRq5kWcZOsQ8nhHL7mXvVxLGj0Sw8+Dfata1bkgXR30EO
kW3RpeKY5A0svqqdKgprLr064ZN7tdqPuCOdnFWTcV8fwqURtECO7IAk76mzMimp34jsEXh3Fb2a
KpGNhxFcYwS/sp4/SVbFJ25RHfiuKHbxslIJRc0mH7CaComJAt//zQrEYLaZFmKmVss2J00eiwOk
+M4KwsMcz1FP4H0dUIoyOERiGYRHusFInt1mjIpqcaHDhjw1ujwJ66MfuAopCZCI5C6Ns5eJQDaM
bQWyqpgWUrO4tJFIpHqWG/lzBS2xMKPV5xTRKKxaGw2DvBwXdKfLsQaFAAgQwhN2iPtluNdX165U
vaWNmMwO5czYqh4KH1ZlhxZDZujSJPptsUAm1i+RdlowzXSn/Q1yvRm7FHmArT/o4vKDGW4iY8NF
YvTpkCeJ+ud8xcj9ClwHVDNx9vcucOKnnATHB4/wWjihkJ6bSTAmlGJFeTN3s738OQ0zK6lT/d3b
9BnfdUXshI9NEzpsMluccrHvWroWj6sgyq++sz4fqvEragAq2pZ0ZMlmNK3biDlcss7G89gv//eQ
GZAJyIJFHutDVOI/NKzEfJZkztywkcFM+bCwT9kzAjzmq5WwT0r1fOXyY6V/ahylKQEo2Td0LEe3
DNwCbnUX+6I0Et11vhvmGZ6fSft9/9C/ElcJI/X3lw3fwvFLu1WxCMgiUS27b6PLMvSSlogXsHOY
5stZ50go1VkZIimEiS+mXxo4kOq/rhLGM/4oiyMN9y23smcrK/b3bu9mdXxgK/TsGtWU+EZhy98k
eO9U9eUyYwmqEFV9aT5kjUCkyR7HcMnxSTT+e/szUpQUYWaEpbpIbpgp9blc8oPKPPgJ9HTOePcL
F0vcxHyYbj2n7A2k7j8mIa9yVesneX4R9rYCyEbQ9wX+NLkG/0NkuItuS92UUvbyyeYE7hyONhwD
cJLOaeAKEWhVIi3GLB3o2u5iyfba0PKPchYzQzcKkNIq/g26/DFHzPk0WH3srHkMAWZCg1lDsltm
+Q3fkWyjeg6xmbLJOFRgdFFLSSR103EExC8G5u1/S5NkGEbQdWdVEU6cHG1GlDWtqH7RA3x8HCjX
LoGIMjrxWdhLH6dYDtnIDTKDme6l+cyMr8puBruMmjtzscGmxBGeM9eRKDjRtIM3eGHiBdc8lpjY
VxsO8mVNRDksiwwXX7BmF/tXaMFqG6/ItsM3TLAmP6ybMatDjvaYKTr4hS4fXkLAwiMsR5ZM4DOb
W8GI6H6fGtXlFeqDZ12qIYIQa8y2RiVhyLCJztgOqjNv2NRrVUlVtsnN6POqj7yxj14XGzlu8pPS
5OLcnBSJgbqmaItT0yMpaWk6V/rEd4cf2kS+Z6Lx5tNKU/sHdGgP0tFwq/5Xjt09HTcChWqjT3pj
d1GwEyXA8HZ7wgIzGuHvxComLHmXXTd9IMZ0Kod/DnkExhXpu27QVMdaib7xs/SRymUmeptfduN7
lj8UOQpAqwNM3N5ICgwuyEGwaWplNB9xbxxtxii3qEFOw+HO0bB9bQliAr8oQP0AymfO117qwF1p
nLgC5nYiTTDKh+5PXBtdeDTPbuLdDpF41slzM+iMdXix/qWoS1PIWoh/7zHJKjkSzgQvOxMEocs+
/AuziPEq6TLyCKHzUxVBATtgh7JVXqF7pXVWhVJwnPXM6hIul/j09jkxZ57x+AvDald1Zn6ESbkG
h/GJv2SY6lBUA7XJjdSXH8zFG29OOE+tELLY2N6zWY4qMxugshT+RWKX3s5Zp61rHKEO3o4JaykK
4oFIbQzDCUnTnLvLoH93vqZgD6URONDcPGK4Mtgx+evq1QwtpT9S8tRJv1iH5in1/7s1VGbkZRo3
7mH3tOhONVoftBo1fcdnizLx74atw/L666M6piOZr8RJLVe5v1HmgxwNiVyND88balBUNRsB/ezX
4kZ3bTowBiEOQ61eZlGmvqQVjY6zvuF53+iC7/U2rZD3IINiKlBuSw52+3yq7Myo5oOUAddGjYui
F87UlIe9wXJv2+toDsfsyvlCCQo6nM+NSa2uFyadDWp06UalBvNJgreE4CQdTDr+CL7FioDpyTxA
LfHznwiGmZM5zi4LJ7Jvzrp0pHHwC90vBJ9nIwfmfOMNdeBzwkXH73PpRpauUwlpAxbcg0DhYbC6
/2EvSK+8dV2uKYlqbbOuN8L/6I+cyo6B2GtecmzxSj24XAbJIQUYMpzkFcpcdfYLdh4tSGqByVVz
YHa5I+g0cob65y4omu/OO8+7x2g3br6yZ4VQCMB9/Tl7/5CNPyAGujXewEul1YEVfovMcNdO2Q11
P59gG95Dvh6HXjN8yOkocRAzyw1IXMVFTckR/hzgnQAHvo4lEred0w5D8fuAJRU3OvMUOOVdZX0e
4p2FiId0raqo3sh5ILODynhoHhW8maILmZegqw9qYKQbDt4E11/uw4pYrmZA9HoeiswEWJWySaNY
mcmI/t2AUVhCaYi/c1Ss3RkZc/BhVIT7777SZIxsFx1q3WEWF6gvg/y3qrAV3C+ScXbyFXGwduS3
L0xHP7J+7pwJWemalvfu4mbwsM9TkU5bMccdJPl+Lg48SYdMGImzDYUvfvjgwibzqX4+tJDMl42y
kuvPSRPcYXp1EKLWfMoH9bVH7gNYHZCJthpq8C+ctqJWqPyw/lI3mjDl51Fl+wShqv0P+omq/yNJ
ZSQ3aoIcgduA2CcddLXLR2Muh5XuDX51UYQixgSOkhB76g1gVFdTzS9hzf29Ka09pSK3enyb0uA9
pycr6dmRMGyi3WnZb8+4uSycmk8aGQKfmv9j2QqUTThaRWzNLv68nq6bCJ4GSlpaHEYmkbyGr2Cu
ZPYloehfSswMBpeyxqFoMAQvzm95Gg2P1is9pB79CFIl64SL6NcFUPuPjuBhjU46RdIvIzQGoI0o
SwEi0pAgrtzkbquS4IjM0OlfekpAUuZVS7xjZZDpDpLHQqO2MITb0sjOk5O2eBxo2KWutdtuOVvI
cFClFV2gKHEV4dsn0xOLmyKMk3Vf8MPFibo81VSiXJs8H9Sz5WwBp9ZiQ/1haXHZg7XMgj3d2Ly3
vOpTl7OtQAV0L+n6F3OYNg6c8uABtpTrn9MApWw4tV8wikVQph37DhX+LgWBs4BoIouonPhAQaJa
GXNyfQVxV7U9/kJbnzGBRo4lcXbQXHnkFS3x445U24VWGGefNfC6fEJRmUaYA4khRXPVofvVDg9t
FrIZdjg1H3VpOdb6d8YNUSUCUaSTu7EroClba08HjdEJQInA9PFyR4kZJ8Ckg9hYsvY0VQvehpN9
56IAiz3kxBa0f6N4CpzxSjIY1AI+pJMzTBcRs/1NKc+Ok9eDhXKcevq1QI5S7/2flWfuZgogTc8a
eDm7iBushU8R1R6NToOSrQpLN/8vacSXXzhc+sq0UJPzhJ4TiAYB+Umi4hYbYIAmd0Y9lUEoUCBf
lL6LHu6Q1irBXssyI8+oEs6oTJSZGphbM7wy6RkKzouScoQZEHynTtV+Fiikgs5jtJrx0lo1tQFl
BCRN4Oj92OY9d3W2rI1Te7XhwFO+Gp7C8bz9FvwR5G3kzTgWE7SS7CQvGYXnreNEMbrJfXa74Gqq
oZ2CBVt7oEQ2b+w6vgnGyc5P/kXt8tqDmwA09JAOmfBI6jy2DMiczNQDWF3Q7GkPpk4MC4/DT83O
29ak7P5hSx2vpo4RozePtuHi43OrwEFKG6xQCAj6JTnqWgzSmShzYcOQYEtx4+/kXcP2R8XB2A1y
MGNS2VNvK1KZYtN9tWEHBMp/uwhKuJO2+HBuU0gDXL047twtG7RDVZ2Dwdxv83BjVuB432HXGJJd
kGQnziwXvkT9PK/u4TN1s7Bdtoy7Jvm0imFb3BaSfgc4q1ydl1KAUJoCiDHBKmSvqycmlbtRUoTP
YoSo3Zh1JFwekjd6OzWTTo2ZjPJx4O43TBLQEo5dHfno7pqy5/rNJUoBP7gDPhkvMac+JKIBdqBh
oKJd1PFawVg6BGA6bzUXV0/SlFlxPuqxlLvNeI6gLtyfBJgpeTphAMup43nsgB/oj1i7a22NF2DW
OmXdodoc9OlBVrBavkjytad3HGe0EoVODdeo/7p6C/aC/JoLUGrxngwFBa20JycS/FghGcvrHw/1
YupRf4uTBswC+rrvzqKoWlgRZJ6r5cEew2AN2bztxadtnJXNf/QSzOmu3kuKdbuv9uyCU2VV2MMU
ZliIQiq33W+BUWwntSAC1UI2wl2ZEHvEmWLKVLk0naR9VTyCX8SdfCOv8tCQgh2SPITwXn0l7M93
57ztSJk/DBonZL2ALkM30uyfHV+mwP3GH26NiEQ+dxAD7FZjl9t2AI9bAjP4PEDZNLxXg2wrsBwh
4R/0goAsr6c9OleoJHQ7qwNx9zP9fnkW77BvVzahFyQ9vKvF9Jt5CLoV6gxiqqtvzrOo6HqOMHjP
aQPY26Rt/AXlkAGisyzJ9AocP1i49tYvny06EemurZBFVVgDxQnDk0OWd6LTcD9Cw1WlYrvJCFqz
7T5kAtY/OFh3KEYOiPu5ymsciXpLT4oKe3IprXUGxEy9I3mIKRxm6kspUpt2iEGdqtqqg5VL9DWT
IlaVWr0w8d86oO3yYJVhSa4+bI0EWkj4WOO3lwVDiomDzzwoCaw4QM0ZJ3Iurv1JPNBl7zw4JUrw
gSDNlbNgOIWXRSxuXB20btoLQsD/7WNgA+ZUQsnln74cjShE0hpYVs77pf3WBsYFf85vPvyLgvjQ
ayOzFsjpKMsr1seuLSIHtYpRKHt8sejqv5XCEPL3K5t+QMbrCykc1TCo1tWQ4343RLlMhaHK9wzX
GJQLKAG6hm/AoK0KZMqR/685t1onv9oi74ldYxkDBzQiCqY2KsNWkzuxVoIhAUwSKXx1YRjfltL4
WwEptFf4sSto4oDOPE6DZXKNKky+MyTN51/K1HV33xpXDH/ehSKBVM9+RHHHmQrmlg4/yo2ipXQ/
kSB92KZI5Ingi/4QIYy6e995f0BUZ18WVUN+vQnTtc7A4cSrxzjNm9G3XStLQFnB95GkyXXtcMnK
5UJcR7iEbznp/Cvu98nprQkAxDbNcSuaDcxINFF3wsh0JrkJGJQX3U/KJ4IjabgkOTk2GRMWL27N
/hvTKAptnsFrZSgILduxqtiYiVlL+kBKwQ6f1oNevO8nLaC8jJ1z4POtBtklQT00CTGlr/ZvFQq4
2NTXCNJuM6A60hSuS7OeGQRChlMU8eoGsby6Gv2KW2mn8CYSHx1nP02KkKK/GDzoS6QNKYoBvuIQ
RxMcU7qHPWuAocHIRBXy4hzBGROvjobverGLoYVw0HEL+U+kM4Jpt8H5CquyFrgpb2/CRTxcPNR8
ibbK2Av5ExrjBGDzlThBF9gKp89cY84uQebSZUN6X9lMIyHNXM5cJ6IsNuMDQ1MWOO1gIsW97XpY
365Q4rqy/I4kaP70mvS/K/dvOsAE9uk3jL2beTWrDVGfn4GwKU29A/KJbLZ6fqCPZI164+VeAEVB
WO0yVqIENgzZwOpBW7ZT12qcFsihlFB1BlAhfAhvEbe0XCNz4C3F24NwrQMnhYuu5tNUVW8v9e4J
AWQqKf8LuNd2MkeSEEk9S8FWfNlTB4qXbBd2uOXcbDeVuaE74txSBp8wi6qLkahDWYK1nf3lH+mE
Y4MTr3kVUgcCRspxuy001SunnK2IcWY8G4C7tOUfo83lph0ZPDliAZ3YQjMMVTKnqMqgBe8HUYwe
g89i8ySouSkvrbIU2DS+V5oEcRKF4Vpl6itnZoY7j2Xi8wtmuKx5SLPplRCsoPXbdAc9xclgUJ+1
/CPJXNh/7SA/9OlfO1tdNuRVzpaRa3+twRExVMlwAl3XfZhLkkCo1spR2vn3Vi/XP7tWuipCOODN
Q+rd11n+URouedJRKmXmQwctQWT++xHGO6jfC/t9S2aDEn1ck2b0UUyyRUvhuQZxwwTXUddZxyHh
ELAvFngRtwVgmI0VAFUi/2LYpe0Q86IAk28dcrwpoSU95Po8uUmRyZs4wPwB2rErOPH6cHVAlXHC
1ru+XG+KPaAYp30nCi7pHsDLuRDy2zY9JykmrnchpMCOqEt4XJcjYAK4dAyHiAGKSZo0xiIaz80D
KKe0BUzoyCmzX89Qv1OHLnJoJ5cMme656FOh1JmXinPrJJu3jQO7ONgYgSOLiw6sh4bJtbq9LAii
RnlvWFzLjmDMwXIQIB3BStaHiOwQML4eUUNBQEFWTfKVPUUZ/n1blPzLXIemSnhB24zLL8Qm16KI
XTGNj7IG83g+cAZcyn6XL3AZnwG+OvG2Tupybh3Z4VtDYxgqj8BE/UT3kGQAODUIhtzB+XTkAM2N
V04JPkc6x0PbpSGuZfE+Sb3mgryeFfUKTwGznBgAal9x5T1xUCANgcdxDsMtQFCH4fU3MGchqGc1
ZmHJ8nBmcxWcd8G0FybrcSn3xOwxeKO1qa3KdTKRfpB0YWKqQzLn9LouFipVEZJph5tpbbqx/pvx
FjOCxqc5dBl3VuJ3wrGEn3wwQCy5g4EqbWh/xyEWL9ELuokXduXGGfTTo4YMSQbVw4qtmzhZpl9Y
liBRYlB+VgSzvherkRPscDDBovkUZu3CDuCG9vV9lkfrOGTYIvtKJQlxkapDhCWawADm0Y8YiAib
29CUlbz/Ngf24vcxq/ROZoRrVrlT6qOItcSLNWFgrF8VbQwDtlUzKHWQtcadFXPdAuPOYTjk5A/T
7ZcaAqG1+HaATrX8UMcfvh/4uwvcdRx/jOA6vfXGX9YeNN745yjgWhDwoUDbz+VhXha95SaFRCdx
7Xi/Fx3kptf2putSVbnqV0IgzSp3LhY8cpIPiLTE8RyELEdJcnJau/Ky6aqXF0P4ALZ03fpvUb7X
LXlWY5h56myzyEkpJvw8MG0MRrDeL8v+W4n10Jx+AHVZeFfAhl3Y67GCoYpYlpWCIbIOxb46VZRm
EUhlt/Hjo/Ii1tyWlHBk5XeGTtWOgxBn2wSnNXYnO72RY7DwbpLqF21BF+XER7cbV5SE2YfwVWG+
ON/yc5c1WABAPuyWdWZC+rAKYHHFuFxKvAs0/aMxOX808gRlF//PPMde4H/eLU7BL6Fmb42NhUUd
MYgIbC0KDoU1+NVbAEXOKWwMq7I+ANEEd3bcLDQKeC+qRuqfEO7RvQhn8i37iDJJIwIMfL9qfsz1
DPRiF3ZXEB+NZnvRn7dq0fyw3Rq58Jk05HSz2wJe4gwQKhSgSjTc/dwfLQa2N1kJ4UbFKjT98XRY
rggj/R1Q+AHFq4+FnbzfWgU8bV2zXrgsexmtt0F8nhPBjRN4rN7H6rh4zBoe9vGjcMuNxfbb96Vk
sZXhJyCGPOhg4VWg6Lx0XMMSSEVnJR6TFDC9m1mrIWM6V78hhIoREO9SnTo6CWi3NVm5x6nsEyRC
HILcGWOJ0iROYxa4uWRaP+MqAGBRvi3Q4sCahzk1J6xCBrgTMJyyk9EEXkDLmPmBXaLET4D7g0Ed
7OuUUP1mLkMItmhlkNuL8FdxXpwZYmGNttuUQ33FGKJejXeJA7L/Nh5Fir4PVpISSV8O+9N5PXvh
RfHQ+p1N1aqyEQcT271AfTvuEd4n5nUxUmD6PM69SAxmcM1ZR89mQQFVaTWJv0YfeYE7VyG3B9Hi
/SS9uAglOAL8/h8NLjWwPJOKKgbu4898Q+QEpwhc5W4+Q5Yc5Nd0/EkmMUS0Bcjf/GKliB/7I+kR
qyaxAxL6FnHN3hlsZpQLTGofqfk/ZX470SLFt5LNNJMqerNlKeoZtvDhAyYQxOQikYsy+dySJw1Z
o+IIs0wCnd/t6giYYl1ub+G/+wEImtPx09FtUHdNrtlimJEakKGyXBiWArIuHT5AzztKQ1mdo87i
7E7wCu4o3LlkeDW9mVv+gTl7QKbzUiWdKCg/bYgocuV7igPmH+s6suYPx9Cs9qihpsu5lMVBUT5w
YXDXkkURcO7FT4Or7ootjcwuxHvP2xxIbwp8hztoJDDYWypiEtfO8tRu0/ZNPIXnI1+jUSmmvgaM
nGJfpCriNmj+xnzh0K+EKL14eDTASJDuyS56rAC2Yv0EJ92KDs+fwm6eI9korbz9+ejqBd3YbqFc
luAeH0B09NZyroUcVhyn58WamwQb2iYN3w4NX0UA0apbs1v0OW93ubiJTwNrC4LfVRj9dDTYj1zU
UMihTAqFwUNACI9UoLI3bkEflg+4WgKK5wdPbsRa2Pzd2AjXw2nWxdYjP/tBCfwZ0p9AZtn8OHAY
CQMS95b71+M9Ezxdx2UkoLeLGPyeGMJ8qYtOyKF8pHQWMcvq9OGaLUDU8A58hoNDpqBS3fi9JzDJ
OIl5Ir3oP2M0tAppoX5yUJafKtH8FWHNpDftMi6Hh2RGOgNuS92Sk9sG0wSlkTzuHrybzB86jdxe
BysltCNHp/BE/fT2H+7Dv1XWysk9RMYuL73TS/jk15jRBSOOUvWiCdEdG5oMdT/rT7NLg9I1Opn9
9xpMq1gNKmYXpl16e07r6ZIPDNNy0AdkRHFCOwqf8dSu5cGQgdxi8Bjzmhos9723lOnimNowI2UJ
i7Ghk91Ll9JLyc7jQbeNNfgl6cduC3iRfz+To5khHycpTl32CXYrdLzCtd7yvMkpeTWPj3HfywdI
vJ8g1o4uG8DcXPzg4KU9DtFYWaYTKfWqhnjWi9XhLZBrh1UU6+J5CJR4qKv5sk9OsXKfJ3kEVI/8
4n6Lmu3PGQFQ5LBGUVIewraZT9bNXCvohaaVeQ59/o3qRo8YFVmDVzg0K97vjB4H4cIVxQbf1oWR
XpGtBuXvl1rpkGS40HbLzy0WlkS21nxzsNQHkUH+sCaAdAVRo8muzJo9R5nP9VZttMM6PvZOAZ8C
dHk7vVgDkzqfKLCa0O1Y+lBlngwrzWILvcrq5dgnKYEoUVZR9lAK4/8y1qh5OpyuyBqXsNvUQYfR
0jK0LBVd1Xf6lELMjHjbYfGq1VcfY4tU/MGdHXYf24GHxFslG1TJ8h32GazGjEvYGyi8GSXsyE25
uD73UFJN+1I8dVFGWoAyCmmor1bZMUfnYcTeEk94j7l8RvzMIfio2ClZAr+BbQswx2kFAKiXTIN9
ksOJJPHmLWOIO7w+tGYpHEMwFVWTkSH2wr0oB92cFjtT09ErKJOth5wxzBOB+xE8+GS4SgWP+EGR
24vd/9tvv/N6dyT+GF8W+GimT/ip0/fDK9RFTDa/sRwqv1TEJjhl+5D+MjAxEAlI/COplGOaMASe
wz8mHm/UhJcGkmA8fGobq7aMex4fGDuTULwhmtOGMml+iVH+jQWTUmlVLGtyhjn3UKTYyhVRe9YC
FQrwNiiNfV/abA27RrFvfcZSLMm9szNg7KMhxT1eLtvdMM9mCtN6Gwb7w9459snJ3jo7amPoqEjc
JPjFl3ZovPtMyx/iA2xFgqUmXCO98OK0iKL8lRHZzrX4EVHza5R8ZpSdzskIzMxEYgLhRSU45W5y
+L+27LFAwJ+noCrUVtWfl2cXiy5qOoCYorJvbemCgn04QZcEP6pS4MolgJizHJBqXIOu6jRFRxgL
v+H1ZRoBSpG+UPeCtVHLEZmWufVpxDWAQSL0gxkoHgiGsGbBeA1TkO/acAC4gH0IGU+JS3kuVkoS
6K0Pm9MwcSuINW9p2ydIxX4GIGLUuXeuM4NZCHYx9MOmsbSAaaD03mzcxTZJpOWUZXmr+MdAcnyu
rXZk0/zAXa7bKNU+Y+S7iuMIdcbS0ZpJ6iBUCZ/9ouszvHB0D1b742M8gjDwJk0XlwWwOfOf4LKm
cFfmlCFYktR+4zdwgWiS9b91i3NJoIrYkXte3rLMDNWQeDDpcyP4AQOu+28j/qcKE5nE0yh0D0qH
anrlBnsYqtFl5R3yGjswpsgz1v5lWa9Hq6HoZ3V3vViUOIjK3RoYuXTEzi5zOvQ1N2PK2gXIl2HE
K2Ipz1WH9f+sbi4Lcf2b5f9g+f/MzvrvX7L1JpARIJFSHFdXGatAcY8UY5GX8YIcVCgzxEowhqjU
Nst4oXwSb+gqrY2uYd+DgYF9lHMpJerny7EenI30wu8325Z8crF25qDYmMlZlRbzjWaZh0D3I8Li
F3hR2nonNg3u+4SPoQ+sBYPWk9pny1PpVsLwPC4LEOwIYG8F25qhdzkazX1JeBu8A+3s/APG7711
QU2+P1brSBlWL1AfFMD0qd72Ven0ianl+ssTp6WbmrjgX3+3u7S+CmphoH1hHD9igyQ0O2tX/mQ+
c/VOdYIRZAckD9jQ94MbXfhVxn7pH40nM6vqErD9vvHsjEgPl3Lhj3tGV7DhPm+oUbF9WFjxjpa2
myaK6xQN7UqozozIYKWfkdgn77+HoctOuoaMBlkVld+c+LnrfmurvRvLFqf2iFZeXpbVKPn6SJaE
oigkj2gpWQhIHQa2q8C5vE4Zz0WpL4EZNZdL5WNvyoeVUdsSPk+Fgh4zuRMQ8aPXhLMCL3Ap3XOp
ey0NtAvoQaxzwws7PLvTdG95gDIY84ZLAlxHJ9BBAIljS4zm4uNL7KEiIzNHJch9MNoqTiHALGcg
MjDPbdRxPIGOahUYeIsmO2nKQIeuHlMUAtE1NTyMCDOrff3sauSqvSQ6F/GvwTLTzlKnyzy5ZPBw
pck4vVCEopIer20iDFvXi0KBnWUPO5pv6ncnOYt9cb6hiPS8LiQ7ZNAYxGvCs1l2L+mFLzkXKZVh
5N9boMtJpmH5FkqMS4uQ8Mwk28rno03JQFFpFuaUSKMSWjfx6MRE/PhKpuDmssSSj7XF2rdEEHYV
Avez7/TaNWRUBxd+aoX1XdTOvkQ15ZGfiTZzX6PK+Fgxoz1Hg8sC1eSO3Ieky75SImCaK208akdk
3Zvv1NCBJ5lpXzo0/M3XRdouqA0xH1I7eb4ZQE5H9zxIIovOvSjNFrJxRtfVFYwFSoMDdQJmtwz+
5SJcZiHjrDFSuGc1agSiSBq7MTq9a9tSMX6haLtD/mVwZYX5ByZmowDtUe4hFF9PWBnea+jJJVpS
WUlmk3Xo8sHH9LdfbuF1DyXzSR/lK5JoP99NkqZlvohB7DQOp5gnkySWaVfoZrjryWiXe7SdAbmK
4phgYjgqdgAyiGUI5yLSL3uvz7cEWd9C8nAgaVyK+nfwZsw/nCynjJRGjZph5Tq3RwJHGBHKg4v0
+8310BbrWZ0mvSR1navpKZcorelSbEjvqfUXHjmk7ZC2GNUM5q0b3dFJHFGXJyJTbqIm/j+EO0xp
wKFMJrgmu2f6xiwkfbeMmoY3xHoQ1Babm9EU5UFGMAcX7vjeed1hMGyAEF3sr58hlLffyIt6Y7oD
fCB+stK9499m68jyLk0Qj3u/hfSndoFaIneBn4Id/BtIm+3UY0QkJC0PiyR6bHSz5fCetSX/2Ha+
gJMrZXZn1J5O02PdJmW+k1TSA/WPvXhiplpHqCQlrVfYo35Gpt1ASdKazu9bleDacKGy0d+zBant
4X9ptU1ekhNQCbzOf9Y+zCzG1+PdL5OsmKlgQBfW7dRVl3m6ruV9TxxRgxKSEEIGku+qGSGZ3wLU
otGPfHpIO3mdFng1bhBg5UK3Dx164+hVnmW2D4GLfe9L9MG60/cxbnMdcSBHRkfTB3YG+NvWYX8X
6uGhJ0lnzYWfbTdm2EhT4TaycMhezoFIm81Pgg88U2zr5HRN61LEuUIm1YvASTqj86NDp4tCgJgA
xTSu2EeI1oU5VmWl4L/ccdJMJGceAroH/AgtqhChpsXVbIMNCiWig6jkymN5qbreT71UQ77T9Unw
eXPfSVHVIHR9opSUzUeqHv+O2l4uaP9EnJQHE/wNE1FrrBwIiTb7mvUlnIc1W9waGrbbm7PvGqwF
5ZX6EcoHrqmP612T50mZKu7mPiUpJifjGxc///gc9uaYtDwn8RTZ7KNMb9SSvcb48kgBz2B3njFE
0AgUms0aCSxWBVI8CbrNQ7FUY91YZ2lVg2V/AD9j9IKguyMwnWIiPBuoWF2C45Gpz5hIwFSvMdo/
S9dhuiYfHTwYow0d3Gwt/p9g65JsslCEoRVr6QLZA8/zGgmiADVUYBpCwEOvez2H8GsH0s41UZ6P
uVQVYMqL0q2xbVF8/e/IniEkhqX0/6G3HMzVQSaGJ8bUx+BwQgT3S2YhezYCrag5CaIUZwvZ6ZIE
6HyWvkSlZysBEnaWXggluu0fxFAmzfCG4lN3a6k3EYS2NzPSYNbqfACuR5v1jzN0cMOfMRXMjNOX
CXkJgfVIU6LPHZhQFvdYDN/yD4Nf60qMBTixrhUqfZrKkD+qACA9zcbfHzIZpq93XkoGg7lV7amg
4mDXr8+237w3mMBomyYWytLsTdO8+3UjARRIaStyUbHqQomJ+SrJRdpKrMCBap1pvkJhIeU16iaA
XIzBEFMaMmGnBVITtUm87vJoTKZWT/rv7zf3HC0PkC5U+8yLcrkgGAOoUNT3Ck87Uqf4HPl0VbQF
caUxB0Jncor2sWtnmqMNm2eSWuCKBUmTMQ5mY45mKHqo6zJDJo9g5ESYMQ1oStzuOnJ3Hbm829/u
SO6EJFd+sPP3B3Tl78JjngxgbY8ruEzAEd2j9eXuv6WYDh8w8fNo4vK/ENfm8+g2bhD+W1vVxdkv
/PgTKqh86aKNWpkZ4dCxhA3hk1wgTKt/r2nFAX1VstUTOTOhv6nB/zK4BcuVEK/KwyiGk/7eA8tU
sRHIwPo5nUxSXECaGDh/Yd7IQwr6j7dJ897WQtdBRaYAZUcH9f8TMCsAbx46UGURxzX7qO/humL4
rg9ivaWodPeyM+tImx947T+r70znHNdUmjxM+1TsgBhy/rNIFc8BN3brTdImMdsyIvDt6AOeRYcs
FTKjeVG+CheSPhM0SfbMF1Qh0pHy9xDeW9u2uVRuEl/yJgiGi7bLxr0+3Ylx925CgGHd7H+Guzv9
R0CCofE0ktOn//+ivFmnVk6zg/6uzuMKR3U3TKrCBPd0M8MlK9zP5zaSG1D18t0l+wjclExk75Q2
FMPKqEt4WtkkDAMpVt/kHUy+8K4x7Q1twUUc85kGd4UsJ09Ed6Ipeuyu8kuPwrhmHePwiXvyjbFd
xLcdRG70jL6skOyolxiJw0mGKO4K53T6LFBiM211RHwU/NG1O7otHe2+DCLA+YVf8kc46X26hA1n
F2N2XkufDki/eDEyk4Hb+CNWOFx9kIrWOG5kyb9S6y/sz8IWYvemGbABieIuniTF+19a+97+zXE4
aTzou5haDB7OINodkttVzeVUjXIFQ4cCm80cxbTew5ebF3aakWEV/jYXSqyQfxm0KgBPUeyRTKFc
bksjHfV236bKbf/4SVmVi9LZsP3ge2Cl2PYm5f9SxH9unpEeyzXavT1p5XfmgUIY3tYkIoiTUU75
WneSROmPcF0rPqOyWBISLgNMymGlmdQxeiKZSGylXO00ttPifooMog+NRd0ml3GLc1TolVmdl7Pd
LkqKU2uGtB1YWCecFU9LM35Rbp6BGONNOeMQuzqbfGYwkuVytzLX10XcIQxfpQr2M2zARaIdRNlY
qJnrzdpq9mOFP71LPTa1YbbOY4dvPZSKvqOn1MlcLg4B0VkSgYBg4StGD/l17tsniFvqwokHvgct
8V+k8BU/HTrd3CNE8C/w6LoMruaJOkUEG3aSBClQnbwYABGiXAVo0zt2qnpbQQKd5XvM3dRADv5j
IMGtaWOLHdqlZA3DYdXyRazxSd2/OJvoKAi3ScXJLJfmECjgQYYnba1PMvcsiB70KW8XdqlHqIyw
KUmY1ozVMPRiaKimCcEZLtsvVzic2nfr622+T8psbTqg3vf0w2aUkDMHXAfsTMGOelqPRIma+jgY
cMitRqB66R/y/jw/wlsaTqUfp49ay03AXa3FJI+pdhYYYAZNhTDuzEvCkmgVsk8JQeJKMsAH9qX/
w1coQzBrNAX3eSbxOhWbiTUGO6kLWZ88CK956nSBKghPYLYKYDwt8/rQPvoQ/hBf6lMlcj1GkjU1
59yOm4lMem9N7HsXZ7BZ1J/fmMRBegBCqEzdu7fWILuLSi+h0fb2wN/Xe9XCoQfG18PCdd8sVk9u
l8EPQaXQC+ft4jCXUm28cs6FmkF9iIilxSyF0teUXlcIJ7iOel6IBp0ZAu7Y9OQ6mrj1VnRy1O7z
67g+RGrBNQHc+RsAjM2w/MvXplRgNFXxyIOjYGbMTTo6vyp4eXsNQbgf72ezcehyUF7K/JQuT4Dw
Hptw9U9A9/aQnTU0VrMglNkfWJiNe87HNmdGxu6SvAavNK2VnnmbJVI3RDzqlLeLCZUWG5A4BE3j
8/U1Yeg4h4DCes89SMSKBWBTwmTwiV6rAdLWOnuHSHHo/R0PVYAdO2pjqT/xbPLeXbVYWvwkIHtu
G21VU5/l8WrN6u+uV60+cGePnxyU+sFB3tZSEfYowpXY0UaRLUJDPHU8EE8W4UIi4bgdLM/tu+Fo
3FRbhdgHV6qNjPxx1QxUvL4cshi/CF7v5w+vnR8XnH1ISSysMrLusJoNN10yAIjgpD1gzhuDv/5N
j3ZCEJ0D+nE31HxQaW8wC4o43bonmZpKnAiuLhRObNeySBxdFs1Ehr4KL+OX5bTSXr0HFDLeKFmq
tuVjj1RcsuPzz4XPRKJrDUaOrvQ6WwJAYTWL7S9FzzY69rQL6TBR+h3F999JEpqayBxY5unkA96D
EKITw5wxZc/Kha/KjOGq6VTdfEn++a4E/G6nr8E8ATQoao1ArCOYpM/b//Iy5e4LTJ3ESTpSGCVB
rSflJDP0GPPU23qayjBqDDRnh//f78Z/dz2zAHb9/g/H4XzNODODNhZYrEXUngvrpOULZtvS3tlw
DcYx7V70GuqIu6PJsxUYWOemu1rZNonYuRFjZ/s6AG0dhXLKTFWvikghbOva3VrFYP1ahZ1Zc4AX
zqUQuSoHxKa63jrbMnJdhtUrt/V4IkJ8JkczApWxv2d/0RENeWuJFcTZ1jPjuyfTFmT1uGcFVa9P
HW+OLTju5bi+LtwUks0LNyOkV6nIMsvN2o2FhAy7w1ceFAQ5hk92DsLZ5IQ5D+t/wW1i/Yg70USk
w5ZDas7SXKVWeicXZEKsx/RWv35BBSl+Qr0CnwZFUxGm+4bxmYCD8hfCqE9AvY1TG/Y641WFVV7k
4o5QTL+nugvvH+WTssiTuj8WdrLf3T+RlwMnBnL/sGicz45vHQzo6vlaTj8RRRlYotvblHPNTWdm
jc45n4XRV1Eh8unqyXwzWVcXM5TTfoV7paDa8frjnAimz1dsAR58cp0t6bOZ7J7P/Ie/4UeVyDU/
Ydyu/qM0TX/Mmw9QSrMTZmOMKyXnGhkK067QrYFMsc9GKQskhfCW8+hjGRpGe6qWRTCdAOCi1YRS
i0i6U2pGovnC+oCnONTTsa/fQIc52VVbUuk0Qo3Jx5rbOwSdX+SGpJ0qNVfbcXY49W5Z47Tgh/6k
sdAeYhaVmssoqmpPr+n1MURmbhOAS6vUi+lXmJZhUZJI6zArbRKBAXqE8Nd9ocYv4zeKV1uyzKKY
XxEKQuX1XmVgSogpqoRzbsvrSxGBUUC6ZvynQ+1oYfSE9roSHao8vHsh9g9FXtcN0lW4cNSv9QLK
C7irL+cJq6pYR2SAGD7CdoLewJ9nN/j1QutejAW9vqQUAGI7p6A22T6Vpt/7x1VJEdzaUkVfy6nK
9Il/dO+vKCBKXiDZTlVGKIcXvHvCtF4e3KZlr96wnqZ9ArzZBqt/JGVlmZ08HROUf5Navxy59cXn
k4qUF+spkt+hB5uuChPlnGmYPu8gRAqF78eh6P7T5/DBcR+ZBCOaPK0GTrMWvhNjJ7q020oeB8/0
rB5iq268LgSTKd8yBYYE+PP4tcHFPigMol8SVVqZlyaUvde0eNdBJebqdUhoMNx7KJsvocmJkbxE
hxUt5GwuJC14PZTtY+ik1B1h7h34EJS3+OVoU3O6z2j40TCR04qvpjJmvtPOpc8cF7WXI9SeoLTO
1kw7twjxjRK2QBTZS79SmozUcvi0Am6+qOue+XT6tPqiTS8HfALqsjoT5INqB8oXHMzS2WsMq8tj
An0lXZl7mn9rBvClrCau4IZAQYto++xkBGozIeYRCytzSOrK5N+aqL8iepZdmVuSgYqP0qHuYAgA
KebYgiwzAHC9E1tdCYblyvWcB5ZRlpll8kfJZxUEBWI0BUgonM7dBrCVI9AmiDLhMDhe3eoUQ6C4
UNXEiNXtaSyGoi5GZdy8nrn0MYROG0qzkqSfJHtakRyj3tdDB1p+nryevgikrwJIWa1QiW2uGRVF
lFcSoIsqyOdeWt7HgCVcVwPHfk07FUD0uCzFaMM4VrX2ED/F7HAFMWswBI6FuPJzVcaDx+K3DalO
2mZ7mgEtL3N/dUEYJecptb6riyuYWFaFCRXiLwPh/lDjerKu/AgLrNDFXyEwtmDmREdEoCUt7cKr
2PUEjmaQXol34YCndpUeTZOqbzQxjRrl73QRM5PLXTrqxBq/e9wyjAZrY2Xppdo5liR4TWYm35K0
myRUkGF/fk34Pr72nqlbieKGO4lJueI/1cdbI+DWnvNDCffp/jQCkPvrgBWUga9HIkIEU54Edoyb
plk7yey70QCZFH0VZcnTaMmmoKi8zFelWUWwZtnADI7E5soKbsq3ap6ekQnlCBlI/eV/L7TLjiL8
odEpW0+HCrWC6qsYxG1k+2/Bnd1jeJJ+em/DGh9o4EIhBXxEmh2TASBOyQrzGLZMzJ3gA2DbFshN
aAJnZSf2KVIajiX7HtTrhRNAkUnPeserNSC+VyZQnxTj9So8FthSeFhWZO3mZScqUBxXnMM0U1bX
7UMBLobuCV9HASpbicrD8WJQ1kfl5vCD2EWiKO+DURW9oiSIlu+GHzuBz1ngLs5Uzemx8FVflkgk
GEqINYK7Kd3muF3Pq7ssjz3pyWa3WBTMhfXR2g5lzYiZPb7gQk+VHiJQl63dRrw4cayZCjy0tljH
TEaWI1KhiFYIjsmManzQ+KVswq9oXVb3XW6eCxv7wExceLmoYJd6Avl/Guz2bJEzFUc1+ACH/1fg
GmzNd8OPqfiLijo8L9OfzMqs/suUmordaivXUMplUnzmH8Cw0itTIZ2E92gQ3a3aXaSvjWq55tj3
gV7KR6fZ9UnmydUL7l3E2HH3LIa1Cp3DcuJt1/WvV+d7j/iOoN4qSLT9yWuW3UOk5z1dn7zHNbzQ
oJvTPMEkPeoBBztYeSlHTpyVJzxTPcPPQwflb6JsDTVe9V6E97DzxrOCFndNfzJnoKhNjDDwknwo
ETMZ87mO8yfAHlLA0kbRIpaurofINdsslPURSI0PqgrCc3KKbF/CYc1FbFl57PDyLFVBUL/niKWT
uWix/0CdhUFvtuRov7K4/Zxq18gjQ/9KyFu9G87twG+5E2esuEXfb8Cyre7bFUFlVVnf5AkU52Tk
DdkuYQ/RKVFcJokvmZTnEH1J4mh1VLYGr+AXpJxCGmFB4DLt6LCSwFqVTfAYHkClqRv1a3NVmet9
nbhgJy8vwjwPGENu1cxLvd8Mn054t5A6kc/yDmtY3U49CzUDl62w6V4wBuPrLJE/W77t0U55+4nb
eijmLwmF2dqtvBx/7JEXtuKAYZwnbeuMKE86TB7Ekkz9P6cVzqCpWdkRSeMujlk8sHQxn7Ipo4Jo
+S7UoCPwjrr6SeAEZ/YQxKuQb78SZEAxjeDI1IiIexojaHANrhL78PAFWCwRbIx3k8k1lIFKbda4
E45KHc3V7bgUArN4s6W7nG8Q72S9EGXJhNuZakiaJmlJgtjvrOITj7HXGYXbXVnm5CQG8DEpGqig
571cSXnioYs/JCI6fsKDInkghFt7zbQ3RBK+p6yBy+PkSF1z06gswS4DocCn6jAupwdGMrvbK6A0
wMPC/mVEzn+PwgLA40xV8VYOfLkia1kGVNiL08x0aB+hd2j5lPRe5Un+CMaHm1Hl5/P/WL0cwvOq
cQ+6W4M6QjXiCx+Nh6w1FnQ45Jls/zaR36FZq98s0HEiMUbNwWVBGVB/3E4W51b3Y7eRp69PRQdT
gM1eNmcMdRcHvddtlSf6vAsEMdOpFla2Xl415Ka/yUk4H0RZnH9e/ADBO+2wYSu6mbO9aLIUmx+A
6K5kMzxDQuGR8BypRcnEYu8X64GXJ2DU56Oq3WbtCPhicTpO9p0N3NowlyOfImG/dnPnRBtBC1Ly
Bev8Ix9zOjpfz2NKPRSzB0EyBPkjkF239pipChgXXp0AlYQSYtzQcQgXhy2rIrtrNBeDtmosYMqw
PVNX907/JIrZX0BcuAhXKcym1bdOmDDKKY+OIHceP8Kk/jd+Yq5+EUr52Zgm+gBPSpadjr/lAaBx
xO25Er67nvtbKib3RwT0SKV36deOWTpumwKf3St9PQJ+CnBRhrFpI52N/U7Mmf/mXvtR2nOesql/
9vjxsd4aUcbmORxim749QC4qHSvT6GQNg3+71s6+fypx7nMRD/31/jXp8tidQ52vr8k72zLoL+Yc
Mv6HX8mdO2ZGN60qyGYTX6WpAJvgZmjLuXsjBcy2cw8YRQe+iOS55drILKanKVGzjl7cqcPoLmTg
4CCX2CaAl3fbTU5xLWRgVMHrImKKirCtMCtr1uJ3rQF90JIIl1vdLo1FzQfm0nxkqPL2Hr3kG2MN
5r8XileNqwuMl+wSC8ww3SN55q5S38NfOs2GR7317H5exws0BtsUiWheVM11uOjprk0SSrOXHakm
wYqiP9biWW2GH8bUIMXDDxODjcq7vXnkLspq3rbVOa4ao5aC5Z8OQsqVbrZRbCYFrLQdqcaSM4GX
HagULX/0vMhOEPsiQHYmOYfxWQivjx7YvumbdKyHt6KQN6QsFzSxHcuzFKX/iMlkgsb8PuHOrzSR
rvRy/HNcIEYUgKnXRxO3Kyi/rL72rHuuwLMD/S3dS2TFxvEGblxVu1r6XbXEZC1k3TrcVkpdBMC4
i9TQxCZE37NpfQpkdqFmTv51+OE9tiW90eYjlcOEKX44x19qTrxKU44mZcBz3hcvuP7sWi5227Vs
9wfRGpdnLk19myqGhDc8dHY0FJpJVA/bvtjJbuPf+g/5QJleLm1+ETIRk3T8wq2Nee3U+eSWRJKH
AQ1U+sfcRxh75KTfJRsBe7Pt8I7UsJDfkMJhQ2qg5gem2dwLDaYonU/NkWCuFex0KlVKHG6dGF0J
7bd/zvRmjNc0/YCqeLIUjp6a+yCSI21KQHy8M5JyEGAnNYNO5Zk40OleqYZYHrt5MTA4m8c7iTtm
LZECXqKQUc/TsF/++klXmUIW+234fza3kAxlNS/AV0ni9sbBjXaLHi2tM2XJNnCHK7bwoIxeEnI6
ISpTeZmfh8GlIp7zXM3YSa+2l3naf+q9HmJ048m+ShYLhTAg+Y+HAgXuFNXo3iPQHr0I1yAWgdb5
Iv+JR1/VPdVJpc4oQaESemjosZ0Coqy/AL6eq7EMqTc35T4jovvBzjqR05k1hqSWuS+etzZJdC28
N+WceGvDwSZs0TLMtdJXJu2NE5jN48t3WUna1kcS7K3rmtgVmWRh/ZZQq/l0WEEA5y7paJBhuv2h
3dYKvHXKUfOVFcbr1x9rsGFQ7Nwn0jUI9gtLFmT+xswtqJvS+TzpmUf/BD2SsJHF8nAIr8pUN/Wn
PxnB8RU0dLDyZ/QcyBPl2LmnoaoRtgTA9PIlHPrSpb5gzfC7fLzelwab0KK4Jc9hLh/QSrVXKNsb
8NwaYY5WvJy7houzDA/2neENU0nvhXzMWpvuq59CiWG0FqVOeahMZz+66aZA73LZNU+JfMmsPUbP
G5tyOqB3MvUt0Ld16LbXF1LN7m56wxyESeIScIvWf9Lnka/sEkWLovqKe8se5tOJln06TQpTmHmR
YSki+/P6ML055mBwRozoOwZvAnYKbnjYC5PCs8P8WcHEApdGTslqYAdDdYuhDwayZfNEd6otaCU0
gyx1QuHtbcYaOepiaPv2I2ZlKuG7lDzGfJj5fTCg+jqL7Ro4mNN1TYTtym89hOIOqpPQ8qUu4N8n
K6kNtCmk00UAoNAwdqRKk6GGutQP7d3HiuCd1r2fYWQTx7c6IIuMf+WvyF4450ElCcdK3B+OjPYh
plx0XKM1Qd+Hp7dxS1ygXcwFT7nxamDCqU3UR5dUnJy3xURfFVxxaKfRYVrMt9vqTMw7yHrvwfZs
Q62tX3+UgVjMEvYkk9FYVfWG8YPpcogMcV8r8Oe5saed/YmfBSbXiGt63KuIFwCbg81VrIA+9F3f
NEwmqvd/JB5kzjhqene5IK84L1X4oY8W0UAR3XrIxqIUQ9rY6Y60npQcBCEPJgHfAzYeyiVXAnTX
AV9XrsK6lXtJCblT31Qslggj9INadwFCr2jf+8iZTBv106w2eqVjH1MfG85bGfwhlb7g4Bjh2lRX
4MTn+CyWlkhGb7ViEq8xrqrlKy8VBccttXLjCFAPyUcxDMdE/g6xgKXgaoZwYmsmuVsWY2caTGDh
Tuzp0PEvbTX8KCvl1Wu9t5Kjib8HZasAqHtM2TqpqnzhFeH+Ku3roSNJNxYzyoXO+BVmK6Y37ckb
2U4zI03ufX8+s3X+ArrzeETkEIYi6+e+AlezRcJZg84sBhLv44+F0x23ZL7bddJRqR+QAF//4RRE
gc9eThb80paqUVg6aIcS74GxhQzAzBsXfyyWnOty4A9pfuIB0l6AVODv9Itl03No4qOX0xcicW8U
sfiGImgbBPKtTb1ZK/uLPKZ9ky02p25rP8nUsyOz8qrXD302RoQWHFRL0ep/tYgpQqStekhRtAZo
gTQmB6uPARRGnVQn4LZMZ3y5CjxvzkkIful/EMutsO5R1xUvfhW3XO4L8yZCiTNWqeAPfQmrrKqx
MGvzEYvxGPaovLPn0+rRwl2EfTPCXsLxKxHpf+vJ1lGAw0YXeF/a35cEmabnzDlb44mrXksCzoVm
zgpCtHB+BhzgvZuCLw4APiUPM6GscKFwp2TkgHBqpWwpTP3bM1DWnn4yzpgFMq+dfRh22RpgrRVi
iQ9VvwDhWB6xfd5IvSpl/rcthqulK3tfDdDpVYHwB6gevF2TUUQOYbAwnLO6VpbDgTJ9f/4uBiuE
W92iYNa6jX53+EnqnkVJO0r5mw6KDszK1T/WAgUiui3wIiXHkmFTKY9t4WJ0aNU1e82fSS7W12bO
IQD6KVUXEVEXo9jRMZ1a1Dkwa8eiLnMmwacATzKeJLbHFEA/lY0852wzgOVL7qqgzhIlYRU4DwQe
D7qUIWr9Np7GRC4tJdUdv4uj/nf/eFbZ8NcQoKIDeV5kZdJHNZ1fTal5ZWzRM9MUqcQ/ScomnMFW
hTjb+wqcvjfbWHcOPZJZPHkdaWxVuT0H4eSGTBqc5pOPZIs8Zh+5J0Y1uLiddMAE1QSuBRgVSkXS
y8ZJZiRKlst4RULr/Ns913tt2M+ITIp6WAzCWEyCzStVrZMgwoHPEJ2NsVtOZRW/5+QcVYqUUunZ
fFvXKePjcqwE+OKjJ4kR4NtW/4iAF4QXaf9v8wvt0siRkf96cB45Icrr0/tRPoUg3RQ9jCtKUlAr
YH8mGh/r+mEyxQxIJuwmqsgLDyMwgh3ZmriptHbTJ96F0KIx9hNMzbbRQjasyPfD27GkPGRse/DX
dIRQzba6XXe5tKA6Vv8yzGrm2AwOwD1asHH9m1Z6pSMSTJ3DdMIn80izyf3eAas12SBQlZY85lA0
tf9e7EkJRiLH70MrFSKsKlOu7BuwuvHV10LSP4UbBK7gVGWfrivD4jylY+r1m3hVBNkojwHuyvH8
cTXP+LiHkXgFnCJRY1U+gD1UulxObctJoFsL5zL/PpmdjSaK/A+ibR89RKsF/FBUI9X2VCeq7ABI
vtjz8gEfQrV8b8aE93OMURqypT8lhPayG/y+Oxm+wS3z0c+k6zdD49G/FRzjA86ptiODHLjwHRjG
/kSkEzCEOELEZt2pgm2I2tlcur04Pq/Aly2XsO5B+My3yoxFEYKSXQ3INxUDydnHYP3M70i3AMY6
ks/zxt43pk8WudUL2lJuy3slF2lHRe/BlKOEWbWGjatWbrr5nJBIkQJ7jys66Zxlx5Rp4xKUrdjc
WQOvXti5G0QRkLIEY5lLQ3LDOYgKttMFk8Ul/m5PqQkLJz+WvT2Sqi0qykSUPTqfuzXvU5cKGVMa
o6Fmu8T23viC5G0PuWYfOe/8/4mDVvrtEe5hFFgAsZ0Nq8dBRPqekGclyXu1n0dS16BNa02D2eCE
ZwKvtiNnfzd1utkJJ26egtBWR8wIR5pNMg4kcTLgBaZCr37aoMT/SGHbRmbBH1F+s29wpogK81uT
8rKJaYtt7WOt2YkyFUOlAXz9TEveQVq+v6dqkIHbH26/pfwpenne5l1MU7s08OMN2ToEe7rxMGGu
2mgc0JkPZteCxD9I/BKS7rMDbOsCpGSzASsmdgCvzFgO9qe3KWY4AR6/tJGJ+KDFXR8Cui2MkrXi
5V1CSudg3rMJgeYQBIkKUOn/djAtHoivmCCCe0Adw59Le6bq7o2V+5z6OO5o64Aue1ibB/hsvCCo
qv6nswA51eIvdX4fLHATY/K4FFZtsyxt2DPRn0yfoOS9/zb3XmCoWPoPjBtRje/GPn8IqVtPS+sU
iwnmrDmLE6sDMnEIBX5r5742uDucms8voM5YlO3e+IW6qj71ajOS+mPNgcgMAW4n9weK/mSMZXSL
nezqo/8uQyMCwu4labIWy0fINxt9W5ArHJ3j0lF2aSWHE0TPsO/GM+SYwXLeAC3fStwGC+HA4rQT
31ToQJ98nH1aNXojAp+Ul+4t5rR8TDk+gQOLhs5N5vN8wHNDj58XGtM7Ay4dvorbaNbTddO9gj7Z
6lZQwYRrDyO7PIoDxc8EyeuIWBOHSK+DY0r9otOuc0YFmk2OptW+DGT0SzbbYEzNjtCRHFLvm1uL
M4JVJ+BdeJrbG3pUkvmCqDWn3FmXuBpsz+V9zwsJ1At5ixT1rz+GLBgWkAh+wl3bS94oIkg1w0L7
QPlXgUq+a/EB7GEyS/nq7Boeik+mtKajMxxLL19ItL+lUNsPeNwFK0p8smo7pXu2RAu/c9lNhplW
VCFdcB4itkgMbeqjy7Vt480uFlcXhmIEshJYsQE+10Pfexc8JviSf29BftXOhZCJHFe/4kK4ZgR7
C0LmZ+gwlacvbMnCeGTwAZyyuk4I3AMzMhOTE24TCWzJs3YBOYDy3ThOgXOAXQIhB9+z1B8expjM
+eO6RxXi7hyIpuRWD16GTaOVUlOV2H8K3WLov7IgFxmWuKmLFQqTgR9EE7RWrObRqorDqnJ6cZv7
ekINky62WjGn2lJKPo4p8Zhx9InfdjJh+M+v4rkClYhPeKOVy6hZCBlcH8dmQF6wHwyn1rO+A7x6
uizHM/KqAzWmQLIZ1zeGHGAHQ6070y+cBJmAnvFadbCx7WsPIsWHYHUToQVrVJee75voGbwSPCIq
AKovdsW8wsIMf5VvSaQImHP4s7MnrLr39YD1xdn1FfdZIYZhN3avhcsLlFxye2UBbgLPFI9yKSCn
j0UqQ3rpJTbNDSpRYF6NOD/1IfiI5MHq4IPpkX4Ft4dGfT0zS8VoMlWn07S6bvK6PdQdOcEM2ZLm
+vx8LzISGzyE9iDHzLBr9fXPNFlSdFXAiYRYbY4PaDAPjE5ztTd/zb1B7Y8qcYqDOKpdHP55yZax
0kPcUXWF2p7TK6IEaHCBBGit8vesmSZ9vD/EbV6Zt7obGVeGsQaOkJqyuGzkuuuwZcbHJ8QFPNaN
wNoUVc1Z2vlKpO4humTulj8xEMl0C6/g7Ldu3ZrE0vCpLSKqJuxY8wV+rVEl7TOMn/Sa1LcYonSc
tZbdnfltt7vfLOd8S06AWeS7o8rp3A5CbnIdYpV+Atat5VbRN8ICWXE0J6kWS4OP95PDY1ORHck0
0OxQZLLU8/UyeyeVxNKD4lPknFmgKZzBRVLQpPsxuwVlnuit429zb6+pRdlE1Kat/y+3zQTHr2VN
+gzKySEufyn+UuU6S1v4hwGw6S0aYWP4xix5/rVoG+UQXU+LwD6sa4EA+VKwcj0oT2NMv83CGbr9
WDNbLosc5nZQwzKwQolDzQ86G+rxFSPRtbBuksr95WvYcTN34JKLXHQ//r76SLHFlj7I+lsoA/b+
prZDjiyuHxdvGDaleBxv45YpPsOq6f0HSRaePiFug5bcYT7IU4SNzeWhwx2w1Mv+Q3oL3qh2WtGb
WnAFPBNufeb6TjHsUKHTGTLQoAbg51NQ8TN2AexWXqZ4OTNW1tmSNKU9DYLZotusu9GSAi2Fu2th
7HgchHuSaB5fLVon/EVHPC7u8YQbVHcwTaURIVmxt4upS5QEaXlfHBCXY2voAfY30sHwehZfhG2u
IERzOJV4G7174MERXeQsmxfrKj1vR1P1afCjOQK21WhTnOgTsGGhvuU/1RsS9M3836V/4atF3Rpn
nVlEbDokjiH48UYeMCPveQ8UrXS9wGCCR1zIwzUxXkqYvfRNIAXGIMRJJ4PBqx1yVeOxHFnoYX9p
GxDNMMT8EW+MwQM7zUTqzPk1eudMRMvmvd7GDx0pj8/ONJ4227G1Q3A7goVIWlfNb45x6ssEVvQR
DP1CirSlu5ustRfU18acM7iUFFcABYE4fIEUM6+GKvDTGcB8bfwR1KQFgs6sYw4WVxYuDSn2ePSw
tUSlOy5TGG4072wiOqq6wWskqQCoxybSHBL+Q4SdKJwTj6Afo80avO4izWQcB+PXRvSo5hFo/yt5
bfRCuGULJNfpMm8MuLQJEqXkuA24OGMJCFvBw+Nwe6VYkVvtDFDkzbu00mof6mO+NH4BDL+ZFLKv
+Qa7LY2P4uJWRKzKttwf9Kodj4xzMKOPC+1GmYMyAShsrDh4aQFh1oglf6fKQcFDixuGjuxLPLst
lffS1CcAJzBmdFL5Xrqv215JLa8dTRZZm3WMeFfkqhS20P8uyyCAyL3S4MGcPnFh2WCt8Kol1waO
ZayKdn/jIblnxJnCwXmNinLQaeSTz2pHdO8h5RcosNmUxV4Q521JuD0Z3T3Zh9KtMRFDg7CVu2Pv
QFD/2Bvv47JE7+sNcLmgLe4KeYGeC+7yOFVP8tW2BOjmFoAlfHFpIH+4phvQFByMZMiFxgpEvohF
mC4z/47MBDGa+gGvB1HOBPFuQOg2YCvdV1h3flzhAEbnULR9Vf+/g6uw1Q+uPkgSw2fwjqhggTh2
IeIV9KVIMQp4YCbbvp/8prJzbkfmRVWNKk0BYcWMPjZ+STQGQHMYxGAMhcszOCWu7u0M34b2AlQR
XiCi6tHk7gPyfJ2d9aohVQoh8onJ0TrngJ0uxh1mCU/QjrGO8DK3Bx3t+SPX/Jp2BKm/INKWLbrj
yl+SvRqRV9Pm3WmgcfTJ9Lw4GXVcZbSVoORTgm/FxkBsaag3jHTU7hhMOwTXjT1v477JT1Y3aIDn
PNnOtwY7oV2Kbxwi0JXEfNelyBKvwvsvI8hC2YUx5v48KVSGfMkkgUS44m8Kv7CS1M55xB7/YUW7
5zicAbKD0ckyPcko3vIXT55fBoSAce3CvmXh+la8FMy+ZlIMyd196d0BfbtYbk/dx9HKrJGcMZvj
+VZhSvW7+V9MP/EbH5Ln7ejFDDqnkX5LRgZc8AmnWENvUoQIby4tME2ic1BsqQo4e1gBGjf7mKm7
RvkrXc1tTeHS/bX0Iyex/lRUZMtAvUqxLU6CnKmxZaZ1swIhdNSD8s7STkexvlxl4n6xjcsgvNnN
TOT74xsntWt6C8TdpJJ2z7BbVcZN1NF8DlQCHWb2qgaTxfXZsGf5C88AJcnHqcT9rLHNJQzFvSDC
0nY/z1XIzoqWYIRqA2GsnPGU34qhi0To8PVnMy3kbbyJhf6GwT9/a8cZx3IKrAvfZ1Fky4t0423v
N8EpmfYR4XBMvq06J2tf133cOZpaMX/IMzLelFTPUTCxqxXGoasVi6R7dlRWaVr3cWP7/QgQIYKU
zLfm3lDtXOvf/X7Rg33VyaH8tD28Et8DwAFt15rk0oci0sd5Us0ntsuBq+u8cdgTtn54bGp6HU00
6HSWbw2JGSaM30JCywBzFGH4J5mxz7N468eaSnaqnOYn2UZKxBKdfDbUjR3zYYb34Bkwe/W53xof
tGXvRwYl1q9oaxHWLgIu0me5UdFj1jUv+ow+vgUXV72iZX3hmO7EBL5XObMgVMWnYP/PfgnxcmMt
5v71CLfwsTlg9MCGht9sI7wtwBRno/Ib/8xHEHJqzjqcpOetz2PNI20sNbAFMjj0dIpm0YgXHg1s
8v0vZeOKa5YIy4QWmMmJMSadJpCPBcFPtjmbUWhCwz9QhtgpV6GkX6gjCcWab+Eh5XwoGED0gg9N
wGyWbUaShWJxIO8aofiAKsSGwp2/FrMAwI8Dw7bZfHvaN01qbsFocELLSzRYKDbJG/maBvj+T2f0
FdKGCLkhemDef2xUiW5NpwNGmh3b91FcpsMbSUQ8zJ9e6M9xmJMibrewvV+XQU5M85t/6OeBbqtZ
i+m1Cgo/xrn2KGfPFQztvKJCPCnNSIVHjZmqIIX3De+CFsoKyBCgu0HA5jDQTprf+Vn9/ywcJigF
8b0MfB30ti65AOzp0Rz7pmX4TAnCssuawin5GJdHb8st8oYWonB2pI0awee5pzZ6fV0rvBSyZKfG
kS+qoPGlpk72HuAQkdmycZ1mo4YbyTNATS2ZaK58lLsLZ03+6edpfTMiNGRLp6Hxu5ZMwHEahsfQ
wNR/mw0OgiWl99yghZTG6RDrMAe2OOhmMeEq9c9HDDgJGYCsowA19rIgDnlIxK7OTwRLg3SCHnJt
NbEgZdWvoNI1yORPVW6D9CMYPMhLoRRocGrLekRqs9yekIn9BeLALKx49JJANCedOWXXuldF0t/b
MIY/KXj7hs5ckDew/rtp55ZY+SQkOj5qZsdXVay5FeNuNWZXBzpz3Jrc2nLyjiu/Ka0Yjj/Xs82u
gdDOHvmg7CRG7XeuqsAiP1QnD4a7b8ncP3sqJRChH3+RxOCeF6c/vzhulFSomd85UIkyvt73pnZ2
7bngXi25s9CMfzWZQF6Eiu57SvS2Xzs4gLIkyVUTxEoddX7iYx/MSX8+MZF5xE25rlt9kLas968l
/32aSUTk9jg26aXzzjInejAsIXJOWFBG/MKAQ3MRdbIgfR3ydxMi3jHSq70SGaAlfqQnAC+lYllB
dYaGKqcpf+D5u5cym2VvyKcLwWDavI8lqlAiV4oacQFIkaGZeYwcoPBiG7iNZ9ik/4R9vhRz8tiL
RelKuTAYRrmteiw0lgO8W67WE+65FebvCz8Bcn9nG51pfZOdXSjjI9veMQpiz50Ygq4ht4pC7AO7
4x/bBR9Q/ZvMQ26fyCDhecIzpQm1LSgRCRHx4VRO3ODVsGnsAUOi0H0NPuHv2CCJX8xF77p3aNAV
JLzAYWgRpGkk9iEMukbjjIVAUbqvubCtn68HRukMXfs+IcPjdtZ1+O8cXAcTwnD1BaSjF0X3GXjs
j34B5uFsy0w03PNQibeZvj+qk3Ai8h35+IN56uGbgwZ76N1rx9pM/HhjlIUqeR4Qqe7+i1uvEg6O
Gm7NGANizd/YoUJVCSxKCLetD5hZWIXQ+S6WF2T0HKTPtMbzjn30tkD/t7pTRTBS9pMWuR8Ta8F5
P6CogGHL8FgPoTRpipp6RnLmfYWTebq5HTRP0NpzCCRGQef3DDX80oCQ/SMxktMEvY5EL+4U0Oj2
GL33ydRmIA4ccfVVr8ublhm26WNTUsJYwo/Mzao2VsFDqY4bUDTAZvkvb9umzhuAK013kRIWjRED
62NNszKMh3J9aPunDdez32/VZ+W26dwzfCvnRYMZFBzzSosnf4T3F39UqwewwHMtcKfDNLor6ylR
TjLdJmqqEz6Xd21kQeJ+0SpBXdHu56hmlMUIdBkqJoyCEUsZ5A7hJ8kJV3sJYFCIkL6JtmbeSCT6
x+cnQ24fIsFIsp9c5FHrmXTcQyGC7uLsqQ8LXnWdkZFT9s2nrXgLG2xfJ9TbwjlYfyR6WZnKnYP/
m731GkX1WZc+Gdy2YslEzlTdGH6evwDYR+YK26tzPhuJ73MGMiEua/PKTcLpz2PhAu8b2lH75nFz
dCJqRfGgVun7LLzzLEjpP5pjBJ8xS9vAZLUU8sc5p75ZKabuDh1qS9O6gwJwSrk06SWnmJOnSVLF
0EQAvxTDIe0DrOjv8hhCFsVFh8sPaGUEdbFEMJXSREyr8YkhAdeP3vl40WHYkvpUSZ66ozi5WPie
AJggLPUJSODsqxjjf3cKn6OB9OFObt0jo8TlW0p+bt6zES+73tcPh5PgvK6X4owMmFNYEfyepZqO
ADuNKnQwonVz6jMLfF5QnuDo7Qp9ORZi6L8ge81m8SHsc/Q6ZjpKSfmbIYQzGytoW38ZjUUoaHaR
nVUdnpDgsDiOMbf8y7nmQgUmx5iBAVUbiYN4o+BVFybvR0MzhDqx+L+4x5FRcM+I1JkkWb7ES3YV
GcXT0fmdEKZSChqgoKSGOT6qYOg5w0sDWde8nfFz5Bd+gSLHNufn/htpFvrmG8IEOAw51AvDGdQW
0rBekQIkY3OoF4k9I/K1jdaAmSfcj5rBvHOKMhXZUQU58tfN97+E5l7/LieREr/UANEzpKn2lolW
MMK5Mq00L5pX7e+lJ1uAZ0FRe4vpIzDqpDLi7e0OQE8tworsZBLtsAcQ3TKMEY59HYO2AJLAM3Ts
+augewsOzeKnm2LpbQylOsKKFMvDJMmQiXM6yNK4fVAEFaLrP0h/4fUEInbvSlnYJbMBNRrhSJ9m
aTXL5CQmeUqdxqJG5g4VnN7CEXutWpkxf2An8xYQnD2N0k3a2scU+tjQvr7bcIPPr+sAH1nev2b+
xz7ZPOcOuyE1FiPBzl7O/GFeaW7HgqmI1u8OnTQF6IkHevLvZffqE7Hpkea4Lv7rlQ7v4YcshMaL
a/As5ysoNG5HfpOV67tQ5n/+ecEPeblQGpbbaEafkfM0TbLpLuKveb/6onMet8eGsP6dx+HYY2QK
S/chIJJQwhB9jSIZC/k/qGDqFnRdiVLpoAqw5XGE3/H9B5wiQTpM9P7AVPL4WsTnk+NkG1Q/yQNU
6IlTzWi0V+10txkP8bggaR+60d6DH+jcKFNp+J8kuEZuhVjN2etjZ++yq/g5hcD0nlfYTZEV0+b0
05VRgxgHO8fx47JdWIzAolA9R/i3VFDQeuTg7TUzkkvLhA1M9PssAOF7OZvzo6JR7vAtJ8V71pxs
kvqU8AHGaUi/0tHbyF7XKOWyVGxUheOHaejnLZcka0pPe17f69cH0D2yYZFK19mvhIF3pG7R5lup
oqT0IYdUIU8yQIdAYQkj3r12D2u5ROXxJXIvpQSIJN90FJa8BAzkMsmhNd6VSnoz9o5MjJcYJZJ0
vGOItL4lylDMVfIELJgjfh5OxsJ+C6GNOopruJP9zIjPrZ9kM0HO3KJHPEcuEQHUVf3YIrVnSng7
PU4p5Ztmq13654n/K/GVssCishpkHpL6jvVEO/zQvtXIQNvWvh3/Ce5DK1VrNKR4D7lBJB6mTRgv
l0aCya+9oyeBl5KErURJgX2DW1J97wpA4YLhwQlTn0il/7xPEtaNjoTaRl0O85p8vI2e3uDWG4Eh
Sk/yX2ePF2w0rPzzPwrPbxl0+6RGMpgXKS7JAZt9tfbhpHxL8HC+ZDAgb6mW7hAJ9RR8vRvcO0dm
FJ2A1zWh+OJSRwPvS8lHJrngbQkM/SCVUsZJDFvSe6gb/JL07vAZddsD45EIM3I+O2GxkagwQRHv
+hn9BVw634VVWr59aEYqvwlUS0aeLBI78J8/4DxlZqqH5TAPLW/BwCT/9j6wT6qoj88pn13rifFc
xJlz+dapSxYd13ecRwEmvLRT/jON3us2aryYIag4Qlpm/DP+vjnzntAXCXH1ZHZJeXGbSNmQLH6A
6DIZgyZK/XgSX5KCSTSb4WYJK+ADu3LOcIGhG2KhKIsQpmxrwXQZIqUEMItnf98WepAkbaHszU1G
QeNA20XyHlM85xRf686EPYFNHO+mLHP7JVq0BvFHDLK6r2Xr1nE/BuUDsdQVT29cV7qAjENCNtJQ
4uawk+Rod1xb2C2EaNO7yGprJLFZNjVNuSdo5ovYDLh0fMu4VoscaKZVQrt5pZzksfBaWn+BPykS
3kNYz7SQoT9Le/byawUTmXYLIZexA80wOd2T+ynbBr57LkZp0X+N2FoY1EI8JQ8GcFTpaBGl+3oS
5k5OIJ4wlm8/xrb9Xsj/ApiCtyJ0tnJr3BLfJ/VWwqyfU37Ku6xld80fTeH5xnCUBYhGyN2ixLfR
7XEB90s8rhcbEn6jVnJM3iTn0NItnkvI6dATa9VhEJydDovJNFOuIdo592m/DjU5UmGUVZ+/ZLVa
EG6K+O//CHWdAcu/lrDbxUuHNfht3dvAn8dDglSGg2KY8690vXSEiHvqkVmqdDc8gLcurN6r3f2t
mbFCoXUAQIs0LOH7JwhWIUUe5807g8rLEVEod65CECVAzOKMAiRufpl9aA1SZbvkDHA0JD4/l7s6
00kzcAYZKt+zx45goj2Q0D620+XV5G8U8ijoWMjTXXIwukDVJRitseBwbDSrzJpUyfxx97uCFy3X
Y2kgoao8rd4L4oeLYyCvwTtgk/ph6O6ouwpUoF45Q04Fa9WYVwTogm/SqL8s5d2YtE3DO0HK6SES
i6EFOfuuCIKkkcVfsF0oB9yE4OcjF5oSnfVpIQVPZ5XYBqGEz+FBZ9LiYZ4HUlNwGeH4s+54ko2G
cXEyTNVZFk781egHASlJAEbIemwL2Z/NCLpMIOfKP7vrRBHXhjqQbVIXLhoaFeWvtpsBGGcWLdBk
L2Qzrvhn0S+W1aLI4jMMx5QikO6M+tnDFau0or4meTY/uw7PcXqMvZ+1+XuxOuR+s62s386nGnVX
1/5FDCpmFEm1sG+7sV98TsWbp3jwVR3gZbZ1fGYxciTNMHBzVxpdU7Ai1s327SVKXHHx/Dm2wgpx
HRNg9xs0Hy1qsgPhG/La6EAAiKSVoV1GJXMwUKFz2j+R2EoGQwRJAQXi6pSCBDZTUTI2S5vYVQwx
ZfA4vW9pFdA5wTTkjS4UTKtxLTXYFfmamS8R+BL02c+q/mqdw9JRw858x+QrREceJO6JKLQz/zDE
fBcFwG2WHWMJL3puiBWqixy5UTzyPpnOBjhevcMwmxa9Z+zxrn5Q8cXzlzQ2Y8PNXGPg9Phx0sLz
zz97YJ+4MF8cBzkvZhuhv0lLCNEYcCpD9Y3iGbaDx5vpy+FsKOS63Rqd8AFJmc6r/RROoD91FKS6
5rHuDT6RomOwmtvgg1hCToK23sBYEvGFdWvyvXF9jkISp7BJKLLevwOO7HPgJuF2cNaeI82nHSAW
ezxLPPeNwN1NZCPVQBKf3E6vlNRLv03EkGeiciwxTSJ5UsXdNswrV7qRq4PpPy+yGkJvtY8Inx1C
tWgsWxFwZg8j6ZupsFmoHqSL3xrJyP8daTv0rkrr9tEfR36RhYA3bxAqDCcIILNWfn/rAFB8MBSB
6XBOR9RzABXSPEpolchnN/iIJbuAaHM65mELCeVkuY/dFFhBiT9YXWlCprRpW0jaBvgOQu5w0xOv
A/osV6UJ936LVqe8oXFwSNpKSVR4I7kU5oUa5LkPEdjKy/SJ36+S3Ea0NDHpoJccfhN9wRxFQfx2
5sXaWWkWs9h6pjsICQG4RH2QZisLqoTeoGivUl+P/dPsbx5VpQpt8bQblPHIYZIbt1/JHk6Px2tp
2mMKfdyBwEsOc/fAin4C/BMrDChUzvw50Qe+oWjiPhiop0ZkzjENWUmkmTglO9Ocli10BHjgPMw2
7/pP94MP6+CPzZWe1y3f1qx03WxDcBX3VdbdfwJdG0sOZNs4P7HHhHqn+ljDWuI/S8eY7Fjs2BcY
JE2+CgtnuDhrYR0VKYVddCeY8PjzFT3SuP7UcOzgKkMbsYZT4TTXGbHlfdg+l3GpjZ/yL1FIx0OX
bvZkcz97uTFJjzaE0s2cxd7KDnXMhOLpqfg+Ue0S/hn9s6Zkgo3ggea9JpOMdvqOo+xKheis+haH
XptWwSmcYxNrqfKBdXTW8AJFDz7Duz61cguoHQqoa3i05GenQKQOqhQQKLI4eJBDSCTcNemCvRU6
IgugLNxXxQxNRKkinr8ltZqcz2GJ7riyJcIpatFBz/Zqcrhna49KqVNRTAwphPlFbFLbpkJLTFaG
1ew3P/7StalR8qX8Uo54l9TWetTdVNMEGCDBXCoRy1Y40QFSsW2Fr/1YbV1n9R8l82QrOuBFA9vK
NnjTeFk/iAmEQMrYpF4Jp9NJBXGuQPCbqcK8Ees87zlCMH3RW3483ZJYhksgjIKGuSt8O6d/WuMr
MTlz5341Uzm4ifwO5He2IOhkInQiVtQY5hQdr0NKG2uf07mLZd3rS00Qz3NXvF7UynZl/yS7gBjC
pB+3NEWxd78fuBeyszAGCQ0lnXgG1yflhjv/+6pZbVzFDMWEXk0qwmXbVnJCx0BP08UXNgk8IcTB
iQ9V1uAAD8gP8jum1SwVPr9qKdBWgnsI7Gv9VumfmrnreEtUSsZ2tFpReLrLB0F25tpXfPu3zFhD
TeQ24frgDIJY+wS8Q4PJ/JBFEW8hlMTWtTSU0U0YY72sbx6K6/l9ITqb2uTdvXEi5kLrcZZSyEyg
DTuo6GJ7RTZ7hFK3YjQMq0BzYulS6P6RLDQXIgPU51zQaqqD09zNYchlK8ZH+GqR2iXc2Ur0uooH
yvIF32O/JWVsbeqLtFcUiOFY94jshXM6RdGrU7ZRq4EDcUoh8DGeenTiDBiGLVu2gToqIqzYZQvh
Bx92+HUCGUtpbRvW+V9oQd2No/asMENLJVa9e5wvBHNI6c5F6dIO7zzoLXQLlunAR3fD6VMQX9rb
m/q8jic7UA8FqPVUwMWC0fnIsnJ4FAk2CcqL79qBau7OpIpryq8Iosw41CLhSObTyyKvQIy08QOD
f6AV2Vmgsqt5fRD20QcnYs17DqlFqyjQWzoNJ9eqWAv/VIMDaNJ5I/ZjYo9Xri7xnUA/the8t6uS
ivGJT7UNlX/qKS0tluS86kb+NcKmlkte8LFUQOEHiXmOukjXroXsj+hy5LeEDR6wL7DPlUPWUEY9
e5avEjNT1uIwWfC8oYmC/K+mRB7y4ocKwPnakvrDqCDd1bJVYLPiiRMXJNgIT258qtixUfTOpHqC
awOg2VikUm/s3pqsEb+4nISNDb5GspuDTpn33p5fCT816MCRs3WB+XwYIEOL7U4zN3XCqQmwiREP
5W3evtwBngfHaYFE+QtlvbV0mu2FlkJ9TkEm0JLNdQRQnyYCTK5sfcbPRtKQkLAb1zEspphXWgRF
7m52FY6uH66z13asD/KmLGX+AQelVAvS+8crwOll1zgoyvG9y22Py9MIUzc56Ul5UrIEGLOCYlMX
eWYfklopXjJ6HwQtviWyPXTt0BGPLRQeo2FOkn9Dst5jAZDCxTOePOKubmnDJDt9C20iln01HSh0
TV964HBAURrfJeAIQasxIGOsOfB6gWoc2S4vKdA6y50IcHD465S6KkHhftAZ7zlMAD4EbJt+tk3p
a9Va3r/Am6ZIzAhGZYanIg9jiBC0upjK5yQEZcDa4ztHpQg3c3lHohtPUoPZ3kfAU1gFgGWk41Fz
qBIJFtNpoCxRwu/LUhJw3psZWN/ygNQ46qBrwySuH52U8u3DNYcZ3seq9nc9eAIdKSpN9B8ru4Cq
s39RGoHPWJ/VC9zpqJD8WLN4hOV9H3UxeJTLkXu/E73BpqODNj4kmbtELnCGB6M1DCLWanRglE54
LhGjo7fOLMdFUa4p0Xh07O1nEzaNM3fIseMNnxwPctZ0grYT0tQY2Mne3fkgwelZdHicQsREsxzr
Q9AxMYP7tqG7UMo1X5iN+cJMCDhTiiwnPBQVWmwDdoludBPM1CAaPsEdlH5kIG0+TR1qfKcF+yTM
J80vxWpckdtRcaeNU1tI+78KGiL0Py6QmHXRk2sAogxT8Ygg9s7FkxfKB3y1cSTgTP2ip6amxbGT
LsXRL8pGWQ/w8/FnhRpXt/9ftfrkVDDca3h+yHoIicW1i+UIxw/oVxiehZbIWp3NoMn6+k9rO43R
OPkxSuPfnUG/hM85nVboOiI8SqWGkoQUrNAwKoF/yYJwDTXfEEJpPYdmI7OeOqNcO8re8ELw5pQZ
NUAtlblKc0YCf/1PKrgzX2rtD2qpe8T9WNrOpKETATRSX3ysVQtepY3wyhJdfs0Pn3HCF+w1ri9e
lnj2gb5qAFd7N9LWYO89HYLRNKFYEq37LZcht2jImev0k7A9ApOKaPto3n7qxtiBZrZ+tXYNCeKh
yH+dhG59rmsmyuqo9nH0BTOlLpoWdDkzHlu49vrAFpbmKxCSjW9M8YSkoKMH8uO+pVl/hpCNELoM
rKOxKCZRuZBmOEK5nZ6+zTDxm9cccBk+AOqCv/JJtJdiUuBtAtkUPln6PCBRFfuh9PCndmdc0dz/
pOQNFH6ozEY/Uh3Wbpdf/RXMjcKbm0/qIoFmjokqWwbME8Hgd0nFtEglWUv2DBhBIUIEdrWOuVcn
KNS9NW+7fZV8zhdpaGj1l6W3BcM3nkUrQbzcW1F9hwDvrt2gyKn2KoL7s3tGGXWxxHr577kRWafF
pe9fF6AClucMLACqbof6M8J/11E/wG8TwJg06cg2LCV3AswVSXyNMETZ4F/PR5xUAOFW62pmu5vp
YzXlTHphZ+VXeGA0bO+9kfdIfHWTSySYvIn0783dMXqwbSpjKh92q/yDcDonyv1MZYZIMX9RZyaj
3GcIcqvBkj15GM7QmLzbja+xdaf3+WilVMy8DVMxL3sHgHN3JyjKKsm5Qbl3S0E6PoDodbSnT2cB
4lV+woPjUzdh3nj5PA2Nz2kP2ZU8Y8lGukjH6hCfQKe5WiX/v8RMu2f26CLICS7F6V9z5PMVxd/S
zYb6xBz75rG5qN7ySd5mVxxrs7ymyIcaqixecai4xhVfvGR2AV6G220+u+GDloRexZXy2fNR8Xpo
qSuShnHHncJ6PgLuPKmWzyRlhzOtBz1TNW00YUR0aqd0lBlPq1OfiX05MsPFyHVV4Hn1UZwcV1Ew
BKi6kdZAP5PJQWWy5trMqkW0sbsIhHQcs8lCteHSWynHBQf1CzsoIsV6QEqBL2vR1fhTLJhPFOon
iIiGVpdOUUyvaK/7OCXMqw4eu7Hb9KDhXGta70j4zTcbrrA2FMVVaRbBKc/FgY404W27UuaQ7X/R
5kJ/K1acr2iCal1adwY6B0XyYNUZPgQJn3k8L9OTe8Ax+WHyO8QwNAEJyceEuIiF/oHCg5C8AGh0
2UFRlJ61V8tLeKzuKH7zGWuchzw8Iu9v0ym1yOcSKotu+wyq2H6xurlkVKu5XGgnLTINwY2RENsR
ujTyiEGBGR8kU+OOUCPpjurg0mUe382AZuuMzHaMm4VyBeW262Tv10T2VgVk2N5PCXFGzSVNDnkg
0S2Q0apIRZRGwIswoygdYJvgqc9AAjc/y9Ues2ljAkcD64EAFG7Mz87ExqsDDhSvySjYJZKHDCOg
T/XB+n3fEjSzjrenaOhkt+qcHHgTcx5rzzHlZj/SN3Prfs5JH7bo0R3ZjtOgaSW4vMPdAHY6ltox
Fyt0m+opkiF1xGe2x+8Cjs9Qr0rfV6O9kxWwK76V3XsKR049YtTXbGX0IW66u1F8eTFXBTK+mifR
j5wQ+7Ahf6DJCw7F4N99JcbnJETeL4QYQ4WoAoxiBUQHzOI+I7NkT/7zBULpGjyhsnGDOpyu1whC
ei8jNTpXI2IRzmOfHLPFwkp6VWzeIKirLSQdHpdbqWTGcvxmgHjxpw66vTBNtD8kHHgETdpHCnWx
A3+47G+N7VT3FzVcv0T9/IwkXI8Pp9LbuiBurPyke8dEmySIxymNS9CWeFmfJFkjALKS5GZnN3Pv
9oPaI9v1MFgi36M862t/gklofncfah1KUL91gP+ia2T0KD3lW5pMxwVswwqWrKyUQbuafpcks/YQ
+IBYd3cPrWtQQURv+XtVn+FIk7H0WP6NgT955nVi9jWiffslLLvhv734dmG3LSvvkX/GemsCc+JU
KnMWmgcRR6UNqoHtFAxVWONPVH9MBderJ4SzJnJ9dDMm7+FHIZqRdA+NYsyb1ZKGcJd9hix4f7tm
WsQvl4mVuZdecxlhm8lq5+Z9ILyQRkJJtGaINSMcS+S1yscBviL8lIObOwnTf5fzLfpHcM17/i02
S6ONuONw/KiupF1qyo942DPO+zYO5IUjrFptavRIiEogkYqX2AOTPK7J8HAe6Igh27t3Ww4rU7c8
P/gdq86zKCuJPkI2+sbjL2TfUw6st1lMtUTob1t6arCGlF6PHhHiJb1+i6mc1VBdw9ezdzJHyanh
NKApsrpKPuKy2gZIAvM84seN/sLXP6nfDBn85jHhRBG0VlKC0rgDweDBg4rKmFHD55UdiSNA5m/F
0VYi7emjq37z2RJh7S7joticj6h4eBnFVoJCQDX1LqbyTLiu0nA9uUpmCgOAGF9Jw0R3njxBGpwY
i0IK9IJB54MU6tmV6iDh3+ek/9O5IsqpAw3JFsPimPEQQKbCgAvqrAmCEPTpHnrAVzaPgzpLeCyZ
Pw+KXrQWCsPL1f9mcr5rNXVWeGx01b29Zk2lEbGFjr7TWDsca9sEz9uOI9DKu81mmtM/MPPdCh7r
zAJRvOYLfs/6EiSPEQ5Qgm0W7oZ7zOXXX/b6lFYiJKukX2ktDyLM4WCU623AJFliOekJujdqkWSs
cxGNxOUgOCidDuTISnjR42rhQtFypzvLdNlk6eru5fvwSMABdt/Hslt1dhfhy7kgqrvpZ2X3YSZc
UwAgSfB913cG6IV8rmI1FhgmCg/yGkVd+Jevov19nTxGafeDk0qidowJyT5LeGnryBLfCUe65GDl
lElMQhpw9hejwQLEF74XPJGcWPOc46XmR80b6qRlXkmkwHeDz+iw0wFxGaRHdSt4kwvoIfK/27My
y38cmJGunFYqiGVXlNxspsJ7vcRxo2r6feJTG9lPHH3QeKXl3s8CCMOyEAFBbO8zoYI3kDw31R7q
4uT7F8mDIPeMz/GWegDNT27ZgP/QIvPARm8dB8Uk4HlYKX50GbqIPWzfOzjxdf59Mr9NJNdwZqVY
hQ81ApXLs9r7YmDHbUUD9GBQTeU9QujCR3IwaMMuJSBDFSaJWMLk77w8gt63n3zjff4PabqcRaEQ
6VuXed6iIhGh4Pz0HOhOatsvnE7VYim8qfwdwfUhUfg5HhFC+NN+v7V4fstfk4+t0jYWbGUm5Nke
SKqRZX9Y3RejxqXrc6H+YnLtmz9cPXPGiZu4xtsCsZZ4qJnUHfQRitfFf5wUvhftXzeFX9PzI54B
yZ6mCTrTghcpEhQco5bdk0dq3gDNwye4xby4GVcA7FMkOt7AyXzP7ZKui8Ofe6G4AEapa4yIWtmR
eUWDkfyyc4ZC09Sl1l1LP6yuAp5hyBbBbaaHfjtNEzSIIgvaGhtPDt89VZEGdVdOTY335P/BRPJu
jnQ+VbwJqJETJmpqSLuZe/N3sisfEouj38WxNrMHKQGjM7BNv9qHHZmWQHB8gqJlzHs4oJvIrK2J
WD8aAQ6pBRukQKvLRpXXe7zJ9bUubRIp0eN6K9xRbVKqmsIFGZdvVmxBTQ8MykcNnwsJ78LllOg8
unh8/DSmc62g+BYJnQZM8eNlrGAl7Ce7RciTrV5x7g7WjZddP+v1wAKhiG9eS9aadNBAx2DG3BLT
p+RA8huBd3ngsXROXYiIX2hE3RL1Ci2g5nlJ7bmnMZpgvgxblIMEQeLODzOalSRp3ju+nGOFnL7z
l6Z89La6qhA2QTggu+9rxS5QpBq8NKyOVESNKY1fc8aJOH0OLHgrhLrQ5BrmxuRbCGC0gyS4ryp+
yT5dPI/5uIVyRYokKxtCPG7GEjLsYD3rZGl7KWU3FloFivMgfqphxMeX/zLzZ4yZS6wE8V6s7OnX
EDgMHFoUJOE0TESCADZFKx4EwN7WozRh/fQYfjz+xyPBM9FAFKcpWIu56LchJ5Z1DLcRQEhouy7m
E30YV56R70GYlPZVxdRozpgyYX7VV5uWtYHfYxEPtzMxyu92Wvu8b/Ng4OrfK3iQ4z9T5I0O+H19
V6cDrajnHD5JRdUmQhccnEpFE5nSoH8wmE3L8jzewY1d7jgNXlWkzkR0PcbrnNaI+Npn71BjFiCW
sGp+31tvejMXTWjghv8TnX5geiZGq6zHEOghoZ/wJvlYeerQMaan6QA4//CQBRlMhzrsBkXOB2KG
thtzf3qlLgAn5jnKSO9aqVxoSxJP8hVMgCYse1hX6dTTggalFV3U3V4c4WZuO1YlTiZnRTTaZTMt
GWlZQhmDmkwUCjxzLbbAI/KF+VS9Zvkn/d79RITm4J+hUng9tEoUZGOahrmixAvW6bn6bj2TvMq8
WDNwwqY01pa7jhxLH4qCxYt4omWe4c7ZhQFoQzohT/3AP3qsPj8fLSV3WTZ+uPjBmIhvWR2DAR2D
6ntGlf/qrtqaIOAO8z+phzQqN8YFUu/Zamvc8FyYBEEqnHKQAdV5WWGc/LiGhhaFIUrYO7w5hAm/
arxHA32J6SXZZ2ZZoyj3wVN2yCXE7r+b03n6lKfMSl63t9FmcCj9Dofcym/Bt6NkYNasmvpfsT2E
h7PqHUx0thH4eBMaletkmVD5bxYHL8EB7DP3+C/et/W26kVGJdOy3xoKo/DLECEXZp9UsdW0ll88
HPTwsgCWiovWLQgRt1y6WCiqmbaYenCTZxFxAQzsZCgBe7O6b5bkaVEU4rapjuPXUM5zflrBfKWy
1/UJNuIJ9ctoUI4S8zDtetUKXEUhCbrdFzL3xYIHt9dZyVTfJ670Da81iMBaQEMPuxSdv3xaEuvN
Tc6G/SWqpExusVwfw2oS1FMCrXmFH67OblhoqiYD5tzhWB7tFa75pV6Sr3z1Z6sCwG/KtZ3hRdEn
iR+XaQlODByg8enCLvjIS95JNMeahdK3/7W2cJzA22ulmVJPPsDNhGimo83OcJpO+01ijimMqN43
81aN7mV5bbY9SAn2zHKqKqOqbnYV8sXyQvfx6MxzsWo22JY8RSo23Ecsuag3tqyJXwMN8n3nou78
a3HDNC99RNnB8PZpMuY5uh+i7pu03nsq0d136pH154T91VSQSZaXQuUk5DqTtI9hfX1SlxpTqeaG
5Wo3YPj8f2x+lGPsbAYYb1yeQMU4bXikmnqYfvKdJuYPm+/La7W46Xmuhh2j3EKT8ca7UxunBY8L
VVmECRP3cEMO7Lt3iqNCng9HJwdzUbX4X2a6MC/2qJo7lS3XggyVUx7YCEB8Lyp/HQSZMuvOxZHh
+xwIXISsY436hQCMPK3ICc32wUs9LJGC3sKB+alw31sTu1vS1I6oNPLHSYW9QAChVXNcDEaIsfDl
e6xlphpkBUUH3QfGwNY4t6A27zg/S0w3TkxjPVlNcST3ZZjLTLXAgpTuvtIZ/VGs/jh7uDPmM9WI
492xUDQmyk9Ljyt0y5eQvTd1/gy0JaaQuLpst+/M49GWmSeFrJp0/4REyqpaH6S11TY7iiXsWvHO
fc70nHPsv/QJozvAGg8iMjWAuTvEWbEZHNkkbDsLHD0SlzSmbWsmIcdwNgObiyQS+9nnT5x3kUUl
5hQU2I6YFyDt0cxbFOp4++qQVSeuwup08EZzxgCN7DkMooR9Jfr8tLSzoMmytR5m0DI8eka6TU9N
/WXzR9bQVW6phwBG2QHA/MdC6m4Ak7eWIf7BuGKvNFCGSSy+7SwZrDyt1I7CkH5CM2iaHNNM/JDC
6zRnCF7DRSPBsjKWyttOMv8ZBzWC7DfCsYbkhbrk+kUKdZMmbmYfE/mFDpXbOW1IcXh1MUhCj1t1
R28aicDh0PErQnRER2aaqa8ReO6V08TXAHG9aBwUSfIu+fmooS9Jsc4TOGXWeijbGOo4hIsv2/tH
UKy++SqgE3VQLXorRRsCcFd5gvbMFPJnIwX4Bq93SPkTUXzGbfIhc0FykASbBX7W07/L2Vusep2x
SoKkOHKPoFDpf5gqfsBLbx+TKUkSwgPy38CfshDWK/l3tRAv5BITjqUx9NLPioCJ8S4JqtnC8Afb
SwumKtnJJMRIrv90Qjj9bTxjYYeG7mroUON37lbgs1uq0QhOPnxoeMsANdQnBNDhchAE3NUEA5W8
6OGBQOK5LPsJgXny29ICHDh91rAK98sFwZnhyYuprE4NiRuoQBc9Wjdp+xmx2qybCsCCmjMFjWI9
FX5SHLvBAEM+m0V7asjOQQjcyM72DAyn++ilyiQXuCE/SXYFlkx5n/SPIiQE7tvKoGz6+doxGVdz
6qwMMzDpfCqsyjtKh1ce7a/rI0YmgvQDsc519xvRX/WJ0WpPAaML3TZ+jOoy41T3Dx/6SYSvLDOl
4qPfPBieRW8xTofGVW52x7hM3x6G8QvcRumEA9y2sxDHF5PyxQjmZmmI72wZz+kIegdHlyfNys8F
xj/P9FBA3PphmwBGnlznZ8cKQdpj32MsBQs/eOo0DgGiaEB1mmWzWXlLQ59eXGFrgcSR2bnkiwgN
/RllpdK1mdRg5HpZ2RUf3fCR0bzLuFaQvQ/Bjmfq3M4M3EwuRSTZZ6S6Kwl78zb9LHU/BPNwi7yR
sNJh/pMt/XDUpXx1B9eLHlZxBCbv/ULthz6cCcRs8tho2ryS9KjzTEdrHEuSRCXouonD9UlWeHD2
glChm9CR8d5oZqHa92dFl9tgjtsy/o/Nm+7du8RpdYyPL8tcfTPlNJYFgWSzQRP+Jat6yvT2KCvI
c8E397lN9jEQlpdhcuWCp84Y5vIutqBLq3xUUqDVPKFOhxfA1S6wqQJ8kvjswhpG0dfeM9gRtQXP
knddjvFlyr2MlDzXDqxjmUEwFIAwvO+/lr4xuC04ehJ4wKHihtFCgfbzXZXMsaIvUrv35s5i5BJP
7ByhE4qacsAIcToJPQEbzVyaTbTy2pQoe/00sx0HuxryzwZ58XOijM9TP9qwCjCT8Hu6v4wqIYDe
8slbB32qu+iRTtWZmxRsRyomOw5+KHLYwpNHmgwk1pc05s6eLehaFxC2YkihEUQGlTwJp/N4G/T6
iAZKXA7JqRPZ/Ool0oOUhKlqCzcr0E/eVaS+rftFS4XBv62GV4CfwdBxvsSQ+JSb4i60SRwxZqcZ
1+qAnK+uwfbg/hsorqXgJYdE2s+ol/1sOmVWjaVufVDuSQN1aMjQYx/fzHkWV9pcBoXZGTvbUttf
63NuoYaD2N09zGzUghZR2E2zUrs3wiTzdmAuA6xYcV5eFm+LlglLbDTk+87NqPev56Lk4W9xCllU
NyLrr5Oq63FpWZ3c4/lTR7qqb1uLpQRd3OHq1DyhvU9m424Vtqs8Q0zjV8tLnbRa66Ja3LJU5sOL
KAJkPe0bFVDiKcCZZEMhkIN8/KYApmSm9L0pblT2d48KPXM0+jbIPE2iDLHV+vXRr8CtE1UrGLKa
vZM+YM991kzYkTtEXfs9xO91lVe1pc9ZNMy2Y11Iqtd5XBjam0wXwi+XVx1HMb1ceUK0GCTkuEdi
RletzUNDZxHOe+OjuQNcrJ/JQ4nzPiG4Dq6nKtncghX9IfUw+OtvuujlkdQiEhNHs43otobzG4IU
AG+qlrEn4TtGLAsj+ZsC1s20GuQ9KAEQ1/2eMwVWd0oh5UuB0xU2IxjE3yXaJUOL7E5izweENaTz
iuWGxAORVtQUGX8pA0eVts3Ikh5699rF1Y8KnkFvsawWoukcA9BD3iIMHL0tWzuyRPGvlcaQ8rRn
3IO4wYjJ1RiHPAWbBLpK1G3hHGwRzrYm+9nzwnRhJLpwXHXtST8BOESrOfHna5q7HAEac3iZyrXL
3QIATVqVBr8zK7zf1HXS1qFpTkx3vyxsuWMUveZfzksGNSHViYxxZ08uAoGnXiDdmosZrfwewUD3
TT1mhl0hbans9NDUF0MvTN5TAIKvLnUUtskM+dKQCCLHI7Hi7/8kkM6sbJia1G0qPb95W4w7QjZB
6D+0FFr193Wge9AOJZUZwmfd/Vpx+AnVmqE2lhSvrfxGPB14vLHUsYGlWJ3L3GQ7oQ5x98QS8VwK
eToMafDgcegOpDGtbHBL4+Jtyb6GLU8/3X/ftixvtO4IxNOWd1wktCbUrGC1AJ+MOW5pTnH3JJrq
DZMYJUXfcapKANAP/+QULGB/KqvztRzg/S42VvrVugkyxUk/uBFbyhxYLV2FKjj6HWjX9mpTt36Z
sU0oZaKjNCKzxvlQ+CP07+f4OqjSWElOheoapx8GNtirkWrb0x84t9x4hFwzRMlQZYAgLn8QGage
NtbJgf0ym4lmOxDQji41nvC9TPpXUdrfka8UwpRIP4O3UreyV1TnwY/1EYi08boO775eqQsYZoBG
IaBvl82mi9TV5/v1XbUTJ0cUH5p6wLtSSGk5I9Y0Ky7K7nj2zgFl7F60+BucYYg9dggQXM2mfQfR
x5Xuv6mf+cBWBjD42OqfZSgliW3iIknPk6PJBAb4xkshIuyLWo4BiugVkbel5Y57xYdnG73PBQ7b
Vjwn6dbHIz/hjNy83LurJ8ZD03lFCYqKXHDG5HcpktvxFxHXzTtLdlxIfFbUdSHPp+Reh8VMGKBw
915fngJpAR2UAGieMoDBFCfOakSA2JmS8l3NSjaD3oHaEQiq2es+UWIVQECBvrDVE1DUMZoUzh09
coM7sK0O9PTau4wtDKJJRTzSSvGc22wgFKpyuxiMOLU/JTZTSA6Kybdu0G9V7o24qPTTANmSvlYu
Cf6laMgm9sCtfvFozKVMgyjO/6Tx0/tQ7Ryb6QcWcOvfF7Ut2fq3Cwc/xRS7wvjLLtWjBZ+9W9tU
4ZEXbW8+JgAk/C4LqtC6lOsao82iOVwLyX1F5VzPS0s87aQt0mswHKW8+8rspqV63r4H9jquQXXX
Wbpze75zp2NB8UM6Q24AtWeyhv2RwmpaPnQWcL5gdrPQ+43ASvK1Pds4HAgsXY2hovuaLPoL7uED
uKlx2Uk7Y3zQh+p7PplHz6BKv4TmXMf1uq6WMQ2kjsdLhYOXHWA8XAKEpEtw4PJG4AsntD8mLz82
IU+NItDRS83JCsBF7qb+5T5k5lRe+W6ENzwI6AYeufjpiQgZn75wFevlB5hS4nzPfHuwXlHyagVJ
amTpK2UcGr066rzuI6CkQ4BTAj9qWxio0MHi4Tx6mTFDVKK20LcbxFmDhYJY+fakQ6STfcIMMr/S
1P7R8LFrHhfxWBRUltoMCADnAOXb49jsi9q56UauIBflzfIeBOmVUGNz3EobThBL1pT0vIaxr3oO
kEjl7ATHbsmzEloD3SjqRiUy7neyXMTR+G17L/YB4O4CGxQ1gpu6/2Sxd9UUAoe6/MpcunoLk0gV
eQak0Dgz9m+YtOHj8mC8dtPHkb8KupHVxkoZgKurrC5gX9Br3rRh9Hbqrslp/zDhrCBJbXOQjMYA
e4FX1lqIs/5gnEwW6ExvI9bBvVEjF3yHjHqKXuFwW2PHkoMFgqefpNekA8cHAHmoSmG8E0DMttw9
A9jbWSaotNBczR1m9zsZpmLUZzO+3HhocAcNUevDyPX2wxcfduEQxZFi/HaXGyP4lmw9Hb/g+wlz
UHa0geaBIazoQbp/yDUUm9LqUAQngCWGDHYDnTVMNX7Qy2/zix4nInIZlFwz9rtPN1m4e5Fogdq3
MEi89WcqjEmXX+qI5FL0Spwey6a06rZDBSEzA3XbC7Zxkndwa0CfLXbB+Htqo8mcEMdo4UnIbr+K
qorDvTNh6RNiwXbfPqcRZW09kE79up5YkHCnVs+KfZ4Kz+4OhsYVf0dRD3KRSc9MDIqesi5AnOqu
VBmRrxysh/ryG+GDP4uEarMEofY0p6XbXnJU7BfySotPjF0pCBENaaxTLOHnQZROyEYCZAIXA3KS
dvxllrj1fZV6HjBbiILqXwZOmbVI8LlpAt3RAAA5PS7vjnBncrHSb5F2ZSBnPH+JxPNheb+BI2s1
W94p9DX0iE0cz8kRTEHaL/JhWYgLgsk6p6eGYjEL5gllrMEUy53L3VlmkfkORcTfR7QjE0ToR+CH
DqI66nFTrD+DS20kTVkhxZIRubkjAkfKD+Efts1VdfJHMELE1oCNaeJccdmsHYyC8cgFZUlxMOnl
0vFL/8K4s5khKN0M6GDlGCTLYKAFVylsXtxugR7GHaD7Z07SXixPkF8PdhOVHHoFE2oXtiYRWmhQ
Dov4qmNfaNg0vcJFrpPkB+wMQxkx+bT05By++qL71Bltz9ESQqv68jv3DA2PcyxmhamOQPVLpAeB
UDcTVOM8a/q3MNxJ6gcnn4W85pHSKR6InUxfNeE7NBPaJ8wNbVXmRrdwS05My4nGzVXJF7lxFPat
1x4Pmcmr1MKsMYhnJlAcNsmzKQAasZ79JRFPhzevHd5soDRYG8sodNaYJjKbZjF7gx5aLrbWlUO6
SMWfMzAeFZkqLG8svg9qp3amD2ikVSP+OXr+KSkC98YTvvuMpMYIubRBAl/BpfwL7GwqPet5rEm2
BmmgRR9t9YORRT7mvltgSmqfUc7vMuN5mpWcdV0QIDk/KgYUZ5ZolQB/f7x24cqM6IDm+qb9c7cg
MA76lWPzipDISxrdnclGzWhGy0QcsGXGrbWbNa5sXGLAscZoj9gqs5V2+yKOHuhUtBMvMVyenmub
vtEKtTzZtbDuS8abwSNGtQFTasKSGHsbDesy8hYKKPZLvh/h3hmKHkYoSP+psBkhd9c6VkVCsRdp
P/0KJyT9+sMV98NIWe1cc6lU2vHwGmW5603NnBzLWkA7VYhqdoy1euTDQHiKalmZQ/pTABKapOET
SiX4VfgLuZ9CfRiM+13yaU9jwQc8YJ7lR0NW/0sSmZAdiddslImzJZ6gLqJDFBnnwryG7LE5n3w+
+3LcLWAk1zsuKvEFcyU80rB7acyNp5oWYbzIGr+Rx7znPh+rMCj1vOcmqqcBRE8k6qqS5CNxGv+h
juQP4BToVjIXRjzwxOjqgfld9TjMxQv4RMyjZs8WpYXyV6YuhgIwUeT0dumZk8VcaWSlrh5Dsy7u
+wa70L1wrCQyTggtuxlgQKuHdW8G31hm1IEm0dqF/pedBbva9XhYYO7uONEbM81kHP6u5ZcHn/CH
mXGj95eYWbo/o2Qg7WawWmwHuD4aG64u1RSh9UEjBOWdhLwidua9hazleHOQViI3nni6SO+4Q1ek
2ktYA9gj2pVaaTXrDI1Mdl6TLMfzMUnwxr9eMm3JYWY7wLZc6vbqDxQyWF8cKwu8SqmkayDWhJzH
K+594jhu+bfo11abvU9B/5Up8dQXf4/95BA1sVccsRk4W8zEKhb7wgzQ0pF/YlBoHWuuIUhv3I7r
bBwBueupYs3nt1K/90TGWpOKVS+GT7OE/lX6MlWeniM3789559VY0GRpvtzzNc7gEY/xJiADdiUV
vcS+ipl9KqWBUKsII9Kg+xEZ6MPjSrys3CuafTAdmkfTFbUoW21ZRY2O+G2SNrqTrybg7tCiphSy
Ii5x/VLKQ4cJehYBb7nEQlGpiHZbB5IrT1dUhEZIRWXAZng3B5HBQYhvp7jFbAe5CMeHM4eYcsEe
WP6xbJ/QSLociXs0IReOtJgHjEfE+K8swHOLpABLT6iUexmtRea82wMV4Ffop5hSOfvwqNAljx+n
nX51Cx0QhFJayK/IAnYiFDjAwQPMrY5drObgOuxtZkAwgkNbro4WEsJbSSPnQzHQyhOPmqE/649l
57QsW+KpzTwxSN7zifIMVcMiMI1WcTmrnpByeJ6OMx1NcCI9FNEEvCSFSllrvulozUCCWkzMjuvA
6QQCB4a/icHfI1AwDYAOhGplurSdyTtWn9PtJFUG6fNfCgvsU29492erH4+rm2xeImxZxUtzCLRI
lScyegPXvmCZscvyKO/f2FEQK+H6g/60ubQxhwQZ+UhPl8kN9rbuqH+viDrpNW8keaMwW5gL9SlP
UZVW6jfkxgwqSL2VapHJHzwXvBGAwSTEcBOS9QkAtoU0mYUs0LentC2/BsFKST8aAVtZGPTXStq+
vNWWOxomjRJr8TIq4Cc93xu9dh9HoE28tRidxtp5InMEF2ZG2lG6fYjuYW3Yv0agFbV1rrlLQ0lI
4JPKDsTq/Q37NsHdFA7LLUpezIyZ3YggvpdwwptQXzZW6RlxU2wmZNV+r8nq29GepcDcu3/o/BfP
OdzAbnI/Aqb8QNaDzoqpfSQEFsT61ha9KYsW2TRudwlGKb2qv7ScoOFHzhOD1pn0s+DbLI514JGP
Nr/uObs4F9l0MYT8K7Z3AkWVxmsL3D4s3bOFcvUsjBu4p0XvIXHv5IiEqkoj8ZzwdryNT/CzTslw
eoRBo73FxPo/L9DuyaEplg3RRYS4T69TyRj5DMrq8xZW9flYSDWWoxS+RgVgRwlJWH4SeptSNoFV
NuYX4J+GPoNC/tI1rgeLmZoP+TtYdRM0+rj60xUkNPMRzpm+gvIsGcp/sbVv6c14/9P3G4fmC12b
4U9pcWqzgDb2Woqe8PFOpEfTWbMCizZ8Q5UhX2mNkn17WdvCQcy9Yl7iw/Sh1LnFYcEDBWQVrgsO
IZnbK5ZB9t/CW3ikFNvsN89N8dWmzOqkvd8hcBah/e8//tpiXhd5wyIuOOokYrpq4j+SqWX1wMMm
Vr9qeshr7ISv5q43lu3kEBYp0uZK60h3mLB/OHS+trDAnoXkG7XC8Q76kfEPsOnKGkJtsQ9b9KOJ
yoMlpp9RXT1Q+Lsfmt/88tuquBKQTm8FnepYsD9dk2jq6M3m0O5qKRylq6+SpqfFSaPOHkjo7/yn
TT45zLatBbRgYKcSS6k2AtHIAWagb/tt/mfX5XZ5NnLRmUrePxOGzWy7tmP8twOcDZMxg3DXi4iw
vx28r6WvZgfjvDkIItTOGKnMYIQfwhzpwI0eYXdXLmmlYOdnIbBgYzZYyKq64DCDNsUZIcMwr7bP
jAxCQlIJ8aroOzoh1ru7ThlQi6nOIFYCfdSOCEjgW2pcqqJZt0HF+cP2DpAYHvH/K0oxnbTBIWVF
J2aABdH1eGyNqLrid6Ed1M3tItEdRDr35I4BCjFdlxOar+gf2f2JuxggfXgs8IE9MBLO47r1uLYV
rEf8sUYYnLETB8nyiAduwVT9Mz6wyHYQfcBacRo4BWUlSoum1VQ/O6n1+0jB09n9iCEf22oG7WYB
E4i9CUw0Vm1Q+HU0j9OVOX/h03XZGDCycNNCJaOzsRej4kPXHR3msaAlPEnRvUdp1/yErvJHlV20
s4XCTZPDGbngzvjHZnrndcL6wKnnHPzj4Le6QWHtaVvooVrdHcijGumw3b+pE9yUrac9Htt1RhF+
JjaHE1jn94rT/8sbdievKTV6iALBHerF2tMVt7f4rW9h+rHMgipHE2bcr/VRI02eTP8owCReyqBE
RKwEPYO+GVu0cBcOypJrTtgQaK4F4tf9M4HM8rfDf8dGcu7x+Ouz+7kaD9evjKrhHDqZt9DdK+KA
O9J2RgS68w/P3uHl4sEIuMyRPr1ACrYP0aPrz1WSjF7vG9/V1oIgnMZt83iaPOp3Ir7B+1DJ5R2I
RjjdtvvY33f3zRIm6VNivtm3xkgX60BJXSFikAj0QeBtl/i75NBxATZEn27CFMAUVzDr6VU7pRc4
ZC82CmlsZ6X/RYdfaL97ExAk2O7MiCGp492oct7pBgA3QcP03D5w4G9gt8TDX1zYEmrn6FX0S9fZ
s0LVnk7pZLI368Rclw9VnxrteC2OORtCjhcxq9I1k01noOWssMYrD04hCtjw2GzQKuV44RcnUpmh
LkBJsFy6BvtDfjUkSQlQ4i1LTovAAx+UYXzJk6tuIgYfsNh8N4Rtmzb8l9hljpya+HJOS4Oya6DR
t/1GITU4z9eGWXTeyDutwxq3t3rMKwARIfXvCMHQAB2F44Ce5QLWnNrVHZGU5vtJxdU/t38te3EP
Wp22p6MRuc+v4+JnffkJE8eeYZL0PpdA0vVFdcYtkAGpRhCmhfnmRKO/FN4x7cn9EOmacHmc/8eN
/yWDtOvXy3oAUzXeY4Lwuo4xWIKu0cwHYN4nI1vEPvs4sB+hi+Dm+1m5lO/gbaaxDcWbCwnRG5tu
12DearAVdC7uFH3I6066/54jtau8XGW5zVcAWT3xck5YHQWPamUrIwatd1dS/ueCkz0TmCv47Ybb
rkqGlv7FAfDOHlKunk+MJ6ZRFwC1cXdz1T8UOWUoYkp9YNBBvBy1xIDCEErGUj5hdP2LJ+7Wx8Md
JHL7UxtRVt4g4CA9zYXYTPEcC+fyO+gJQdpC/58gycqLLKIRvAk4af6PoNmhwS8W8jY3pu+Y9xXD
JGex4DBVUxAcCVqiIrsoN3B0dA2weT/NqP2HZUjFU2W9ummH93F36N+5X14S6uyU9OgwHN/Ksf7+
1EaD+6ChDVc3OKSuYKtPdN+iK3Fie5/O0a6i3xuVdbhO0VGQ/Nuc//fOEKKaCqudvVbvkWUSlPe2
sE/H5OjclMqk/cOHLfb2TOIUfyW3C2Mr54IsoXs7a9f8VlhA98LPVnCaBHzGt4uIJ0UFWfHzXDgq
Q9G9DSVwkeV0i50lnAsDRtuT/9r//N6QOfeky5mNwB6RVSecbOiDfV9o89rAGuu1xmH1ukMMBu7l
t71WP2DBEz+KvVR5psPoaL9tTFADz07mn9Zps6YqbzQuYgGyisP+gKv/9DFbU9A3Jk9a73bXYF10
98owJZcYYgkpURQ36ySM78jGYXyG0H5CmIjk6RKbcQy6tuUqMh/PT3i8mb4YRG1gVECNUmQcUGLs
qD4H7XV1e4cSKQcn7hpXKBiYZ7tJ91GkdqybXc+L/lozoIDY63rFfnitKRvM0IPukRpdF1MfAXT9
xx84VCefe8PhYKB0HlzdoGMef3u6FOVP0PfohGPs02TwOCigHWDTjOTNCZjfrejdguAkl+WAPAEd
rE++YOhsMLqHzQtET5oxqAPiqvmgGDy3wRhSyPghyC1oT6KB+9scP1MIeKHc5hLbJeCZ9BH/s57m
Cli/tXg/bPUR7S662/bNdLovvjtq1wO52PHwxvnnfWQd7NHR6GJPQXW6yTUf9pDBpRp9nFAeG1FD
m/Si5mPRGruqoQx2VGc7EpvYeDoA/Lc/9rJ3duoL4nn47r9kYyRvxd7NTvzkjkiCPCcvLpSkElNJ
Pc0PCq2SyuFBNPni5bCEkonZCAjKVyNhsCTTw0MjNhTycK05Y3qRSAbcLz3F/Wy8Qm14iAP2aPNQ
KaVD8/Q2SLVpe7PlkmrBtzgWrG+32MI1ymrN7qlpFmfssyqx0X46XZ8CJE0BoPiwVPonz50P6dns
WgmAyVmbn3UgoW/79Wd7K8C8ZG6KhXXI+amuRx3ngQrS8JGxJB9UYd/kuGadIf8H1uAecSHgjGyz
VPdeEav1PGK0UWotcCu1NIs673+VHz7ZJwzSJo+MJjJO//i+YnMeLZFh17kqLNAocNh+I7fE178j
enIBiQwVQyBBUz7i6MEmPhj4i7FRAFL/AHMTiif9uTVM06OWl1xEdCGVrclz0XevkL1aAHs54YMU
KCohwo5yET0Xju92yyJYawUnnc6cOfj857aLZ8miHakpudYyiMW2/jZhLx0SnlGmB9nC6f83umq2
cKaw00h84myL8gDdLOjT1qM55FeOUFonY3uCgq5uNI3SpX1oR06elvded3/n/hheEN3JoMdzdTqR
ku6z+PHHUTFvQfV4n1cFJXXnxPc973bemrTPwYFeeVGpDpt78euBEc1QqNKQPe20nr6tvwgGmJQe
BTMQ8N0KQ0iDEbfeH7S/R6kkLKJLA7VGWn/MeyCQZ1KB0orn0mKHbhYxDg4AsnfIzVhnlkQ4iYEi
qt9sIIyEa98qOKmW1V4RcndMv/YsdXuzr9aTP+DaBngtoHCiM4zay7ApqWNM1Dn9agcPknzBN8c5
VJ+ivLjRr45VlL1ax2OOcYMAMEjczAax2h6ygHLYU/9phu/Fz/jUxV7N/dCcMtykx4+c5fpWm0ty
suoxjnI/np+cjGQUExT4KS3yAJEHDe40HBiUlQAiE80/0fgwEUTPGC73dGfIKBDQXJfInlJLrggb
ArCmU9XrvqtN3zOjT0maqEq4qBUm7Q2iGJ9vhp43WdGjmKju7RBZduQxz3kgsdr8G3Vj+9odFNag
935BiJLoHyvQAv+hWy7UhEQyNheJcEFlNNtH27bPH4MddGsOYuG8NHUvhzNPxhgZiGhzPiOhrHHg
P3At8my2QBovzamI1XW8DGJT43w75PR2hYC5FXdrGreHvYMOj4h4rroeJoYKqFw7GRNWOdadysxn
pxGANxhHHqDacALH/W0ZsVUQUkQiem2s/zSNoavGHAsR8Cttds6SOOtjwcHw+hKvvNUDmbfiiLcA
59yCLZKMU2Ui+oAby59Rb6FkBb2zYC1zM5nnaVEKHH0sPvOJz+gVmc4msWvZYyK0wN3/HghsIxxV
TePKwtjYWvwzSvzm3yhiMru99mInzoHPSK1/EY9eOGwzboUzj9lE8yYAV51RB/UJYMRxE7OdRcFn
ILg4UBGho37n9rkeSjF1eulzLTWIKs+PTdeIm4jV1FymkDw+KWMeMCAgW2a2Tmm8aJfic8oD+XPz
86SDAS8iV1da/BE7NxrrcAUXbxpKai5xGqSdi8uR9MjOvU9b9Fe5ozgSeqHmimT8CbwEKrbZVKOt
M+mYl26UKnvYrl1n+M4pV7vtcHX0lmUNqXzfCrkiIKq/r2cz/C+0M2/prEhLst1dOiBSTIdV5CWW
e1LwxwzaIy8HrVSGZFo5WAt5rqDdfYkb/er39CE+LtmTcUB0jB7c1C9+tZ5oPVomaJbakxyoO2xM
CTjmgx3qKnIy/AXTBtNNJrqYLWY5HfhBZHTcRVN/cpn2fYVJ6Bhyf9U6qWEK88XOVjmjgV2+HXyY
vI53A17qU5ZyEmXIy30//lhqp2ruqy7WDwcf3/6/n0SzwwdGlGYeJw0bt0Dgr08GXrERWHg3VIeV
t6/yL7R/pqvnCSaXdtQ1NrEA6iyQIQBplCDyakpLhB9F4um7MWF27i1YqpeYFGVNtHT821xGvANZ
7THyuZKjd1ReRLyGyupF8+AxnHBMmC7fFkwkxgAnYknSzH/TTCh/pqhpsOcXhiOywnPJ/s2mGCTZ
SgVriSpY6LA89PmPO6Zj8YiQCkm1pWjzAQ7Bz7QZPcC5I8ScsXgdx2uWhEtkEUHSFkJCGpN4T63A
3p4S85KpUeEf84Yw+WpzRnc6hmNW4nMFt9rlNd0KV27JkU8CS4fyOcclURhEzyYdKPgcnqtnFV5b
I2mudjpinapq/fybcWzWYNpi4heL/c+7EygQrTeRFoY6NoYcc57TzEtvXFASTnjuXO4Ha1mIvXa0
/cHKBbrHNUpP6r2Xgqw+/pNlZaTr+oAGDxeQ1IfPRjMFiIWj+HxXAigGejvOQdq4MX9pw16zM8lG
nCyrwoyXIQ/7aaDBp/FadL4ZwO6SqEE/OXKx3TBiP5yZR9X547FiUqqm4pG3tUruBwGijgej3uFT
vOsCWi/UJWstTahbW+2vBdnrIJgGX5YLEe3ETN0lurMCocxBG0pA4V09i8zybWA1tT8GVq0aGPFT
IdL1aky7xMyDkjlARb5ULre9P048LwszO/uuWgg63hjoyUQFCGbqJXaPLahGRQj70WZ5ycrhEAuc
fNUPjtiH/4zzloEsO7ext7gNewbziyREUI2vCbSom8KzK8/XTWVZIYfI/sF/8ezdCo4H2rnALD0y
gFur7ZcCIwRzJCZEl9Vp93GDDqtfceplcx81JCgRggRZmulr+lBkdASyZ4gpMh4F83MfH1oIsO8W
/HHLAESAUrm7W17D6P4hr6ML0boRpNBGARX9Q8hFaoHn7Tsjg84u+vpGDZ7mGsSuLS/ITwgl7azT
z/dVZEO0rVKp8/gI8cNx8/tWOEaLPXGKTJK2/RyUrtlW/Fvays8GIkqWGABTGOTsqIvTiy1DPkbg
nT4dojt3HMVZmtG93Z5ZphWOEwkwxhhklSxlMOg7IJ7UzeU9LuYPY4oaX2bI9slD1LaSt36VKkHi
ZE1DRW4DkqH/hR4TG621xMxvPI2Ms6/xy6vhre34Tn7Xbc7xJBxGlp91Efnb0RI7uch2jRfI59s6
XaQVbbbebtsmj738MAXiYd++fKkDcCWotYCABfWDr8bIuT3SXAK1x/OwtGExoMywICHqgFgfwPGg
+oEh1k/Pd+X3bsKSZOB0HMKPdUgi7JqH8cMYAh2lZaS2HgMtjhqcAJO3Pnt8giUrgSgRx1GsRbXZ
u+nGiDQN7Bjdsa02TrKeVgpOfx0M5051PimmtZDWLD/PpEm5VpVzOYHPZcrz2IEUPIwSCVGHoLE0
iNkpltizGGow3MFXLzqcWAEetBSmPIlfYK4/P9OV6Y0CGfPDFGJoRxyu3Mhto9RVEPE9HmhHAqAk
xLf7bmq7tjHHDhfAGN4TLk7wKYi9H5fqN3iNkxmXoVhTIN0yb0W2bmMWSxHQ6snN4MjXKvYLfndh
tvVs+37BmSFZAvmkFxV+a6FAkSl9aMV8+qlk+ViqJywiUYMYSy6LFkcQWCpCeiGIgFS4rOruLvDD
dEOpe0xbBm5sUrS5vVa3IDli9GIuxFoHi8QyaKeSmykBOnQ5vavGTask25TaGDNnYWJfsop43FZB
tgaMXV0UQF4tDyIGe8+HKa5jQ6RNjLAUekGyDmgaeXg9SmWHrueHgKIBTShnajWpcpkHsaaSon51
26Z9JdD6ix2dYl5vhqAZP7CAnPf3zqkzRv48MTES3+bd9hu+mIloBysH5+Rm7CXLkA6uOAlSd+c6
dnRPjBsNlegfTn4kxsJqZbA8uikIPQFrUDsE7sbAK/YVSFbxL5xOrT3A8URHOS7F2BHrk3ZvildK
rMW/xTaMntXBpnZM2BYCKA8hj0fdctSu3+BXXHLMTOFNpbvhAZCkFXPj0GhDElAW9m8whYzsW48j
cAG9IxDdox95MQszPiZMILojzS4H7PPoFfttseAZXKYdbVjeidXptPlKe4qRGzyI/WuZJYGn2Zks
IE2SwTXWVaIHW2f0nGgG8ACvqTP0GJJSmNu+rMC71ihDOFNqso8/x+s/FtCirvcr50PQkrMrmWmq
u1FMokuvSGW6sUq7WLJ4fS8+4cKy5eu9x/3PWOhME9n1FKJuO258lzJtvBB9uksQOU6Usd0qRk23
TonOhZyhreypW0DCWVT8N1n/79pAJ9o0DDW/hk6uDXRnMFmI0sqYMaEsmL6U7yCXQ+xyy0TPMFzp
qHxLKb8KXVfkutaam+4+K5rn2UYElju59ENq5yKcjVVcsspwBo3NNGU8kmiRMf3oUGJqcXndNLtl
ddzVfVW2LH3/v2L5f1mV8f8BPzd9Cvd8XHh2dptUYM+wCir6kdIMzrSuOddw4b3WqRfwXD2+tG89
CbDUxeXWy4NbEYeoJmWGK8Si/SPz3yOf3QMoQk7Jc0l0XZeVXyCpekiFE+FQQfpoion99eo3Bwg2
GJrBQFwqqkhaEOpedsEfMU/x98edyOVowGaBiF3fpnrSnpvpY2RV10A6VnZrVAAK9u+D/HoInXmt
IHjtvRKMzlV7iTw62RDii3AxvqVnXO605ggSiL65SXi5D/mUpKopVF+BFBkKhpzEsS4y/SK/Ec2S
hngzPOZZ3ObuRgPYdJwdeLh8ywbAtTiEnuiDTwLk7VOELdrQR1gqqoaY6h56NQuvNzLeVh0Yzqf7
3wtNAyd9FQ0ENXHjP0AVhuISi97LiLMg4CBlTWH1HFAIkkjKWwaLP1om7MuytHD1Ltk8fS1RcPHd
edQJfqqlLbZ0uCPu+oLApnhnxzNxtfZ0l2Li2TJLyysfAvdoUreIRcIGCfuq3HuivRc0mRwoXF+s
E5o0RwQsD4FbeTOEwxsEY/F7hlQhN7/TWMmBUvDP3G65Nre9r6wCAwHYXpNLzoYIOkVjBpVq/SLD
QA9OedPpCm2IHWNUqb0Zpmu+F3RV/suIxkK9YQiWv/sN/xvfoqXdfF5KLxu61CQySN+oAJCzJy/2
7HYXZj3Qopox6Ny+8d/CSLIedW/q2BaD0DgKaOvngDjaBxEU+JV0C6mx7ommkwc05HDerhaNnai0
2t+K9B3Pm+2BxMrtvd6CfnV5VXdJRIOhqTDO0Hskvb7N+f52I0itbx4cNAxB87YkGMwJQXyTrm7Z
PHd3D0hteSBvOs7Y7HoXzOP2KTOlvZ4yyhoZo++eYTCsIdxkZVGX6pDYiSpr0QE8kskVGEKoceFf
0um4WG88vMiVYrIbLhUrUXICo2kztRA5tgVrl+iHFgVnjNYnHmNVARL+ye2VBMC2rWRxL95k36D0
JFhHUXjFkXCf6YpTWdNQhElRF7IapX3OnHKmgRYo9XhOEPOjzb8BjohXXjJy6VYkx7az7fJePfCk
4vHcb2Kqm23Iz3bco99lRRfm+UiPFF2fsan6sR19GGKPbNQ9WTsrZK18GxwTWH+xtMIEuKEjZghR
ylPmLC9OnL7netylffKqDZRCFbPS/YDQu0MLwHvP0hROBXNqWCO99EhXEDqIDKUILs1NoXKDDb41
4kOpNTbeE20NIUBQQgrhwNe+20t5K4kDH9Ynj/XE3ACSvLapVctuPp21JVpJQomHsM+T79klcIBd
vwibgrNbv/r90/gi7dwPOLP6ZxRTZvEhCnZt6AqI+WXRiZkPyM7715ONrfNOvup5y+QhJ1XClNGi
QmM3pTwFn6TH9aFVXkDb19gp7oO2/yfdvOt9dYJo6wnNhZvtOULFLLhdIZuysT31DOJI7jgvzVbG
vuMtMuULwSD3Pe0zflgFsZYyeqCFZQIGUM89aqz+zdBcBMIHrtfK6DnrTWPJ5fa5NBHDauAzzWl6
6/D9rYVWO9ykE0orQbd1HQBFJt3n1+O+eZCeuGrFealOh5EBpk6U5R4dOxQhTmFA2xWKP/Ng7QGW
SwMA87McPBUMSX8IpUkB6586ao7wgU1nlDhuwSEn16q7cKxmFHOgrMhBsBbKLIsEzWyz/2PrA5q5
aiffpxnaEF2/fiPTnyYKAnt6d7UxrAv6y0uIkGLe08YFbwGw3QDlBWn7KKoa8VtSSHFBxquXhB1i
e3v0xBntBj/HpyQtY/rxLdUPFpxKSeinuLDOJoqn/3G9FZcsUBNroRX6tLRGbNuN+083FJdwnnBs
+XpDO1NRR+iqiiwMxT4Lv6KPUwsJ2k3YkVPB3k3al3JnrItMNZGvtPTAftpGn0hDkxbhY/cViCcQ
QsdI4cRNkAOnWn4+RrHyYQXpe16jPRx6G/76VhaYHLUt8gTx6QDCIMSzErKgBctYnIXPcSRNjsie
Ax8m/D7T0hTQ1IL0alVro5hV5frQboZUzfYwZ7edXDZ1kLd0BxIo3yllNnP3A0fJdv/UmsOo5W+5
k9b63noyQ0uVjLO55JRppyKWzSwE5Zsx3LGqhoru/JZMXQMaRrocNemxggEVOyB9QroFfIrDT2e4
ctBfNySnVkvJuDaBSj+99hA1kDNxFUSc2/Woq6ewQfL4nWfKWWsDLwutK9hmhZfbgHoGrVSxOhjS
IBpf7Odr9PfLaMt3ZFXFqzbs+xUeABAMct9n2gwkh785WmJL4TndDw/iazjWjfapjcJyPnz24aNw
S8mCF8lOSlLXl73pyZ1E3T00GILndWRSkaKybYZNpO0Av0JjV4Ra1x+VaWQn4T7r+qZixZ5GYv+N
atUwa5ZUekyMAQkNSqx+nKb1oStRkWIE+fxl6l0megenBXLVvLsE3nQNIoJt2I0wVCimXZvT5hPl
5I2hIa+ScCu0qgNR+sEENBZ88gG53tMpC/o9QS1QJd6vSlczIvYgKMHij4zl/aurv+0eUhzTiAt6
G6wVnWlzNp8ocpeUP1aPeFKrWvyUkmqmgmzzD68Jyyt072jLGMc1ax9GDpJC6eK+BJ0awi2ONPui
665K8vm6YZSl33MHfRPHvsIM4tNKPe5LC9TeJtval43PjkENh8DMgVBz/if/GGa6rnJf6lSa8Hpe
g5LxnkNF1Wuj7U4qlZ2lLtj96davfv/i6s516O6C1uvj7C0LXmdYxHDsBtcSgMlRsCofMeYSQkrB
sjD0yMGOjF4ZpoWUadmKgPekrPPdShIf1S/TWnPvjwws8QivoOIeKiKz0OurBnlb2uXwDBl+g6OY
Lgwop54a6RndBn6OYpBFIDpkJ4nN1cFcwNe0X+RXuKhGMXy9UTT7Hctx6W5whZoZuv6FGtx0zH7n
WRr8ODR1XLzU8X1GF5RIoVX8XGLTwvlufxppLrGkqTJAyarzvNtyoHQ/IvQ7ZE24AIcOsSpj+fSs
HS4P3TydhRVR9a0aq9vKXOA5wnXmiPOduMuOtYzGX/kKd2DHA9QdZwRDS3GOXhpo2dUICnrReGn3
kV+MARkSoh3BG5SbsQEo5Dx3hmiwODbmcib1gGqoRbBJyESrR9WGFSTWoAVheXtWnjMA0sX1Yw18
38nvKa3K9MeyQ1hDlmawwvjjp8H8cYd7he1nhUY8AzNWoEOeonvDvs67DeEJny1ARHflU4TSqZ4w
2kciyt+eg2evTgAzJvb713XI3Tr5/2ejwql0JPgYGg3brilM5Jyo+Ucn/P2l1k6jN/VHd5ZVRuck
NixQ2gdq5OOK/U/xouGm2M/DvFczhQQ/tZzQS6HZTM7DuzITleI4yGeGYAxxyiBtjAcDm/HmRQv7
RtmBKlIiJ8vd3i41IdWml9nqf1MwC/jkDVfa3axzuBxopI0R7nMErd6ZT5/xJU6Fxasgs9U92Zhv
V8h8RtgFUEp3JzFOFUsLsnXaNQj3CNk/HedrfBVu655YB2fSSTppKd97i0YWfNKPFgij60HVW1r/
27ERl3F4jKbFKcgtZYKBJZ1/d71UZ2m9o0Laxkkn5QudJXNOMOqDsU4MW5O/EEauYQEXQb85TYyS
iYYtCoXmB1yN8ruuJIyvc8cySsR/ilTwiShprs3NZKAMPH/UhKgn0G0D08ItyES8wVhqI+w2ABks
rwYj4PfLf68Xf3s1RLeO60ZYZc6EmDU6AWEmAaymc2COMjESiVR1aVb1fMrT8cYP1BUItrFVsKu2
UxlUd+zqYAjQjqeFlJUFfFZzwgyLemtJ/Qg0NacFlSWp5mGT56h6HZwpOzsGvCg92HPPhLHGJKuB
iQ+lW/0MmKH92VZnN23qpzY5uDar17eKt9SN5cOj7o8FQ4l9XSp0894XnUMbcEskCJdSRmm1l2O+
7ViiEU2ckztzR1Ly6ob93wLvuj6cFXhBsySZtDbu8JUiN1NMfId1aX2x/5gm6g97/Q60SD2bXjNC
XBbNYn8CUd5oQiYAqDsxA9D8Fjk9bqFGTptPRrjA+pAXTcwAiboJYhcyK89YPoUQ04DXzXWSVL/Q
Lm3sS6dUf8jT92GQVK8pIHHNhbcCOboKrCu8FMqkygyGwy39NEvl3glYNlqixhPAaN1mRehvgMnS
Uw5vggnv2Db3hMaNd2+RVo3j1WBDfKC9Rx8VYCUnGgZPQn/Dbf22eilXvYUJ5Gjam8Zjppqw6YNL
XnwCFSmKxn6uFoHVGnN5/+EEAb48XUCqaBU6kESzRrsXzcgUgrzvk5dVFwCHTWiKFkBGBgh5VmLV
9+C364DhYMCWuVrQxhKRVq3aa4ZnWgbcGn4P3bvgz7uapHcbfyA6RvTmlnZeRGBcCcy7WebiUFmL
B8gKu3wMWi8fgOKHdUn1M60fBYF74z8CAsru8C1AxFX/yE/YJfNZJ39LSZ+6c9RakEDpOTf071RK
H48eSGWGA2OG0OkxACnSsAZfYBjqClB2MWCj12XIIvv+XIUFFPrntMo8v04Whzj4P2sQhAtKYBTH
xpHqwapbyKTIfrygIOXWMcXIklitYpE0qkhHZLYkacmld0C1mcbIgu9CkvsTiNU0YWO/rcj53Bdb
JCyMKCKZmA8omQL2DupsWLExLxnEFjQ1tgWS7FF5hxbGzYDyvjuP7ZULrz6AqQkKASGQDK/bI0Yu
AjV08COGz5+P598ERByEI2PLNXuppeAzQYaM/o3UQ7urq813u1+EdhEIbhQkD5rdUhuWPxvBu6R4
gpMO7TEOMP1On+LUscGzMEIQ1nnFzwi9nNqr3rzGY/4QicFFUMwpQfv0mULxgV0AdXRHBmJ4cteX
npUYHoNQwMbKmadK7qDQFPz/g/XoSIa7bC/CK8E6fs/WPzkyCN7GYIboxSH6iSHPJcnqW/Cg7n7J
M7Sg8/Y78o+ppuhRHK5JYGiJ2lC2Ny0ceYUmbh0o603mu7BnWW9DpHVF3HK1dr13OSwV5ya/3V1n
LvyJedbTW4eM7f5AYYw1GZ35RrS6hiOhXctJmNSBakjLBMnwbY+lr/hsDdVzHX8TOfzp/EcYR2Gh
Ejp9tr/3MfWxls+JJ6bdHOALquox1+PP2nA4+TBqCacirHotc39IyI+2HHrtVKBrTI8W28cSzii2
YrBjMFSjyYisuV7SxBm84NayQvmSgeeRSFWTj62PSUzoaP2/1HeqADtC0kP3Fn7sA9XHoWhYClm5
I8Zz6b5sJkZYTVmVHY1vN+lGTA6c41oTW1A924g+jvfuI5MnAB2M9Mer+TSqRsT5dgrAMRrsq4VR
NqZxgVVLecIcEbKU8ZIP/J1zXNkcDfuWSApCiwlG7K8A22zwt+X1QqYjCmyvvIM7M9+cibiVGUCp
AxRvYShJFsOJ9G9AkMyYdMbdCnO+MuFDHANv8JOus7uHswpwCB61J9Ne+pf2zd/fTg6CYVp7fd6l
MR5wrH5RXhVc9nQAwpwpVdwXnxJyrHQHIzUQiCWILcsuvM1dWgLSVmYDs1nS2y3hwBUnuH7V/ZaH
6eF+hTSYGmVoDMMQ4GVdymkxtJNW0N6Z8a/Pkdf71JVqfdfIowedO/xqjDYAiwJal22QBqcwPp5b
HVg1sBst+SgeVzCe6dQTdWMW3UhWlyU/5IVj344cD8iYarkVtA94cNB3LFLL0vbGRj1lFN+7aavL
QJ1b+fKMVVDeNHKq02cR3X1FbdMC5ZJQwBaD8dAZFU3hdMkkWUk4ogsD3w037Q8YbpMyaDJmytq8
69DZnaBeRZlKE6J8IT5hLFiKCdJLqnfEAV1sig8+0L22TIDro/SkBR/ECk5MtvqDxY/zw6GihW2z
pXLAPJhSh94aN8mtkp6dWCmaIp/KnVRC95UbjzSU7O2xCCNNVJ9EY4tKIBSqVjJy0m/RZBUs/uxw
VNnStVJ9d8GOz8Md01+fN+jVmJS0eOXEaen9fVSSu7TczJTSq43Z3QajY1rklqV5x9Q5nIsXf0j0
As5RmQHIaIrHmd6MEbh3IiprdG/mkNwU8YkJaEGueDqT/MwO4z5TyT4h0BGBnUVx5hVDjyt/9+Ju
YBRXu9cdD7+LkvDhtnrtlvX2XEgNyYcr9wos3BY+w84v1oXTwMO8b4g97a8D2eRQkQXBGLT8+2eS
A1324nfxCG3IMwuIvTCWtivUtieqPszXK73CTnm5a2HDXBV6yt67gkJp3x0wUYmeqYAgPRZ83WZv
vAnzwz2YO4zsb+xG2L5OPQQgsaI284QFpkGTXUL4m6qT1IE6ktUaAlUlFm2JIh8bTs5+P/tGENW8
0118dgF7R//FfmIqBuQ6CX+2oliwpx4thVUZ86eZk0NVsrVkqh8JP8mbq5NOXEhqonN1UWAbML6n
U5uwfeb3ZEU7qRjM13y1DU1beLqsPL/1i4CP2fJrjzLHCDtkAUb/9nP9xsMMUZ4B6P/9lEJJeWzY
wrQXA/jljFlFDCiHAgvHFNbYwDplJguIQrvGHbt0J15UrlyWXlOo7L3xqxSr+axFSb27n0X3QFeN
Oc44+CGAzUFONIspQoDuCfPQVqOJlbpctmibaKkF8D9N6K7pnGs5sZr39z2NVAphB9T12HX1i9my
6ycGtRAJA02dAktcNZsUKIUY6wKFgPTP0/ZbFgFzKKK55zuA1jp1KB4eSCjhq7fVoGm3f7ar+5+g
G806Fk5JJoBA+TdKmkl2M8uitiHyA7kb06/vLZKftEDM7/x6jb8s33WFHnhbtcLJ37gLONUgYkiP
Tsv6cvvFG2eowvWQYwAjjMl0C1RdSMgca+JG5klcTYmqv4+3Z/wDMvrd2BoXXhiQTX4HENNdkVKY
0dvO+jplLQS9VxZl638Jzy5YXZLHML++QidnYW/dLjmkELRdBS7P+dUsACpa16X/xWQJ9oBusICV
QWucwDCnmCzDvEH5vKriw8iLWslqBF2Ue6DhFvTJ9mucFPP3aFQjohhe8XLOGXRcwgXuElpjbz6K
8B5ziGQa+nW8UmQmk4Z7tyRpVkcXNatVZk2DLvniWfte0fEgv0CscGPdxjzlmfScZt9y490P/Fid
BALebo6oFW8iooLdK6fqj9Btd2osavlp7MH/SidVmsKyJOsifOrDFnRtU198AmN9uiMnZH4ouJ8f
s3NRdSMBVopqF/vY3bbCGoHIGEYgOqWYjV6LOKRFfXNanH0fI7N1D2T6gepuUC4RgoWehABlH5Q6
wCuaOhUbiTADNZk4dMuclgAzsOhzXEcq/lE4caQ4MLsMHNZPhzLwFVQkR9efU54fekGQsQrLWqTs
SvS6PmAPA9uvo3FRuEtdfuTHAgmt9vsSfgIlmOxk4Mz1iNPux/F+xbWOAn6L2jdZ68FfDTz7/6qa
DpUdQz+zBNR0kPn+4lRoXX5+ZwZnJ8XoBOZnDEgbNNilSt3/MbHfAQmcWdQUGHed0REaQDzKmm2l
wwsn8OlHNAN2lj0YanL+PHrE4KmqcmiO+tNx9C6WysK54sfg7K0i1BgjkrUmvpolZjD0bVKWfMQH
q4eNLUSQUaIlySlaDmc0i/6LJvBjGJJDgwsH2eFcG5V3p6FFBkGXj2tTM511eO7Aya6T39FrqI8l
OHJCody9tiWppGgwCckF0kvmyPnFEi1cKT/x45WGSGlT22poiW5H4OEudGkebaEtEot4IIE9/Svg
pQs9G2bc52lrvZMO3jWfL+P8fvziMxx/UhWTivsFjgBfYpTaZ6YmopWKxgKZed0yrP4BPFHx50ki
HsY1u/DVpcvNmMulBm7qs/xwpJoxLoF9rcwyFU5FHvm4gP7TnEjZ/JwKYi2zMB7kr3PMPb9Rz91E
PH3IEBqsXPiWIg4vioQK6G91rFxMzZbRxIrtAH3hE7PGLf4b/8wOvRsV31WesE+ryS86/pFpscy6
We3McRQI5yBIQxLR1tcMKBNS4YAhgf8bs8tO6QA88kmThA6T76DzKJ0sNQniXtGKwM7VHA2xcLWY
JrM856hsM6zSpaE2zk7VP8TSyJYqhgoBgefobc/1NuVMwk7uYkl3bxkMsnUp6UyOHQQzVscne4gB
ILmiiGonvbLccu2W/eOZ6aA4/+WsC1iUC4y0b2bMtu/IQ8GQzivch+9lmoEuu3cH5HOEpF4Jy0W1
QcvETmKnIUcdapz0XwEwoOHzc4kLM2MdsbpKqO9B6q3k6sKguJCfXIvpQAP8C/BoXvQEPpWpH5k8
gxNxmljr7WJjTD88DafMIE7dZjEmE/Hcmy8YU5WwtRXEmZTJnDceDRZPwg8fZKjzBTExkU8TO+JI
X7wAHnj+TVwXki6e6brY0RWqBR4fGyWJIXbf8qDKRYMVrzGqi2/S8y10ngIVvmm6ISRuO3FicnWE
tc7CzfbgrPIJUTnOevv8y8oDEF7BwNokjbi9MDEDrGGKQ4la//zroFkna77mP13u1xEVk+5rsQLM
cUkE6K00bHUGuNrjFmGBEKif75fzWq1tr8pEEIexPOTYrRpGGM5ZwdC4Z29RhE+n8ARM6WUvUxBa
ZKf+5iX4A19Z4TPAYRP9Y7ItD/OK3SQoQzU1zWStFJ0e8gtPrc1q4SNgSc1Sbw+jSbBkyXtgzPtM
FGeQ1HZwnX5q2dBwqs8qKxGbTtokE9pz1VPmCLWEXk0JOwnNO4gfEWFZDA6HsJaKLpIM9JQviktu
LnmV1Qglj+idgsDRXVGCER9w1ddVJKKggJrgTkveY5EtU6yTnXSVYDGzWLTOXC7/OMSdWy3Qt6YB
gEFBOvJt46YOKPkF8caj1UZ1873yMnzyjBjSzN6/IA8vzcxE8mTZ9eY1OmUFd2cR+EQZ0v/qxeL8
o5gwRnsy1oKd+y8ZPgKxxQ9EsAot16cS/WOBFIBqc1ins7edQ8QDdbmvSCnVCiqfaV4qquPeRnZg
ZFDzuefiv2TPLhMcA/mz1dBQu3yedXoF3Yoy3SzAEN78WXbxZCrNRsJOZpwIcs14CzmOSgYVTxQ6
3a42/uM6wOe+1gqYtYqbNP2lDVsK8K2AEanCx6X850y5dLCJOeRJ/cj7WIjiVzImqCx11xiW6j7j
Hj5DpD07bD1/U4vnDAg0wDY3XxwfSqSvsJ3zj3lF9jkKsealX8undsOO+bdG021tTdThV8Q4jCgr
CTsGV9TP7rexyXhNuJQrunA8kVtjFvwaCLdR5N1lNKomiXYBsbo0GFIya4ao1o+yEdtjKOcxsQ3N
0njjdtpJu0SB5uqUwtYvvHyVvdqkmtGQg7zom0W+oAwO0ZZgYRxps/xAhZZL5eRIPEMAnMFM112b
EfXbiwrY5qMnc694bFwPGHlMXzuxJ29y4gGO4So+p9rvr0kXgk4Y9b47gBiw6KPbNaa11/Bs/T3P
9v7C0Qph6f8eEYUPD9adhD5WpFphu/r5q8pCujSclRIwgi8NNkzv08Ki+bxl88OamuFaOPR8S8vq
ryzFVgsI89DG69CNg8mSMUDjDfRtP0KxaRKTfCOuPKMB5gWvC2JEzXryf8Vv7MXF4jw7ZiluKGhK
grFBvKwkUUU5ziPMuu2QshDYWA+Acz2erk12BfCzBZiUqWXTevzSb8dFBhjOiOqJeSxv2yB6jPhr
HgvaHE+24tCga4FuxoJmJEPMmuZTVzBqVnoU1TSp1VDWAIQhQVt6IHRBAkVXNDJkOPtqBKkTm1rE
Y8P5j2RSBWGz73/B269aCZ45Xbt21BcWADC3jl0KVREgX+BSv1YxgI0+1tZcifXe/JvauoK8+9p1
pjVfz29Qo3LIJzuy0nCLQkk7QD7WmjL/VbgwSpagUfrUTX4bO0JlOAebPbFYIw9aNmOBGITwnO4K
OknO2B1J+gnGhn4E3aOzsANQF29KyPX9wYRFNuXgrfjGGah0uug9GAPladKes4ZpLIjoRrWnkzbf
tF58nTwZwOw4QPsPKGXXPYMYU3I4HwYFU7UFIy4kUAytllyDj8HsK/kvO1d/v70eX/zuiSMPwcmd
mRF8vZ9bOq+SFhsZ0HthYP2F7kXhTG2NcsVRqmOuv2SWUuXBFKoEPFmm+JIffv+qI/9OFf5q3wD/
zTlosiW/Vl6xKGt1icNIYN5R6gTDGGAD3nwtPmVEKlBdz63A+iLYWAVl5vszFJTWWuusuvcVDNiq
/FEpLxjjlhUfdM8BQ3T1xFjsaHqxKAQaB7jl1E6L9Si59q1N646WFGKclcsn7/sNK/8tGO0JdE/E
6pzyJEfrE8Cd5+C/MB9giereXQI1Jr86rWj/0BN3X1B9ejN/o55kXoNJBnRqi0zWQ8wl3sfOUV6V
RGh3xAPTZEXXSuCm+luuAnnNHR+PjU8p1s54Ao3aJALQTXyEeQ34b3IXIZzg/WyeTJt85Fx2vgEH
r2m05qSH5de5BgUg8YyDxsC0vId2P2JJynfBXw4qO85NCIAyMBgQSjCyjsIk3Qf/AuxgOq2iB6s6
3yqa5vZeJm3VOk2Z1EtKKmoOEO/IPEmd47iG2TahTjhSeISIaNOcPXIOCdTbwT7eb3HXiXZJaSjK
bilecsLwJVA0fsgHOMNqRL7v1cnvC5gyXZe/ZiiO4yOjl7vdUcT9Em73qHVT0mNrsCsA+sFrYtyO
HhnmFv2ZoE4cvKVOGgviZs4HBdcDMuKkfMbavPaXvC13gToi/9wxW0tiT3iya+CuHEcJbzYKma30
d0UODS086ofHzrE4gEyAvOzVy7xiFKaGxIH+8hG1IutA1umD6Cc1f1PxFK2qXOOgjPkmRjfvVS+v
WjIBhNoil8MhCwaIkRxXQA2mepCHWF8SXT/i5rQQatyjAJirC/FnUukx6SxwTeNPVHOlU8WcpIEn
HYmpS3CbO+NgJya9WYKBtOmnwnrMzs8h/EOIO7Sg3ktD/8ELBAyeNKlkERp3vd50nu9DAPizz7bJ
FaK6HA0bIWMQXQLmfbwslUxRxw/cZUdhoKbM3oi2EhelIrsBsJflop/MmRSVS2Z5XvzjfproHOXH
l9v3yTX5nR/MBWTca46k095YjQZqAAdZPeLGCa1RkchWX2c1hsNwEm2WL6u33OaeVU5d5shkCRnp
LqpGYs49XnKJzKPjulmN4dYh/oXG59bSGhdPLe/Dst+4ydzgEzVB6DbffPWdzJCStbRWi1zeV/cw
jHn16VNJ9Nt2UjP6RIL0Za9/sO3SizFztbGBuWIUX24MtAxiUM0tHfJ4sMZGOBfWVdOLU86eyLxS
hWrac3/WNqxuTBVbnB+LZjM3ZcBf5YLSnvErQ7vXiiGnkyAEfN995nvU4ISsr5ING4OTdLLkn7zu
ypNMpDjzLEjbhXnKbUHz89IAqnbgt1+GmaVYIqNSuoX9zgxc/ZxmjOz31uipcYUgN7XJ5PnehCL9
1zqlM++rPH8S6sApfxaL4PlRxjOAGP2S8Zd3CvrN7Dwk9pJ7GaA8gVECfk3azeL7Pv0fhSKwdQuE
oaF3pSFVcHykCtP6ctBHeEqXB+RsXDsjRMit2jUHye94TqLQa5YbCAZVanQkDO7wr5O60aGncFX9
NNo/U0L3dl03oMSsVX59oMtAmjBw7in6s8CqnL3LsqFMwmiwzyNblNrMYAtdFv2A5IYHB62Z0QMN
IvUIPYHVU70PucoKhcn7ry9OjYDz0v3HzVdr4vJUmIzm3envFOc1l2c/16PP5cZK2Ekm8pRo00DT
Lz2OJ4g6/MonMxwhh54sHAbtpOexgOqe/S1+Mne4SjfDlQr6ZR3dsmXIqyd1jz6P/ZLk+Bs0Pej9
mntzAoUEeoy44q7KROnXEXDjbiC3mE/cH03NhTpCZu9ac7qaAr0bUpy1q9Ne9UVV96UbEEbFjWe0
JP1nAf5y6V88DM3FiUJN4uU3g4vBVQr2C6CVlpy6XIUxAFHIVhe7y4fUk2QMdAFUNmisMoVJgBpF
t+jCvSweCGct5vXmAZU7YZAUObYMx6gUm4qfA0e8ExUEzOVlIhZ/L2G0mFyVVPcH6YDZE547XKgD
vv3xeDRs3rNnE/3zplq8oClLglL4A53dKGpSChnHYg5UUDm+zpOfBsS7DGQqA7y9z6gMZGBSSugx
H4/9BZdAVxphpqKqYNox4CiriuHmYNX3/jGtxlQthv/oVTjoJWwKZ4A+R6A4mtZ7+ICWAd9WtZot
elOemyWYnQpPuP5jRY5hLLitSi59qkaf/eXs3yv7Th61dxuCTXATvfI4pmQAbP3IFFm/FJQT4pGs
UD4QtBAT9QgD60GAvm9y6bqiQyHtjdHANrCAwAc+3mgqSnvL4ZzgP80CO6V+eBXRuw1s3ISEMXMe
Yi6O+ieBpyMwbRlXUO8G4N+L1L3pJk9Tf/JgTUUR6+HjFXhYjIfU5ytnJ/lQQphOOwSiitT2M1Qr
joNHtahveKqGbY02l4cjaClQ4n5fOT8t0wZteBXaHnA8yxUddaT46hpjJ4CtlW33QlaRb7W0e0Q4
OQbFu8NnTFgb0w3XCXxi3BxFaxzlyCQD+MAXdokJ4T3aZaxJi8EUL3robSuqX2hLjv+tWxnVzmWN
L3dxnRbSStfKjhF82/70X2c3U2+W1rHfbK/09P+0idGPeSUCbUgyDqVeHoLrc0VaJ0TvgVn+SxOh
qW5Sx/HzkDKSAXq7EAgmxnc9pEIgkKscYoCdWpn3rWpTUbunfi0qF1Cy7Wfk4MZNXfSWcaY4KBrh
zBse4o/ps3Ib6uAGzxRqChkTFjqjGlmehIBiwdjb4rhx0qTh0B84r++PKIXZBW7pjvUkGVMiVekj
ZI4MYgyf/hUAhFeY35M42yCNeUTsAJxwrprs0I4gKj7qwI0lgeT9pyJJ8GtAfNRgE9wklFaE8VYd
wUZymu+Upva49WOx3mR9ecg281R2HxS8fusjaxjTZdHFuJzfbAnnsznCS8AgsNvKGD8HSvrmgDBW
TykWDQly1mAGaHt4E3EcSsyxWcXx15Clk6Rvuo3DZo0eu1b+EhUaZzddVrKREueNitgrg3x3i+78
TxlOc+DFvI495cvvJ6LYFqyjp1cAME2sdlRFLr+DGGGUqKB0HLKMxphGNRsfOGoktROMm49DlYa2
lV43AhU0ItIL/DvTlx9H7RcTlBPeVtqg1HwliNRDbHSCavEK9UvoW5WwPZ8x1RysID9BjLsqfNpn
x+EQNztxO8MIPA9jgjl2EvE08YuApd+tB4ox8SCGb/LbVbG9TcKT/MnQXgsHTH7rROPS8tJfDrNV
1n4rJv+FOt57/kZp1wpo6+8eizKsww6nVwcX8FoYQvzGvzs8mwT8lR3uzL/UDQisqhQ0koj6Zl2m
cRHQjyOcqzEEYRm/56VfdjhusP8ROr5EEYk452jHMgJGt0d5L0/7xFHdoG/YjSRpayyA63TfAAPe
GAQqLUfQpSO9Nr/Axhrqe29dLzMBTdYzR8ecLfuYsU7I0HCD+542Ddpyu++fHxh7/1BKznp/0LEr
M1lHo75q1IIPZpD4Of/x1M/WHw00vMJurBrpT7WTLsRrf57XJjT9w8xVtG84sJlM1+Q7aFMqokra
3jjNngfYJqsUCC6ooy58ocqkpsUop0cKSv7RAZ3JQ2U59VBsjv9Dc3brLIXI1OJD72KiLcneituX
m76inUDWrjA5C2Fnb+Xd3oVTOo75rHZhcrvtdT3UC+eSBAQc8zPBm+e9BcbEYTr6R/T1nF5j40uR
OMWb3ZwDRkcvOcM0h2+IHxmFeDRXx0MwsQbgtPB1pyXCzpjKJigjC8sXiWM9Bgo5VKWWAz71v313
y0V8/P+fsopMUcuEU0CLQhEuJv7hdTjFl8/YQ1LjZwHR22g6XX00NQIpE3poFCywqIuEH/FN1tny
TJIYulYpJQGxum6wl++onVwh6uxwx8h1j/Wcvzht72oQ5z/rgbxaPBUc5kMN5DKdI/kpSIdMShpz
SSXsfVKK3kpFAyEmV5NLWvTAehwnvE/f9c9PLMgNA0p0xrU4o7+1mmSwdoneqKd9IczlWoEZls0l
+MNb7ZqzDiOHrZzNdWZUnTBXZv4zgZbusPbE14aAe5lGcRI/4tUAVNjFFPlMAmoFVfGcZj7YCG+p
rdu7aywaPoRqgGr1Wc2VrZH99It5RfiByms+udT8ZnfZbFcavThM7ZGFMA/h8MtuXAkdEqj4OseG
3+IAANYRlmmFFZnRUhhhlrAtnTPn2DBiq5D1DdOz3YTgI9L5RqASZmDJr/42qxe4fn6vkbjdx0N6
ooJEiZPsWqKnCGKXBwawJWB1p9PdhSpTuTQzsmzYdYccZZDViLYV5cL9gjcg5EzFa+e3D49jwk9d
BHyquhS6zjj7LPdek02TXNbHtOV4AgKx8UdKf8HUHQBeHYYHtwfg6xe5yWSAmQZG6hwO9A8b2vec
qiYhfNpx318NnXEaFzj15d7WADAow4HWCEPk1t3t7DxeLF6M1Zfkdl7ZBStyZjySTNFANVUHGYFi
SYC0JO83HlMR4YdpeMce/oG5UiUyC1Ihs3+DfrNq2DW8Hc4Mc07Q7XgHoMEfXtQ4qVwyETlCbVx7
+PvNCijYYfCADgp0C+qU/pr342Dibbt8erL7o3D0lZaPicGc3Qell0LZM/xd6MYUebRkKwHFRsGZ
PICBKYZAue+4k7gzGm8RZ7kEnhr6KL82wzHN7cQ6e7tke1wi/5crrEfUc8hrv6/FY7kW1+YinVE2
PB+VJpzKGeW7xGxfRg8RCCti0hSZVftAG2PcQFp1ZiT5tWkeqK7KVlxR/bGeUXtb+ig9tIsRS0QF
DKWBMby+E6e6PpuBKcxgv1/srnAuUHDrbmk+HihUp4behLrkxXAljHzOpsl0dMy2gewD9xdwjeqR
7noeDlTT1yDKhJ7lTPZYA6wgksGGOhxn8nJz4F7rqRsj4WVnRxhaIk0h1na5cEKAqij6KZgkJiuB
kURG/9Zn9zbVGabNwR2qRLRt6ECMhkzruEfZ0r5UMcm9o1ROpp2omGrpf3DcSAjAGnxAiLuP+QTf
uhuhsZaAxObywiD+zSH+SBDESSxQOjonJ4lUkZtbVivITjRJoT5EXswMtC6Nfid8nYgbdaoAWIOu
EmKdnTvx1osQQUi3OKxILGMzA8ruKUAzDDC44WDh0IYEGA7H414iyy+RLgROwHW7I6d2A7mk0YUC
GE15TJ+VPMrwdPTsCdBORqN2pJ0wcOMXM3iZFhGBdvZBDK6YE5FKeCalBFUfU514tZR0zXVoXkmT
BeGQGVlrjYHR6DbSHl0gO5wqoa4vGoxxUbSafdVGnuhcpEFsW38ywCzPqRriJjEJXUWon84QavO4
YIZgymgz9Q0M6CXIy4SUNBZxrTLNgxpGZ9QrHn/Brp5gm9oe5HHtqDdhEA+qBFa4TK25iYxLrISx
b4ePlbaENuVYvC+UnMaVNiRHkHH4XxoO1DwySSDJkNGNzYSDMCRjD+F5zP+gezrk9RjYjPEjyXNP
I9Q7lxWtPPIdkm7tSCy9aNCxK5QxTGWnQs0nAZ1Qv6MgzWGMt5vRMBw51/I/d+HmKZPCo3kALmNW
zEFd0jbwBwlTpTYweGOuIFCYFOUhmcJgpo/nU+pRzMSTP2dcC9v/EYSnMFILG5XZ5BdWHdAhcuuv
izbP/50KP1j2UYjrzGaqyKyQ/hzuPiYQlGB0B8LIr2lqMAC6YM1e4rXfV2IQpHoLXSYoK67jGzu7
oa6qZvNYw5G07zrjQqn1hOLLnz73hT5oaRz325+7ETZuOl1ss6B6TXwKzBJl7aFOPa8cXLUms9JB
Cn81iiRkTpQOg/wnQ/jwD3S6EhwNwfNl8ZEtrA17A3023p6J2ICsC6e0YKFtN8xbw5Wcz1FlRtIA
NBHPobQYi8NziLq3tncm05TxJ3b/caUZDYqodqeQs3ETGrupvoymKWe+Djft93p1CFvdIv+NLOii
bpfOJR4o373j5duvDuZBEPclzFhJmLODsrcWZKRw85wABm2AorvN/6wJlAhz2jjReAsQfHzVeXlT
CEJw3wzCmF5PVoXhErRgFdtDtyFKFkMdVwDo2JiYoyMNZEVYv1/9O6g0gqVydtgnqCmOZf/O8fko
XRsjob/cxwt/ewOncYVvUgE36SDBS97zXjcP554FBIpRyMXPbnX48xjJ4c1DRZzOFv7ie2pqvjkb
s0t7mzT7ZVLt7CNWoY7TqfAlkWDM9groNlx32NNczLzGMhmqHliGSh2bcZNEbj6+B7AHvMlonkOn
QKLtEcqLKm78Ia+IFT7uUbfgWZfq/391nDC5xlB5kfPnvoRtdeOFqaqHJCsHliBHKSZ0WynN7RVR
yOTZoVi/hhO2RKe+IYb8R5ha03y5TmD5zwF4BK+8OiUhSy+Be8QcnVq9c0j5wcQjmsWFy14dX18V
gsTbO3shr4esTHAxJDx+lmnfaqHhkkceAFfHrhRnfEQG827Ccejqz8MJd/JzHOZUyel43H7+8abd
IAGwV9Y56hTMmoSsKmL6bjaUPLM9HIdoo0ohsllSRljMwl8cF6QwWr5hOz+734BGiGl3Bf4aYdE5
vZB6jNqWh3IUG2ZxGpvvPRpWV460fbGOZdhR615/W5iQz7EftMYR+R3I6E2a8edBPTnr2292EEA6
LNXhhM3ltK/ryd+C1q2/X+tdWdeFGTqIqmWtyOz7msG6i7YLdtXihSjc9TuPJ0jSaAKa8wAiEP8V
YuYjmYGTPNYfd1emhwkmEkGeX+FsnRpw7WYAi/v3rXvHtbjpd7tYQEadP4dU6iANuz2Ts5E/0xBe
tS2xh8S2TyhMGgDrZv06/V3tqTv1wUrY7RZZzq7aJ/uWmLvgBzAIluwDGy8xWG/3rDZSvye2EQ4+
C/BjOJnPo98PrlJ7hdrJOxgHsIbXZ7yCTOy4vgipZ7zuxuiu7zr05KDTsAqlX9oyBeBD9d4ZcPoR
Zh7iXTidNphJYX7s8k7/ND23sANKrkly/+hoGPQrCgJj7NZK0HI/n3lbyFFa2XCD3IYfYiIvWeqR
GK+iW5TRvpqt8pEIL6a+hd1zxK4SCKXqZ1Q+yeL4zxgmE+Mxkk6tLcVAold6ak5VcLvrbIPhpkDb
wK32r9ArbgLuPPPnNERP0xSughIH9Kz8i7nZNDt+loGVISsGasFvIgU0evkE/e2uG63AoB4QrIPC
qTZlXjq36/ef8siw0WGxob6wa9te101ZufROw4hBgLwORg6awnfjfDsY8P83iA/Vx+5UYymrsXAy
Sos0I5McfgDA0SBnTGCzrJ2lF13D3L7shoX4z3AsL0Fa7Mq7XtraPNs0E0THU7v+OiStCK+KcVNi
eJrRI3uFWFmM2k+PEIgEGzIaUPR6VK5G7wkZNAaNXJ5r4tJIgrd5li8vVJm9V3NxWFjddPJ3ymb7
Yid//jAUnYWFqRGua+os3paRBZxCE0FRI95R4QbGWhJAoSW9WJEBdGyUWfI6W/mcRBAzSNFk6nsP
QAw/2mTwDy5UPC3n1/rcgEuit1cISK9yopGjZtcxC1gV20LEhddugmw+izpG9JS2a1QIZN67HEtH
VL+iC5v0ByEIrgiTq2BdFbHOXu5gT8PkyjspvdQHHGqgroaro+MA4l10okFI5nGyHHIkZjxZ/tWX
y97L98GakjAF5nexvgmomXOx2NpcWF9e3tGbez9PJYkCBocQ9RsJ+iYXcVHR3qO+r7Br10PTqayg
c1v1KTBBZTS5lmW3an4ekEcI5TNs+XlsTlUBgPQ83GH4y8GU2n1z8cSqUGmUNFVnqfSeeeuAsa/Q
EkqMqzNpV2oRslLYoYNpmOaw8tzDtb29t2XXuWYMl+SN5HUFljpbQFfJ8C+sDthyhy2TwD9JIWhk
EzpJmtc8QTAIAC1YgejNvzpRogWrTkhQ7wQlAIYkO8VIVxDilBE3OJV6HL1RUmzLrDIDI5X16zRN
j37mKQ5W0T4XVAGake0NgswzLYhkXDZalizvLj30RxA0W8d3JtgX9DdpcuCNNtqlI/U/pN1TBdNz
Tnlo7NBXLxRbv03DU8/EyD85RPDLl+cfkXCieGMp62EgXf5OXHMiPmXf98/HT80BXfGsVWjUsgfM
4mzGRB/d+QBf25jSSH5d9c4N7uWjsyjwEQSjUNfIFFzKXj7+K449tTg0O8mc+GQ43ejPCIGr2X/u
lcYXzRpQigUx5ipwhSAf4VS7k8SWEwyfL+WgiSJWIEisTZnZkLOBIX4bYMklJaDlXTpjmEkEICg/
y4LE4HxPVW1WlYIU9XHpQpUy2COQmQSC4QqbEsHOULCMKGnKKQUnYuUqK435A2Uq/ZBi8ZotddG+
8rPYTsh4DIABfIx8R6VyVpXwJc5qzdzThAiz2PBGx31QHx5tdKK4ymkcyuY7fe9uBOq2W+nODngX
B8gbgGAT7u7ZmUxICt9XRj5Xr9ERc+FmrlNjLvsZDveSZKN3Moch3/ob+mwNMlAXaHeAwTRpQgDB
mV0I5hGsc1/PVdRwFRb2/mpuze1/N1Uj1E2KuLn8uHlfRIsq8L2YOMyBqaibv/Vgc94OIBYJNKqp
GOXWY5+z9lrveKPO/ps0DvoYS6u9UATROh+AJSiv75KMFezHGBI84it2NJaDazlPOATNJpjD5qw2
XSt5fasppLtiCtkf65t2wcVkFuuASGvtDUxZwK99ay4kD82WN2fzohd/Z3LuT4JI1oPuu4QukpqE
6gx2ycMNtlU/KVnJz0jBqvD98Bqu1GQCVRNpfoQmkju5RYIvuabx0oVeApg+QkkSdIdbQReS2LkM
Ud+9LF53Wft0NCy2U5fTiTqaKV22TUsGFkvwroRb+X5HQBPXbc8fn/YwncSidh6pLr49Ypxe0ifa
ulIQlefGSBgmq72vLCvLw3XcmrH4pPHovWnOXb3Vhio1F7qlSbMfTPTICq4r4deEBez8n6WOQRB8
BLzPcZuInmdtyce7byJKesbzv6PUNom8JrdaPx3VPbf9vr7DNnxXVLXl10WY5x7g8DrYtvhf3vFj
itju2Xhl2U+uolNJrlDUJQNRAPvw55mNCbSxqLzypNGvdW6BCHzYzjyMhl4Z56P9Nxe6J6dnO4YK
XQ8GzpJZhg3Ud1E5rrVcHkMtuOy/0M/gm1bItGLvR6/N9TNgOjwHMaB1Ln8+l+74Nhd6zn5Pz0Y9
W/84On9n+RPx2cdqrNdMtm/xf1huXWf+Vti/SWb1QDxjACAi2n0S3LcqbVBia9FqK4VyqIHgO88r
4F8sIAnJkUBwLftnmhZDSYdxNeEAd8hr46FYSIZZGz/yUt2z2ciQOl99Q6s3Z3xpUTat4zs0d/Rh
WBaNhaer2CYaxZEDUUnSfaShQuJnf8uyz0GjWNNm/f3i+hu0xNtS4Mk5+u0D84/fqGBHpPO0F7UF
iL1I20w+VwoZudbMbO7xja+PQ6TIoUtjyOJxWKMcxStWQfvfY+R8/C38rqvkaUyd7nYfDErfMAY0
+mZ0umLXULvz4efoVOkJfVpvXPJM8vTv4jG00LWZkKr7TrfGlQarNFoI3QmxHNBQgcX5G58vrptf
Tssmt0vhZcUfElYbPiA5WLzEk5drseJ7qQl65jpsWxwAjl/EXxUP9yRHgpI04srQbU5ZfLfYS5cL
qT4ON/La+5UT8Mcz94hWj0xludmv1LIsonghj1ytLpGbHjF/ZAV+BDr7RNzna0QoLhF8rdyJT1NT
Trug0ufnoa7QOsUeDV7FMN7r/ngLCEuFkTQ/HrP9PoNBEkspGZowzYtKXQi1xfjv8GQCYDkyu4Eu
rZ3AjRIbUYEUr8qDyVsO6oteFPYEgfKVXpF1KSKpvcaAGvlhn9ZKccYsLBeH6ynGGsv0LDROVjS+
/KyHxGUVU91zI9N4XMJOTIFTmkouhpVh66hn8k1ZzONjFZ5l63a89Y1OOk8THzpbE2dZbluSyfSD
7aJeXIf8ED+Ddt8QNmc+wBNSB/LoX4lJ0LpcVtOSiEvP6H/PnitSWn0PCQ4JLtxcgDiP8nQN+hSB
v1Nk7hdowodTkVwv4V88a9h3n2uu0NnjwzHgvHyEgmQkK2PQn27oylE3DlksNHlot3TOgmBRGsnk
banZHMWmgKA5BIpiMaWCenwPa4sTuJmcV7aTns3UZQQMWZIt2UV7xFq3I3vGzNG63MtBEvM/mZip
EiTDdTGxQyQOVwzxhpqLKS6Pknd2MvK2uC42xek6CH4UOXUdCoAhZjJAwrUJL1rYvW5GsphpGFDd
hGJm4ZOe4ZBnJTAS+5v8aeL4JHSeAcyKgutLJw94LWWDK0cWra0f++hbpUas9fBe+3MbqnIsJ6L+
zo2uPXAC1MbzPT0x1ad1UVxMDnOM1+c0sxGxPplw8FwnbbREeY0nE6LceN8QJme6ohppv4ZxI50s
NiFwCUKE/Y4oqV4hh0xTLQcCjDlIED0pK4UaJDZoNMSt+K177dCbkCfAlHgwsx2vzYNG7UbtLJsO
GX34r3kET9RUAWqm/8B8/VfmdNFN/IYusFlLVL2ZyCMAJT1AX0VN28drc0ysJ4nWaVyA4hkp+2hV
vuuwnzFDooDO+PdOQKqK8elCf/GxQ/SrrQK42WyxSz2xL26D7EEiG5SOmpaMRt/wRlqrNmwpM9Z5
na1b0Es/UvixvpvwrJ9TM/dSV0HHgMRddwOLIIprxR780BfgT/NJijSmwfpAhe1kg6D4IRvvShXB
S0ptLlfZIlrVFdGCok8pl0COaLq25kfzKgJetGrvHKsoHcVo3J297h8xsVXa5TRQsdDwoKHZJZnA
6CVWVW9D8XoCItwQINNIbZ4VL21oHaf+W2YwzE2WmHSommuyWdCjH6lxSR37QVDJqFbbcUooUnib
DGtjT7FaWz1d/Ug7TsjaNbmZzZDW9Lcbu0k9vmth6RiPpgEAj0UOvC0bmHtb6YbzGIfSh2DAgc0B
CGv+vQIPzcwbaZ1UDVuBSHANoLqLKR0+oVGt2xVWc9GFXKpRZVDjWgsVnJlXAkSvLPLHq8VysKuy
Uolo4V80lih0tmXcaem+XUil6IDxBG/XW0aJ4x7qKIprJ8cxL5+QcASQoaY7NarywrYrwoaV7clV
z13ypPz5vGhbNAnWYhq0nDb3b4/g6SDRIljj6KZSUS6Ouq+zb+Py7VSOKw8h+w9YomfBp8Rs1xsK
oF9VQVJIYgAAWBB/QvkvxDuzfr/BadVtZPoTmj1R+Ke4kYFjDmVNzVs4dvzWd2a/onYwEqgWyFBC
HnwD5dItigstpkjdD51lK5az5iJq50qf0X8BIs4VPZ1jZ7wi0QLQjq7gS6b9t6/enWgTFpMtcYdS
ivC69Ep+35C7+IhtAe1o8TPVVNAWIZRFbdSHxwAMwAavWrqBe6A08z56vOMgC4EmDlnvovl6bQoe
rsgOytT9mGdH/TS5j5qmEwwHL5ejN0Ea4p14Y4AZIsLpsio2AMiLbhGR04/7f44gbP1ygORbP/GV
vgPB7+0OTs315i3G+dXI43O+6YmxBECV3MpIr0XDY+CfCs4U3VgBQrODpKt8vFjfGbFeznifcM/V
Biwcox2fiqMWMG3Jt0hXmNPdaxHQaTVrMGeRpVfy0GngvWzZ/MWVjOhwPM8B/2jJTMWVQ/YOjvbx
3L2BT7edHCBifAfK1ZBTuZ993crpwKQUjvLEG1BzpX4x96Q+iDulmzmuTLIeFnpIX5uPY3xc9jDY
FG+UJa9wvIJnAvNycE17VsNX5fgnn31Sg3K/mwFqMqScQMsK167CFebZCEI+npSXyT3mvLQXDnjq
y8cnj41YNlCZZOYxVTWHWji68YwIsIL0p2KNPFXYSC2PFZMopKs2fCfrWjkmmfBw8I5qXYkPPVou
KMuv6Yweb82IFxP46F/snRSJynVwf8SWslnLfZ/mwNdHuGQm4nqCd4uHYo2heqxCsmHTrKI5m3XQ
sLtkrkorhCRXv7Ao7J46GUTM/rRngYB3HVc2NKiyRkIEVakiSXIn9HlKA1bvrflLAO/vOdqZHsQW
qYAd1SrUm05sHmoTGpw2ZukrGDLALeKmj4reJIbILWERLclKUNF0QbTrOw4TAt8Vthp33Dao9S0y
BfkZSdDpu7775ivOoHY+FaiJGQ3aByqTgcMrf7GFOw0bPjjdKtFaKpkYp04oh0xysDdv91917T1G
NlysgypNnMwOINGqRJNBtdNNBdC96DJ634Yyl1WoXwigV31as6+WfN+Nhyx2RjB2vxdHRg1s6FQw
DzNF0SCRUjeRwh0QB3KFJUWOJaumljqwSXAzPrx1W4oRWebXuknf9xP/O+FtVBDydKM+NjJBUmdn
JpnDKiowFnDuLOkLdC0oahZPmCQVFFIwpkuxGdeQ67Jutjldh2oNNQhTr6Sp3nm8i5RbWRk8UBoX
7HMNhz3f3/hhl567YXoEibNtTVatpUfs8m3Rh8+Va81m9HRwyCJzURqw4Y4cIomhNIZcjk7fwwn+
wYqZtQ6i7oQhIJtgMxtDwHkIlxcgAIDmwAiRxMqE+i5JKglyzNrDOn2IPVycai99wrlMQZ8e8I/i
tNrILziuwDzXpADOH5UmJwjSac77Pipw3sD8g0ePlR81TKJ8yS2tpDz26RuMKUeMqLPbUojic+PI
FdWZibM2DwxMorTxWnc0fI9u5/5u+nvT9zw+cUFYKWqKxxCAhxTQ68rPUOjUsjZVWTp7vuKYynhg
9hpdmEujsevSo6WYJqbe6hGyd6FQdgKU5SeHvCDWDUUs7o3NBOiOZC2tO971P0DI2Bqw78NYodZB
fOSukR8LAZbFBfKtCYD/GA1q3Yu4PZR95mflUznPNXrxfaQF7kAcr1x5QBD/yKRV9P0c3PrnA3vL
hpZLRanDiDc6NBTPbQojkWwpMD9PpK+fa5+Ep0AkAqGt6yhmIOqOIAsOR5dGieKkjBqctj2H49CX
mOwcrqeHDRgCimzDTh4y4GyFIZCkCv7W+MCp/J5bQjo6ejpXZBUB1d38qV0jsjrnlNSxxKVA7gnq
eS5ujShXBXBTDrfxfaUY/s/M9xu7LoACd/CW1nwU6y1Z8pNq2TImrf3hoFafzNXW6mgHi7kBvfkS
Iy73imxa+ddglebSU5+KUr1XsAYpoYlAvrS3sXsEOMzzisC8LqvTWh0/OKh0d7CLptRTqiHO1e11
8yxe2iRVA+fQ2iTzzPSnQyFTraktqWdx6Uuw6diWFhLhN/cypVnEl1k9jzJwphC136yuPhkZDuq0
UXGMFy3kEL5OXf2FBGYL0X5UHCir4WDxR9+ozyg7tMSBByVe15vFj7SE4RQMAM6dHX25wvrTldbQ
r3vpe/RwGu9N+6sHE7jLNSpkuKmAqdcqpRBlp+ZARUmABFZ3LXccujDIVOas8T+bTrCfiWwpgHkJ
PqO+jsfWHlj8MKQV/z1dUrMNBZBese6DhKFF2ATJrO36ZuWKdZv3cVRYWIN9OtbSrMg1TdAyNHs8
Qr7wvVu+8Ma1LN7iRheWEcAYmFtC7sHDYgVJ+OA8yVvz5GCrxP4VhzHwseMYyTbvGl9c2pD5T+3l
W/exZj9pd+EcPPRuE5KhVZtUPWGetctSJc0MsCQBwaxJo/VWBd2BMGC23UkWt9+RkfoE+xs2hTOr
QQhJucQ8LvgW3akw/GRnPAvLD3gFuIJ/eEUmzaazmOqj43VHx+BazzY4TeBwFKcv7XP9fI8zyb/3
5aOGZdc2/tW9tV85661dg414K2Q3ObwesQpm4TTdMS1d3xGU0axwu0cuDCegek2G0ZPqn+tBqtgh
87ZwJXFE80s6BbVEUukI8etx30axF7WGopP6X5JzOWBWP0FgWtpJ5ceOq9jMieDBQ2n4PcA7iEpR
i8WqbV7eKSkFumKkFN+wx0zFcbyFkDWUNcgGBgb1D+ZQKxcvTs8pwiDajeiQoUVerpyScil5VXd7
oU2vjXNxpB0/CWO2Y0K8MfCB683EVPG2agJdiL2sE5uSo207/5lxTQWCkXfEMP6ozn29jbkjAU6G
7E07JcLpaBGFj//H11yi8dY3F0NDKBccPjjtiWRac9zbUr+xw+Tz0y4QBaSU2g2FD1PM8SrG4e26
5lsDrbe/yEw2+JpusJ43IVzKsK0Yb3GKfiTRFCnGnyb9TiY2/7uC5OzonhhiowD2Bi6oHvnEeoGp
QUtZER+WP67USRkXZRtLzyHHhztHIa/hDgCwE5iCy56+c5bSe8tg/dsAl8eDUR4zugA2THx3+rYt
/nxTId9FnXpnfPdi8XDl9kZFlIxx2UdVgW+S9RVKeY16flaII/app97kHblyghnkBV7+1tsT3pah
6EGb3bWVWFXQhacQvG6MbXF5Q5D+YJXGFORPxO65zbfFcgA/bESZqzbD9HYnbkux5ROAGd/nxRsl
6AELnru3I9p7Km0qmba8E+3yKVyOsPpFYC8stHhGHmWZY4DIHDxUvee7XgJsES6PkTBsUPn0qwKJ
gaV1Kp7rWZNNTD5Upu2ocSSMu8vLqit2VykDGbKL86oLk+z6q7JgoTAOeAAnjO2RVJRrCFF+Vuq7
8BbfPvkrB0HGsbMbxDNYR/+HwpnZoE0BbdbPtDcSuCO484Q3JI6pfJ09Gd28aHHSbqzhH+psK5cG
pVqXEd7kMvDINYrnLTbggH2DYsa6aoB4FUKfXNOC28UB7nJCMkdJCOq59owWt7/Y3dOViwVXFPgT
/yzZ2Rwkz9I3ZHptkzgPSlkFAxOxpQHhlKlJJVqdmV088z1Bf8oJ6OKbxW5Z0ZAYCMub3B+/RaOC
bfTi6p38PkwlIGhOY7mFjh5Ex397Y8d3vZs9gjmFRb/YsprRoCOX60rvCRr0f2jSTWRZq7+kIfF3
kdA6NtEc66Lnb3qH6hMAnOTWj9s7zg2N6xORZgK4jl3ecLdNV2NSZoGmfdr7EsXSZZyNb4j79ryX
4YXu99JNZGYizMnTCGklS+90iY6FaqNmiB5JfwcNJk2kRPEZ/6Ap799vj7ENH+/X4XyYmhNFwGxG
4H377CLU2Ht9anP6iRfNtY4Sg0i25TsCO8V+zNVWzSKdPV8l9w4Vo2TWx6WQVjD6Hq2g4z5EaQKx
H1vZXgm8W2gy+7wyRULeC7e3mPH/lGkfUpskdk4vRO7mQIG0vj0Cb0AsRG4OOkTEkRkrYUKq6yUz
OxLQRKwRa+puu+4t3rIuK4piCne6I6BJZMLIdLYftS3ZI1UnDxArR6pFIctoJnbUqOQQRXiDaZ8c
y3xn6PgHdV4YbSmlqux+7edJWZr6gUrZoL+s3byDdDUFM2UdOvBx5go1k/uCx24xXjKR6eptxci9
gu2t7DC2bjE9hPHXallVz9JFtWYTT5NuPMRgwPQD7rB/yAek5SBEn0AsRyZLYfW7uyXXQadG8tV9
oMNXt9hwCJs118FbL4nJnJNTg/DMAUA5HaURw4COAgzXgDZur8e0RZlizquNJtOD8s9tRfK5zhle
qmiQXFHZVUubz7TR1jKz06X/hBf/9M+FHmyq5tr1hsfcoF4aksnL+h2C4kK24VCeiyBFx3ctNt4h
rszdw39xi8m/zIvNJeb4l77CDxcDqrGeKgTBjtNcV6LLFkrzhaF6l2IDBPnbjSay6O5G7N89cIFS
Cq4iERGGv49KygbT8UyN7gfAwAURK8eXmwGmQH9vwPspPhUHy1DjBcZkB7LcHtB3yZ3kUxYW7i+R
ras/V6KwXlf6A1BZSKGz2jQZ+op9xJaTDIIiLWJZStkWv+e1wwV7SnIpRVqFgEm9+zdmzK8twgqp
lUf8QLvMMLZx3rwH9CrisbCCppRyf0GxfYB76fhn85TTiY620x0wWLO2PEbEfPWG1rnyZg4l+ccQ
c9BXigk5crdCi/oeN+2x0Yq8ezPrAVvyeEzDjpoSQWKZ/cSnpMPsw3PjHUARt3EEuZwfhXUzHo6b
WETJA88R2ISPvtdzhZ0AqQ8vRIzABOKGJzZXJPS6F13DFAKGc7+KGd8ENCsOO21bFDGYrCYi1EBy
4zZme7tVA0ubGCdI5jntEh63fNTTwu3Wxbo+uueSDjSrwWR3u/EfeiA6AKjdXwe3/aTCe6HK9nx2
8IjOUmkrjPXhskw/QIeUDBj9KMoPlPbHbkNaDM0yUZGgTvw+NZLIfta2t3pyH9+NZjcKUW3wBPKB
qDwDoXClph6nDZ5JuLRBbmR+QjYSlKydqtkJMjlnZjy4poXVvn7g+bMRLG0PYx+kr9NnLLXDi0zS
3NksFlHFqSEFCsP2XvJsZY4bbvQEY1fkM+NCaFEvzFc9CmnxoRb78mZFtZhQIDow2yQ7Yb8VTTMl
XL64mbY5CbNyAaG0l+olu/rBaS0T8s2d43NejP33m7W2XZ+gNxMbFhNgXJUDc31aFRM7q0lIE8eQ
DY4YfkcrMOXs5ou18o/n0DvmE8saCR2oXdTn3xoSTusIQ4ZRXkCRDd2GyOJr45CghfL0rPVGRsoo
gLVbIJYeZ2ug2I9wtUPsS5Nz5OetpJLQXf1szuFZTRbpZKE5waLva0mg8bp6aSbS4HIi1MxnnUFb
izw1gE8syZ+g3MYc+LHII51Bx0YQ8VGXgQoIfezbi654eaTUCAprMEdlLH2gmRDpT8NfGsmnugy6
820iapW7dyWTrxfTaAb5Jo8jJMqcc6+IndNdHb8sZnHKTdMzGzyq3p23kfLR1jcw3qN8gZOPCdEL
5paoNat9BsUPcndeEgV57qfV2siw2bBp1Zy3U7mgXxp4qi5QVDSqQ75eTKQ/PNURbWyEHdSmkrT3
LW4V2zpRTl7KVxl9geL14jk4IazM148hMLu2EoPFeb8n0i7BrJRc0nNKJFgXCKnJcaC+OD3uDWs6
zCSTa0KZnS6AL7oGKQDTHhSf3i2x96op27v8dY4QknA0r8FIV1IagBASZ3madNFwfGrfD/DhFjhB
p7sp2mk8gCsYuNm7Jj9Ii0waAlvFZw0RE897izhJw0DlJ0h6TUYvEMrWz2IekFYroVrQQAyEm4jr
gtO2xVdJ3gBoNtOtoAra+QF/rETjztTL4oaiHAISAT2L4/EFiG+ZApkb14u1P3wQx8DKrEA65S7r
bWGfeONp4vn+skjHBcPO7SxDn5GV1671clXdEsB4AI1/QheZuR62kiEhJKij/CgkEd3zfTHofcAA
jroINPVNy3/6uvd4rGXsDvaueAjlzmjdqx5ub2NmRPv2GZRPZ7ixSlzw/IXPRtK2Y3d+kzq44mVF
qJF1KGixsW7FaaDyGh3vIygdb0jIBrHnyrgFvtKSmHJ9TrA/BkhWl3G7L8ZeKm53sZEN15ZFs7qq
79+cqi3vZ52c8cOgnuhZBYuO/H1T5rypvX9VVst3bUakMJ7UOQ4Z/rZslsRbLjcRvk8mMYHKA9k+
iHGdhLgvIF1390BLZjFkUwTKgY5cla3V8PNuSIA2bET2rfEVW1yLgaQJnFPYq4VU02E7QVNoqY5K
3FuivIXpWj+7/P/0gNcdpEHzfCNY5Fd4Hcx6iVn9xEuxfoPTmjBBeLsZtUiaRSUn5xXCQKRciGAi
DoT9YH+51S92M3+h4Z7fiw6VJKXJ8cNRZNIcySGqj8C4j4uCyq7ln5je5Iuyz/Y1xYK31Ui97r0C
i0R9V7cdv2DcvIk7+7QEoueRzpwxStdCpeNNJSGTbM3l5L8ycWa6f6R1OCOvsjWngI0LtFNJaNdB
o/j3ogIEn759/I/pg38BX6/9hVvxHVUS5IQOJZoaM9UDiswYnm9vhCT6oeGmWw78kHy9ctLlIbQ4
/3e57FZV3WFgRhCs8yzacfD61uqL4Il9VMYQQ5g+aUq04eBM8dQUmz/TdyAG9lHrPi1qxL/eL4YQ
VC3hO8/zQC2hhY/IIW8a8ig4PFmMNL8NLjBM9tJeh9qqdFZxD2ds3oiSXb7aGggib9KQnhCXmSCC
8Gj7CUxMcthEVKjpT3knz6C6G934jCOHad5HWFBp+q+HtsrC9iu14Uuvg9J2kpSSZy3KLvWQbVAB
0+LfQQ81cSqyDIUycCNRo95cSBQPAYd5II7xmbX5C2+db7gkj/E//cUR5RTTLTEG8j2ovGx46hBa
pTYtAHWUMh5m/VsPvCNT0jorKKngz0IxJ5RD0nDYfpQaFRq7Npf0mqJ7SB9M2tqyVOS4FYtmT/fJ
Qi6KvMb99Kt9w4hHTHxk4OR+hgLzSHPLhS7xv5We1VLa7mDo7IEGr/ns8l2smaZcBaEuRvxkXp9N
WOoQg/2gc/5hsXqN8fP8Cueasux3zVebc8vzXid/OS+VMHmo6bcmVw/LNGRSXId03PsRwTWjkAyT
DMjTuPJuPitG12DJ3oaz0jH923B1KAur1+nDfzT9ltGzEfuHCuSL6r/c2AxR3SFV815tdESHimgr
oE4p5PIpIV6TU9dQsso24v/pwi+YvzVFo2/+W/nWlrvsKTk/BwUxUVHKdM2UHnT+j6DZcHRXG+WX
UjY6Aazm9RM92+ABaN8nZ8FJ4uWwlDHzTNmzRLQYs9HfdrWJFoCNDbYxT4Y+fXFfK87D3caII5EF
yoipyZZm9QXFbkr+dWXYm5hrqueif761dRDDRvbwEoNHjNW16xmpwMW43lbeQ1DzAwSLPpeNdXZ/
gbyzij5wC4fTjwQmNj9apsd6s6MzV5idDt6gAxVowDXTEtsvhWmwQtk/Kk6KYarkRsHaOY4O53lx
33DxLtNbmOqr3J5j5bIdgh+PsTgVN024FyqdE947wJUT8XPwK/6DXZWYH3Z3t4VNUkIxnrUUIy0W
z061CEV1PAfgz0daGADgNVnUFTRkuvP1Ir24baGi2MFw8FjAckBsCHMDm3HVZf8llw8vLE7xJLNz
DznKbnUJY0OV6pY5o884ilTD/jHN32WtKCZCJba26ii+cmQ/PX26VKSlQd4c4cSxtMjNvo0Z9lW1
Xr1/j+TqV6OmB76CZ6CAi8+sx3UPzdMDD2MZ3IbDgP8aGE30y3t1t3binvoNgtAkjxSQDw8SKuRj
2t/LMR8nBJd5ij9pEFTsURPkw4oWkANS4+4zVjiTaaM0LSRyp5OqRxXyZ/k0XoTQTSsa5EYfH1Br
WkaEm4asH5lMtGpclzisToWA3AWEt6B2Cbg7HAWR/ZKFkqeQSk/J9Wk7mZMlQZ2l6ZQIaCR67uxQ
tLseeae8pq0alt4HRmmKtHr+zobLzPVedU7w+KYIJ1dfhys1SaOZj3vHaC9EoIJ7oBEA89kjefXN
yOAX/y+L+LNqjyma9L+2T2sd8Pn93G2liGz871rhI+UVibehdnribOyZH3JLwkeg4Ox015a1XYHz
pj13zrAkDIXRIaAZSv7A3Xrve5G7lbRbi8wFxuJ2yq7qSG3HYAhMvGJLIbZNbnMTM4TASCziCeM3
JTixTn+wA368I1hJAkn/M5jUlnihrKU3Z9ESUnxPbNOgXiq6E4azGQ6MQNuS1Xmo67Tn15wc1KY5
kwML8xfI+MEdM/qGprOukra9AArmD6+Lw7XGNGiseczRmrdNRK8a3vOeH1tO8qeHpil0lpBwc8kH
SC1yn8DdOSUGk7HWLDUUQSvT7Iq7GIAa+pRi78gwuVMFb7iSdMPmIn70i0sNJhOyWAz8TGOsL/N3
osfVGrx4VxhaAoE3QHxDXJj7NYPQQ3pje3goll8+GnS9XHA+GQCKGIAQRfkggRwa7305I9RlAco5
AP34vkQc0bsj2/VdfHPkp66QA5WZUQRRdjHUbOOjEBLCWdBu6p3dFio9DS9ZqB7dEKZEt5DZywzJ
vFOmlxc3rn8fmUocVwq/pVfNLSFzvkD4q1dMRqcz0HQFe6yvVerpnN7/yA2C/ea3SKIB+A7Saln5
lAX53q2cydwrbJQnxqO/aWuUsqEMwzJc4ETvJnyZo/qyrKciouY7p70C+I88WBiPRWdfDvTuAVl5
n8OGaZc4MS8vOV+j+9LT8TfazfTH+A/eZfrYaYfXLb7jLN1RDXamVC6ybelcMlVthMbRL/BKZLX1
j4cp3dz3C6lL+cjToRZtb4M9Z1jXWJ1AzhRkg/04KmY3C8BPqzYNsgi8N7m5Noiq1ZZse7ZmjL6V
XvqfpB8cv+QPz9leWFRn1tKGCd3cP5EvHhVfHU8CzBZ7JzuH8T+l+dYPGHNeLZwMAriCUgoxUA2M
UJduP49vBNgclpsi3fM3g4ynsHw/qlu2KdFAoHpuBCEoQhxarWi2Nxkt27YrhYOg39jkimltQJBC
tqW8eGTsGwl+yet661UCXyCaK3AUwAIDpJUzsN8Oaij3Xi3LsDuu1njQhECL4RO0htkgpUpJVX+7
HdAgOuSo7bOXzgZISRiZ1ehEndv1dJrz5Y9THQbX0imkNupdrXSzE3UAUCdf6is5OLfHfGqfs+am
2ycAKs2rUYs4SCy6y/uqFFxrxp3HfZtibKd3DPytqJ0ddbhJCSEsmN6oQyNlQ7Sb41WxiKWAfBnQ
cVQMTvZWXIlbY8pvROXBQMM+d7RdyhuPtfdcQRqjuCybxO5qM2RN3d+AjJJxvy3Qj55DzWMo2wBq
aBWwHO8Th5CNJLp9quF/AigwIpIHK7Jbmsb09Jg4Ce9lQMmSRYhXYVgq5cSQwVuoit0uwJFG28yB
unFm8D6T4+8LBZIWF7LWIkh6Di4AaHBeLjObC0i7pTkqZiXNUiAjGt56vYh1tTsPpoeDNrsl9eqi
Ubj1ntjEOA8aJf6ZXcpCf6ywKFqzM85OkaPOHKU2GDFPMk3tcD/90GrizdUfZwy5b0yJHycOi/dw
v/kPNphx6JLniY9MdiC3M/+ObxbUoLFKbeM1D/n0dKKFrip9ni3NeRkbDyMXQfkboNKWFydU0SU9
vle8GDfD5hwzuIjDgcq/enQ/JWRegF6T6C/t0ZQXt/DR5yoLI4GyGsZNaVNb1xvN0zVSc2/fwyIP
fBp9bnDHLd6awsZQt7Xr9VsWsWGXTJ0RLyaEfpJlrxug42uQ/bH9hOVCaTAa8t/eeNKVVKB9lxGV
4FFPkWNgrhJ6IOpF3jYC640J1cJ1KrpBfFlo8oBn4WttOsvPnWuF+DCZnvDvjzpWDl4VKKtUjRsj
f8Gp5a+AxMNKeEBjWCO6RGfPD/lsYgbTX7VgaOBodWDtx+illaHK8WOrtt+E0gkRX5GDcli0KlpQ
jOqfLp4xD/WMW19fjaBqil4K/VRRwKH8gzVQ7BzBaXox/qPUOAig8vFz01KDSQUJV2OhMgj1HNkL
iOsLbWheHGjSKjky44qTKCzm4+WIJDXJ8gO3V33plrAhZTGsp1COzT+wPfFG+mISRjK5Rm07CY5e
d3L03JB7wFH65biyiZ2bcI1RWEKen9cSOH3qfiaWJqoQnChhqOy4zYjJRBdnp2/Lx28A1xshug3b
U7DR8a2jlQnoqXlX9QXrKgy701lrFAoceqMnn+D8f7VI4UGCau3n1m7vczy2AmGB3fok0QwllwkJ
Al/CAkwjmIBRLn7vX22oL339tcHEw7AmJYE7hQliu9R0yRhJT6cKNbJPU26RhpMkyi0AOe9fX/I6
KGtm/cPEDXE36I7YIPYNbqjlf9qlWzg06kHRUYGH/D2PyFSYvuJSclIQqpx/gmX4kFSlWmAjXUT5
t2A4FcbJFG83pN0pVxFqoQskdAAsYifZrrJHT9Lq22onMEEq121MDVmQ3OGOwCVP6tVDgTL3Q/I1
1gZS4hPCfp0TYWT5pJ/StBQPbcKzOWvgeLky0b4amwxXpumkQmbaKsGfC+20WpijwtXxYjrn5Ph4
SCaXD9XOIOBI1Jj6kaLMz9fxgaua3V6RJuVXWNVYbiLhRlnTJ4PZ77q08uqdBfFfuntISHen3cNE
KJGQnyhiY9/adXGfq5CxDI4U7mCNh8WPASLYv18lAdjwh97uxNnBbPLMOIdTT+lUBx8LYr2k+W1E
JDRh/MsBA8rNcqra+V3hU2P2QIJ9spXopK+0quu2O94xHRtbDpKBkclVJF15XSYeHexN/5niWNFV
JJnxS02euJOToduN+oaTcKKKI/bZADvF1OLjrp0821Halkru+lmYDROG5YQ2kqoRAoRUV/yuXfmY
hGhfFg3gFFUQipSYMFCDvs8aW5hFdKIlhKNH4T8u7dTSfvX83+frP5UYC1jHg5P1+USI16R4ieAx
k0CLdRN+YmF6RDseEk//KhSEg38uRsJ97yYu3hvjBP6KIDE65fqdEfEhoaHnED/CAF1rlePx+59u
eQeCN2ol+TXyrKwGu0xICADnn2SJPeRee9F5IEvmKFwRdxDSM/L31Xxy01rP2CDyERXMYuA6eTzR
6Xpd4dYoueZ0U3to/6kHL2kRsjPLpUTGV1GqeEQDXy5YepWrLZYH8YMZF1UWKq08K4PSMr6+SyHW
QULVYc3QxjFWTdfCRodLUdMLUHrzNgDoc+30kP4jZ2FwVIyXxcTQ/ro+FTzOgignAgoJRbigKA9y
6/qykDgjbam8nMCVw+dicHvXLwR54OcOTuuBJ1TDAApK3gRffdC1fWTUQgwnVhIl/ZdH1L3oZlY5
MRj0qLk7lvC6IRkZQ/V2V7gjsmP7AIJ0USkHUFYns3utMurMAJCffb9g5BCNoQOim0tHFiAIFLmq
BnxMN6SHC3fcqSycPC25YbBWXm3hWVdSaRbAVcfxnFkBeWEp71AdMAZMCvaRlnyncC2+6AaZmjPx
v7HGDsVArKCUYEbfU+BNFFvnMYMyKUDZ0343qAVv09di3x1TPaYca4LVnSZIAlE3oHPFNW/UTjt3
OVfXVIOJv/L2K4elyt/Nrdcydl7mB/fU6wwDAUuOpVyL9nuKEWcvnnjR5FK8DtWbhLkOnanCYZRG
dFcmnVdqsCPGIhb25Mu3jmLxWDYHu93tU1z9Me8Ugl7EXUI5vcgHul16HNj6DPfCeAErKPEszRL4
+I6Y/zn5/WloCzBxpbSGgzcUZMru2aC6LRfP2VF/wJhRUbNzQOWDI5ozzohW4omAPf+QRQQ+NTuo
tgt75SBhjTFCn9NpsUFY4Lm4dNiyr6QbuCb2s7FGtR/UMBdEW9AUAk34t5sM4vHmS/ceT9ypbmi9
hpYIzjE70wv5UqrAoW0Uo6okkVqy9ZmU/NUIj41cFBbRtbHmrjsFYxqmgvpDxmNYnwIHcveipJAV
KvjW6+OhH+D6ctFCC6uyfM7rqZqbN3WR2TPSyNhvA5tHWgr+NURAVeCurPUpkkuim8tPBU8C633M
ZzDZ9KqMO0L4rQ77Dojpv+Jwkz/m//ADWpJE3QWjACmVQemDjXszM5vvI7Un0fEPltiAHRVQWDVI
FOFegCDR+bYx9LK3H0Zy6U4H+W7uL+AY0x3vpRFkdl8q/YgdH41swpEVuAX7cuVHoh8whoEjWAtJ
NSUY6GCU7qQgxQuyfbzTcHniC2ef8uam7sM/quFg2/m6oz3ANPWZ5G6OOxXY60fcGrRYBPB1L2qE
l1COD0/ktiBiHopTABEPKAgdI9ZOhifRvji167amC2YTujTBCwqKZHsiU/Eg/WrF7PgJNlZTkNmQ
kB/muBRfJbyDPrQe+SW3Zecdf3TwHC7nzFpnzlsIzqFsvDvJGJSEoRKD3Ohw4TZZNM7dYZw+LBJI
3Ga7vCXrUuQViCG++O/jC6pNldoGDckBlLgZ8MuSNTLiALOiEKlzc1Im7HgZWRyzetB7LimwtpGO
i5SiMX/5Bt9cF6fgksnSeW1Is0yiZwTCl3aqAkO9QIxxy63/Lq6bnzZPRijCHQ8KIaEt1zNFkT9c
SHNzEB2Wra6+pKKky6Y2VTEBZxsmRuC7iKgRGmsokmfdEb8rA4IB2sHLVOFQaP/zyo1CgpocAFF8
gi8F02jMmxqaw0H3MAPo9odHePe5eb6Juxe5xncjOXxnkRKRZqx9pWKTXMBNW4Oer2NZAxmt+06g
CHdOgmSe87ZllYeJ9BL7JG+mbaZ7qUXlHHFAvSHAjxIYXMGdAxp2myIVlIWh59MbmOZ7K5KoKNp1
NYGCYtcUhDC/SesI8K+uVxAtN5plTE6sbzVLqQmmsFXcNOnjLwkP1a+n5Gfm8ViaECRv+Ry9go7o
r6avN6fLTWk959okgMDajkr4OtW661qSpi9y17k6688u8BymKodinQtH5789mqYRN3yfajX71HQJ
Ne/IUNDY/oEaHbcvydhhDLv2YoJbPNJe7QO0dwCT+YwteCA6QhAw0IE6bE6li9PvguLeopmnkjDp
T2W4Ts1jPOJpQV4NUJTU1oZv+4FrFgQCvlYKlOXaWg6CloKUsby/NaHrWkmpUftADm7cn54kiPqo
dCwyBr2L19h/75xwyeeygiyVmvTm1mququCGrddzFgBdtCIIQyvwt9R87fSTw99omgw4glzTIY04
NmggPlxKmrEjG+YFEPhCON4Eaa8nvU9Pnlcevg/EhCIkoMd4vfFDF563FVQtJw5i2Igcw6FomJbY
8cdICax6TIXkyJBhdx6y/xosLsiUOtGrmlSer/DQqFXUVCHS7QDtbj8bFOd/7fCMBURJ+Ql61y9R
ifKwz8QtRno2k63VqMcbr0jQTrIAPXl0PtX7YiYedcIna5CrGzx+QLrYn97IiKVcW2dL9ivnLgx2
hmDLPmVCSVumEIgET7RU7mHsnhLNQCPTGO1ieVtNBgJmyueRryReZiwMz2wxeObq5ixX86urYGag
Yzt5yPFSmMRWaEXVBcyFnt2KLpyr8mc2OPZE/E8Ad0bWW1CvUgSFGRhT1i62sPgwonyc3NvMzaa2
RCECOSEPRn0VRt8bXRLqDdoJM5BKRj5ojdYlbzojpglKlJ3BltG7qtblFTkmO0eFs2fVlatK2vt+
DslUtJ3SRHsJDFjVxx0fXa1ShyIUScijuF+wZWfxuPRla4IS26BUsL33vw61z+IhMDqxYO974/aL
TV9ENGw5VicjUMBRvZgbkU0jn+zjN+jdAj/y52at8FXtAXBMSn5bVZ5XEc10EAfVtCOKbdF/4vZ4
qWeHx+0z24zkB48OHtRPbRgtYNYkFsrLTgr0MvKF2a4oD4iH9/HeM6UrxsTSPOjD9UlQkUSC7gcV
V2JiZBaiwo0tKY61LrLwRtnhHueaB1pBAreNBkZuVRF+aVuG/wr9/Uv94GZbam3TPto576vEOZOz
X4Pd4kLhEO0uE75iVHa1PJWkGKtquY883KdY8Qm/5wh7F6/wRGT6cbe216OcwW87FZRXZT2UEFLy
ejHSLKr2lrxsjXs4ZQwdmnkbigaNLEQwE+EiPjNAOZRH4KhWkxE7ABZYcPbOcOXvczVXbGstK4Uj
7zMtt7uAmQF0c5kiv78tCMCdWTqhdcGcVbd2HdTJRx/OQcYruH93UOrwzsOMDawNqMFw/7kSJwPL
gK3yKwvInKoF4Mh9WHHkml+lJ4qKzVluLr03f6xsJrgQk0Y5hvlqzD2yVq4oRRvNXICjEnuUZagl
gV6b7B0hK18c2a+8tJZ/Uz2JgqKBgTFUE9R04wSawbF8Hxu4JuBU44g13DkQMYm2v6+El2SY/BrM
NX9uic6txWV5+HI1kfYlJgdvdhlqpUvOfL5dmDqAiioG0RU4ClNH10CizqRjqi6SbO8XiKcFW9e7
jpOJkFjXVo/XfxbD7v4uAmUE8yT6Y72iNLn2CwJCMegfc/xCYHs4QkKFBxn6LI58xVSEoSb2pGGV
2oIFHiLCwkRIP3Wn7FOw2ZSpkQkIMwW+lIsbGnptC4PbWh6zcIa1jr4sU8gzFPGWeKD/1F+Q0vMa
HNd+QH2kpeNJHStC01Mxzw7j9XMhmvxFmqDDrxoXj0LNRBIxkC2KBIhcwiX4//pKFVIgGmuIilxH
l0pZIaumoO3n5fXA3BDj1b+4kTkgYrfLe0EFyyUakdQZf9U2I+9GOvdKJr2xKNEzoWAuD7qwB8bg
oPwPVenmoUHs1iBw9aLTIoegb7rFqEZFGUt+Rd9Yj1Y1bl+jnY/G8R4KcK/glnIY9fzNUNpQ4lRO
6uzMDigWUlJi3q3fbSvYCQ8nwNw2Kd9lvEt5pjQGoOwk6wmzIcLFKnli+Sh3ZOt/pt3iBtKO6dNq
L5j8ejSrkg6rPI9w3Ekffz0kDcUUonrFJlJgjh8osi0T/EaaEWwGcjLTvfBHra13ZQh63qK16c8s
wPb7//qRU2HaoJxu8dnEJu/3hcyYo+a7FxjNd4M/2BpDyTkW4/rLROsHL3nvKelDRewY/glG07nD
8f8044dKg6oBm4Yb0ltsOwtuEQ4+kC1JfnRGMHg3Y7cOHN9nbfTfX9sFY1Gt8Q3m2GNchGIX5L8p
jV0Jyq26VGtIcOm4L7yg9vDZUQQemW+1oryPtckpeHetQ5ydgaLqzx+/3L3sYNqUF7KN1Rkz9vTA
EAIhcqQrjYtqdSI7A8zuKjqH0KBsDiHe0AP+gMSOikXKfaB4hGtMph76CY6roU9WU9VGBut27M2x
+1WdiF+UGVsktWCKbF0Awakt+56i6EtxDk9PRvznT4JwBeEAspm/DUgA3Ol8MAvNDrraIp5Cm5YY
knc2dNni/0oO+U23gMf64ML6HTEEWQZrjki97UsgeN+qARO0FHLBfscxAOBn7OiEhe/540c74pCy
Ttx2b+T3vZ4pta/cX9Q9Zsd9IKChytTpDv5z+LUlu3/wh3y7JEP46gQMBJv/97fMLkPVMkvZFRPJ
mt63IecyxC18pzpA13hwZFNtFzsA8L+13P9ZzwtwdkyLVeenssJew030TOaXRZOMNAYs3GQAUNPL
WVSRPGQnbvvSz0ZGQiQJNgC0Cckz+zS1Z07SDiAmLyKd6q1Ygxcg4ro12AjHFGrO9c17MNiq5SFn
N/3uV6Jn2o4SLKaWzK0EykDeDrM+WX2YvK6IOaVYnLZ0q5bY/nFn3sANANJ5pt4Gbl8zc+5JE1ZI
EllfqFLj6pIJiIu11l2D8WbV8SzQBHI8vyAhoJFyzqFPJoEpiL5yQkBRHwvOm6e2836GPhoQIjY6
hlsciZxcls4oxwTlyxZ7fimtxcb2pOFF/ka7ekn/C7Omx2vr14eqL0GPCOR9hj9fqUY9aO2MEGoc
TTcBT3bQ9yoOgdQtGVWDKM7CO5wtLwu3+ZVGVYl/DA9U5av2Xl5tEAq8kBPjUhJb/4SvsfJ8wtzA
2aI1aD2+VHCh5M5zp6oCCLcMjnYL5An83zzpPN7aBli/RettFgXYyZ//4ZtniVzQhkGtgpT0aWKW
0E/9e/zwijQ+aMNigRAnwYabvEy3u4/E7IcgJDS/hVMuTmD0TMVSnRzIPHOaJALXUDkyn1msRE00
kQeC5y8uWnuFQlSvDqMhYCkV2VYOMhPXz54beQCG/UjnnsifvKp5L99hblk+1DZ6P8MUsCQP7d/e
7k6Tj5DXoYJhXnRdr235JYBBrLsuZ3O9aefkOZ3Oupsny5/wzz0nNs6ro2+Z+rcxm4VbCvPvjfuE
VZujsoPJPaGdZqdItyH/OVxrej/GAhuExmx8ELdhSoa/x2jkN5YYBH9PV1SlHHS1x5hkoprESqsM
hCR2js2jRfYCA1peY62M9toF9OA5guw64qWfFqwzRGHaIvmizJW6yVvHwueKAk2DQg8IwwvlX8sc
sa+ImaMoZDLVOlLpyQ1w+yJBPbNUyJL8riCtyGpQCvlLB9KvoqsnYl7sc0KTBUeJgHsRPQWaNbkW
dshbpDAtympOc82fqHgd91n2MxA1pYxgA4Uv+iRkxiaDGpEoRbbO+FnCH9SS4m0qE1LNQ7y6iMjY
2ZjQF9YMyk8/UAWuF1pHIZx4RfS3AwwKSCOCjVkz7Gxo4bU5rOmpSAP5gQAtvs/sRiGJs11pJEhS
KXvCUmP303YYjbtN9Wple/es3uyJgci3ZtXUsE2hsc4/PuxPHkdl+rHqaBtJ3Df6WZJXbmoUN22l
2D1gseBksx8fJ2LToNx423NnZ81Q1BdVE8FRgcuDDkJpxXfif8oKfQtrCRVAWjTmtM0nMPUXPciD
O4JEo7zgdIYdxMJvoCkeX9tX9xQP4VABapBDs7nZCRgDqq25HpxNyPyu4EAqfmdNiOBGFXIw8A58
INa2yWqkaeyWb317qXG8rs8yMe8c+kCxSu69XScu7hge3Wn35n+oPL7pgDSKMU8TctlPAsBuhn+K
B12pRP0S+gLq2F66AvkjN9dUkoebsHHPjX1uQKkJzTgLsbzt1/g271/82xjlT3it1ueIJ99Swhyn
NgzamAgUkKbbpYpESphz9dFO1YfYzAwpS93aqrTLw4iud/p17pU2Ae/etHAUkl0+T2B689yrNxrb
OAxObGaqgWOhQZ8N0sT1VMyWPvKMtFOyD0Ns/lenMyEs2mAXuiwnLe+h+ROuahqPhA0GK1xcBNs7
+VW+rAZ5l5K1VXYOwShX2iMBbGMPk4NIkZi8Nbo90p9a6hnPVS3q2kzNQ19LmQGQhBx+nsuc6RPW
Djn/dayJJB746GyupgeWxGHn9l/m0nBbVce85WsZrA3Ige/66HYNaeQqXNK2m7C4W0PE45OX2F4j
yG/VacuHSETCIm8XCjqVKCTlTwDLTKUPVpW3zkATiO2DG604jxtwO6WYJ9AUM7A0Pd8KIeoyxFU0
fl2uv7cgV+RPR5kTfTKiGDbXaLr+CLCoj2g2dcau0pGKFqOHmCLlK3STCehpxHgLYkA5SmvQmoV5
7N9AfcbeYaiDzoMcuaw6g5N1uKMfaOZJ8MtfrrHfSaxPehTUk0divZDdWpXAgBXv1GMwNOULnJmj
cIyN3xnuDPmOh15thRxbVs/os3jafn+NdPH2VTSu9zqDDUuKhhVgwnp85drk1yXJHUyGeLDFsFs4
j+SMQi/Fzx/JLKy45jGxh+EhO/ULG/Q63Bt/otDiRV69iDGu27m8oH0Ih1xbGZQUzIh+c6a/msTf
UjdnTLfEyGEkFzKFHP/YT/i/WWVSFpIsZJ4pBirb27g/byRQQ0MVtujaN2PVaW9JC2vQhPykPSmj
+kdHAGLIjrChGRhWxcrU0TJop7QUp1EB7tqaE4nDS/xffVtcz7m9u4Z096bop6Da8J1OGNavEj/c
Ik56otBX1X9Jw4HxL6/xVfOyK2RqdlK35Cn8wD/j4Zxo7CRgukdTDjorM4h93H3H4FOcsr0llcT0
52Y3gC1QkajD4HrTyriGWYdp/z72bgD6JTlYh+wilSTy99dmpKTcfoYIEKuaeE+8RDjqRmZB708b
c7JYG4Z2AmyODGy7hCQdlGvuQSxMM2T8GdCKYNZeG/rKIT/GlqiNJab/Es5nRkRuofzvND5f4XlJ
TdGfkBOdbloQs3LEk1Txe1uV98xOnJNyLAAAfa1xZZTvBuc2tW/6q/sLrA870Rx3e22Z8upF2JIP
ydQTwwHubmfVlRDD1F5YNiv4O1SqqG/lEQRMjneNFMYUWa7jrlJRGMbraDMH5llleusuNw05fppj
/08Pmhn+kVRkko2LqpgzcgsA5HTQst+s0lo0rmUZfVAfb8Tzt5YNtbd/b2S4gcNi8uprBktjLeSG
mrLrhmIoa4kpxsdqKqE/xj/zcI4hNB+3ji4f4DmD15l+2z40UKtYcNN57oPyRCYfG0ZvSRvAkYzf
hr+ItA+0aC9YJ86sl3IKB3/Giv3xiEwdfEPJldtQrKRQXGQizBECc45FDguP9R6h1delzLg5PmeK
6tZmYU0TNzuHt/hAKshMdyZUR/+WuaZpbXRSjKIcDEAREINy6Qw+OHOpHW+P7Vcx24lr0ngNTHlQ
Due8WEWSa5utY3XCyMKYghaR6atymgGX4NkpzjW45q/jXFFqKPz1D+kWAjwpEnbOUwoQvUj4+HcO
Ad0nqOTkGws+x+RXS1pubxPKrLJZGsfTdCBTe3ugDlBoWEpz44EiEmYjJqTa/waDNGuuMbL5yevf
XU55krh1QJR+POdCzpIbDisNUJfPEaF24BLFpNGnubMDlY3ivABa6+N5ymAEGOULvEa2KWjS5tBs
ri+omq4bs83jc0VTKSEBixni4gwqJDBdUdGmFsuF6QOcpioy3gp+NKEF3VUqXzOeCHa5fyZ+4Asg
FmOTmY1U/4CQtsknUP2lsk960cf4FaymzzaH4zE+F9Ikn5K2uTmPVIap8JbSE9/u6rgZww4lR4FL
ISmP/Q/oA6BpoLXxvAvFnSnBej8FYOMPy0CZ06Dim1pb2jPS54xad/73ITIMJtGhXM/ZqwlLNRh1
TPdCthiLPCQ9wy4CJVmfcr3yBKU4qw9FY9bJuBL/QC0GzBlysejHv42lfxptNdacyuPWhaPz4txy
jWVhi7EhkmE4dn0VzX/dkGRME4+RbWOyriVCXaQ2Fa89vKpvihtUeh5dy4MAgkfkKkCe8P2qavFe
MVEnclR8LqzFlpird37L8uM7TQoH4+7EEA3P8OhGYZ+dz3x7EvxI4/0W4aCw58vUGVdmvVIBw58k
CjPYq3npEl16WrBrtXdc/sUVQeYMcBqu38qzPOpCYFskpn2P40JvWDrG1g1bkI68wBQPScZxDjYe
Sm0544W3Ao/6peUdojKGES93H0wyN4rUolKN6KUzlrKEWwhx+h3CnwQR7qaZPBv+nxUHbNJIstbQ
ZT666z3IF4Qpj0AO6YxZ/7lnDO74USk009Flzr2wDw+QxaNlwKzvbk+ugPdH1q7Rbq1XwJMO8Oro
wgq/Kalms3dPAGNEI5BfkTiS8CXRztfHbnTjdRC4mGCfs8EhlqGjBzZ4c7ApZmaTuer8qXEpT3fM
h+b+hrt06jyp7CjgBq/plIp00qw25kDP2qIHVAy8mA88b5r2IBq+vZX34y4hMQqF77g85I6jxP9T
Krdlp9F97V63nVi4eVkWrD4GiIp+tmkmPDgyE4aRe+0ieFyR88xXLvsznreii/XCqkNcg0BS5n3t
xGg0Vb7+WtEhpWog+uKaB8AjmF2dPYkl5LnlJjVwWb1tiNFV0DYA6ta1uZCdI+dNHakkgkcXnpyh
Ad+ODvBQ19gxpbOzo1AD4LGfj1hK1fEs7TtuxlZFGkN0HRzTJv+f/NUgMTgIh0oWjQ0D74W7lAuV
HQJ0QQPIMWgnNj2SPznGKP0Q3/ln6hwFrTIR5OEE2pUkSKK8eASmGysdzXuCEiX+8o0pqjnkODff
NPOzP4OAV2+VpQaPwDOIBgUccczQWyLSDcCRHEBQ8PiELZo2z2NQ5Itl3IfRjusMPplkdIz4g1Qm
4ruPL2ZKJYGpBeA0Gr7qfQb5G7PHA5HNbW80Gb+WzX799pzFPoLkZd6ozeMTtriGtGs1y4Nl5awq
G4F5yDYnz9TBsIGyHZGijB0BGbshDcV6dCKCtDsOVhdzWsBOpGzBE1v3mP4FR+7zGCVN8FCSiPUV
VzAn5VDe7tBn7bt13bUO8mVgRwrJON3dlofX2gaC0tX1QfkjNXQ4ttMHq5ncaUa47MqEY/ooZm06
DKzGmoed5SBp7Dzj/j263LyCxM+gHkmi2yCGrbBl9qbSJZQYte7RyeQDYaobxqKMLiY1Q/aEenMY
C8fRrXgSTWLqNiRRP8yFCN+Pw9WcfNHHnMmIVkFQWsLEs7b1gjFTGZvbEJQOf5Eq/5rLwYIM1KIg
pv24N0ujNHwpdhavRCCSA2M3tt4tOx5PQ6lp6ip/Dw9mZXwgRNzUbdqLqqdT68Iv3HflMVMekIrj
GrhZVV6rRnERjrqjfy3jKsptTfgN8h8iFnIRNVn4uFbZqcyhXUle3BoqYgm4ScwCY5Vdn6zYwaAy
klPjcM5duov7ujDQIWRK0MvrknmkNU5jrPX7+92HcSyI8cK7rEssnf90uoE01ANIKp62HGPD9v87
/q0+Kg+VJsx8/SAPLWLoSPAMiEZYHEWD/26HsFhtv9kwISpS1B1n0Vkjer6+vj4KQsoH/1YzQxjC
lYK0habqX0Vt7C+2ZJkZuSGIHFnRlz7dLRSWnyQHXMIkG5giNydTknA8HvAd7YNUewbIgmEabVCu
CTV+i5QKJ7ihA9vWuMbKFuNFZtFFFrmI2N3pc9kDxuiqHjFfwtJk/ft7D2Bza7POi1EWKQq0XiAq
+vXalWBTzEOjW2L1egCFf6o7973DNVK/Mtyh2/kK1xLkfciTPzRD2LRzJDF00m3O4xcsfbVJBL1A
TLvPGjBXI81YXiDX/T+2nrmCKsxg0mKkSHz9eSSn4BNNMXiCi2BuNl7S4K8pYZgGl/6XzFrND4Od
RPnl/ilfpY/4ZhBRDK+ug2bvDvgFb38/iqQgXETQO3qAuDFmXLxRC/9OUqI9T/bOq93MeFW6atah
PvsyUl+M4gsH7uaJpkPkF8QkDkPmjz6WOnmSbKtCM82cAfbRi57o3xeobLlze7M4FFxj7muFbO5X
tNUqMIBeTACWwdJOe9mQBr4Zs9ELlqlvP4PstKdy40G/+x86nF0y1v5WA0+Z1pE6ehE3hJsgZNhn
6+kkUVshPeXuwyuCQ/Dy3+QNTs9thNj4T6fabHhSNQrZgcHEO1u6ktuKJac6oEN1B0BojfHbXHOn
Ww99ud8TpRJ8CaqB+Ljk4lxja/d5hMaVw7Y4S07jbWKxSFO+ERb1NSKiz8U3usLsQKySBScM+o6y
fHzc0kYAbQTOD3g+PsmnyB04QY7UgGv+sbj/N8oKZkYed3dhzHOJ0T9HcoFLGYiaPZQ/Oou2fMb7
5kVqr3yatYzF8WMAJo7oPGA/zLKm+DrqP8Elbu7KXq9VodUyfdbWnPSCmDiOhV6fhlSdGJSBEH8/
ai+T8rQ4h5rFGQJi71Uda8QVw1dfMBHvTReVTVW88lYiBI0djLnvVMBo9X8l7+Khv2JJbwmU2/5j
YF6cvcLuGFZLHX8l3D2z0alCZop0V0GDifhEplwNBMBMTTVAiTa5nJdLtsJQvYMnv/2vpglHPajr
otVc4FA7J2g7SnfFmXIkpcbU/RdrncWUxXM2ci9XqZfbOy4jQtE8Sn8un72mdfJ5QcNg7a8XYPc1
bmmxxbNu/lIlYNi4KXzh6ZUP0HPS0S976HbvXq2ubI85/IB1KUFpWIkzzaY8p320Ak3+lV82ShtR
zoQPjdKc4tnFM8/I1amuIKWf5hAIHKbpTKVsM9HZ/YjZKzOAfa9fBY/t7bw9EM/au/S8QvK7ANOS
II0EIar/D7tMbiAQyms2tgPwav/UnrCbnAfhwp71ZwuGFkbUnNW7AX84FokLcPPdX9gCOXKrvgLe
W7GyiXFTJ5qMmKGQ5hVe8/sEDICs1E4ypArcw9e9DftF8sTc1j5Kpi+TvCK6jkp0SeNDFNAW+Azs
/czNsJET54KQZxneDAW6rcIi/TkAlGPLngTo+pjriSX3DwpJptHuNJzjXp8nTRg8EmgTdTqrFG1E
7cK2sCbvmxOA8CFcAfRCvkrkEqFNbh+T3uPP+eY14EmD8WGGRli5ZxCfMfglb+GZ8e89c7xPnKGY
6pQQwQOBR6pRemXK9CyJPfYBz3/J7xuSsbFYTTs4cWRM1tn/KDMUFmycB6OAsSG2EYdUe3fWxTNG
SWAPTV7nSPgnKuH0S4v3mZG+SqDBByTV/HtNNkXi28wmx5XDpGxBEEyANsLlp46ScuKp12DFNwUv
W7jZ0ApT76XdIOHDD+paSFi6k4uxZQ0LmlhF0PxObyLfBw56cAi/B13or0JpMIho7HA6z+Bjm0NQ
+QFFtbbyNKwpK65k+liFWLc9JY9kGdyFe8y30d7jIyyeG4E/Lf6nuGxGDld2pY5PNOjT2yQhBySd
5uqPelrVfonISkl13Ak/stQzDypb39ubWwDOgvHVH1qu1bR6Ny4e5YgYDNmA3YH/kRvz6pZ19bJ8
iXRTe5uyR6WI1us84EfSOLc1IvyszaBmY8ZvT9JIddbfDV6QQPm8b4xYzIfXT+C9cuOY38KzVmJ0
bzjk5tsTYrE/Jlf+u0SlFiS5CWZU9KQiEDFGZ0ZRZXfbXsAzvoPNmazIHPbRK+YrONKkzhFJwXCp
TipZrvG17z5/ZrTV99IvM8PrhFfZnSQUUI2PCR8SjJzEDxSJU6fNdEwklehLwx+XsOPI0j8SuiLl
ihAVtqYWMUtBIar7YGE0cBXpyFahRU101kYFMOFzgbNZ/WtvE1zNv+kUgPZ5vPNQrvjVdxv4NCId
7YpAbzwdNfh2YTvGaEpDFNX5uTPyqVz3WEP2duRB/kN3PtdGHOGv0g9Pt5d0ret/RIv/PAVXIGO5
b94mq4h+Llwlv/pQc9tWLM79KybMm82n589+/Yim41173B0yAnho+RAqYhlVpef40LVJCEUv3djX
ZkF60UW5MOmBtCXpU76/mqQSC9ohuIDXClCTNIc22NBCYS8kAV+4r/A8iyVAGOusOjD8qsP7MaTj
KePHd9kRDxYVkH//7H9ADvhW6reiicUf+iFubaOG9l1+KY3fVvqDKvToUOlWVxoYWx2V9A27PXMs
Py+s5FcyIYMtRKhVPethDFYS6xC0XQGERCbVRtQ4K5WOc6DCC8ucoit/4Rq9LxYtodvmdJm/uSp9
WEOHBhrM/1n+RwCeD5bMyQmA3+h7yJtfgVVAMSqoNlPIAJk7zK3xWfRyx/ea9gFqlL9tFVG3F2x+
jTg8HCVmYXZVG3v/eF7itXovTquYxiMkwet7Pv42W++5codNL7vb2Zghf8ctrG4kNqSlIroPoQaf
Ivw74B/ue06WV2mU89w8BmDJtSqIlhpBE0nnBhMnkwO860Kx0FyNi684ZJjMzG1UUEFyV5WXGzWI
tdczUe/Kj0othQkt5kZ+dflrgSRHKinjmg90jq2APZ/4L2yg59lUuwRddT9xuVz7Hpibn+HH960R
74grDUtgOJ63z+i8XjREo4FgWVdxecleL1ZorFgLY0xKj94G6hJi6z2Djk3RrMITFrfF9H/p01m7
7pDROvrarxhxQlqyN3jPQLSt+UsAkK40Rh8o5XZPAjDDPN6UchwGogC1ExjvXMFUnn8JW/4U/drz
ODUnpcSIPSAJIwLcwS58VLKXB4iA1Qm3SsXf/IJuQKhUEIctDlbAulZ90rcF14/7MTkE1Uw+jdnY
K0oHyLFNn3FooNQSWQiStimppJEK67gkDV7P70a7pf6qQSPyNGTNC5W8pbxxv7LTNzhfILEyCDXy
KtSVR4MmmlF8XtP1R6xsC5UApXD0mdIu9tKn4fDQEESWH1SNnWsThgFHZSmZX50zQhIq6R3Auqcr
S+xWBPRRksBXTzu9Cl577zm20FssIqd4jcqMbP9EJ/leqNW4F4MeOyxlx8wvFbEyF/F96vGIeuaX
kulwLPq7XaYsm++mNXJdscQc2OYAgdwiMIkn0foMcFKwi+Ejyq+CJKmHvY6HHAUdJkLP8MToa1xc
Z5nPVlxs8IBioI9TN2amZ/q04jp/weu0S2fU+ww/ldnDj7KJKJ6OIksGv4jPEQyZ53Kn1iYfRdID
fTl2IxhCkLFP8f0d1e7QJQriz/xFTfOZRDaQwiUnWhgAtz+TI90G64Yosoh8n+jsBvqzIW/v/VJI
cUFYzZiqfAD9QbO7QS8t+eXJWxrEVahrtv5OrFAWAXG8BzbAlXrbIpGqjKZavKwxTmWNhGTTzmGG
lHPp9y3/dH391U8i2791wOTKs1mGfmloEHSu5J3FKXTkBBdENVq/nf0enbH7JKoZlNFum8vrSvnD
MC819i6DTC2cihZNx0LKPpEV+WUtZtcxcGfBRFGuBAslc5le7861OTY/8LzlA22S1agLSgOKqnMx
FGGmTT27hc/l3Xl5l+bjSyxb3SOCwgYyHS3xBLqOkYUfEnnjopTcZxNtq7vulcfsCIuMuf+hHDZz
L7YqBwyAYjvgexfrhz41C6Iy54w6PEVDym5udZZOjz3rEwCm7U16OyaiGe9l7nXRa/L2udbAj34V
652o88w2Ctftff9MWNDNSdy/9KR7PSi9Bz3UwLG+ZjMnkqBO6XcB2RISraBBp6skxK8GnuFPFgPX
T6xCk8H48xHneMIPpzyhm4PbRAeaq4zhlq99Jin3530TOHq9Qro7GSjKfnToNwCZW0sKET3IaF+o
THxTwNQAPtrSRrj0Nnzzr6pKmUeAMEbkcbLaCh8dh6KlVld7gZ7rnADb2Aq9iOF7upkicAMyL7XK
mzF28BMjjFHZ5WCGEQjswpkPItS0rGxelUrASYQluClPUMvqkVdgcz+HpA4YGTO+pmuA050KvJug
23ZTMK3wH2JPsopDpFjWER/ZgM0+J2hA5XFhp0huAsxMzjEznR/IXGOkCGfGVyOOuQzIepmSip44
ff6aJS8945tQ8dV+sVf1N5az/K/IDYQT/2GGH4MYXh5eEwTdKqggzs07viaRMjbsZ4WWnpeMXO7F
2QUVoaVqt5dW00bi5gL+46rhd3U+3OVnIvt+bCfB3wuqKFpE70BwzECa3Qa7GORLk9RQZ8TG5okG
3OIGCYBM653Q7HGTlUwQbPta5WWznP37+UM68dRIlUnu3Gbwo5FoYHgBLQ8qQGWbWELCs6xmENHs
yH+ydx3QOTnduuIJYKyEnPmrVL2LW7ALDqlQv1cBrOxAEWLp3LO0IJGkOJ9tB7DFRB5Z5Dt7tjSj
p4um+6oyJE6kuUJaOQT9pyYY0ADrQoZzvh89cL9Pa2E3WWLv4hycUkteayj/mRBpoCu8ymmgE9U/
0is2lz+OONW93piWs8t3QKvDqWemERnc8ivqdJp/fWNjmY9Aq056L2ZOy8Slv2iEF8KCfI+EAaoG
GJGV203SPNgWOnjFpT/1rPbdIKG+giYE2z/p0Z+pQYEBoqSgSgrO7l+goO+en0mc8Mxz1CLrz7cz
sdXyca7nkC6HxD3CXADndeJMIyl9FoQJ4G4rRzvb59q2G9hFIdRVKaRe5y984vnOPPo14l2d80ef
wUJ2C92apajUvAkVJEegnGmJZRRLCz/KSKxWKm3Wz4WHpXltW1EIxihBM62oSjHAzSjyZ24q00DB
amZhIQL9vLaiG6YoVa78leGHDx7d6siodFsiLtvM9WMSf4N5aj+KXxFi1guQuqjIm8lW3xsbApma
hDIX5JlFgslZeibpbyTNVH3G01mvUl9a0rNTlqg8GVTvf8crwcg4P5scuLCM0o/lQzrNr1gh2fHH
12jizjYSBrc88o8bMsH7nmBGgumAKWa/kp/9Xu3MjETec7LqNUOJ/46WpMXW7UR601cQgepAA06M
mDqzASJCL28yTHeAUSBhnIIdxfsdctjiDIjN3IY3a+6OjJ67ADW4Lp5PkU/ZlaZskEawW0wBxX8m
akj3VKzU0eTKwrFr6tbK8iSmN8sdu+j43kgyjlu9dD7qXAM8DDUcmbSTHjshNTkNAbARCbb7wehz
BA6isBnxNI1TmbfYbRbcs9whNcbo43hv4a/ZxyY7etOSCvleFe23HCuegnERJC/W+uOd1FEBKoOZ
Nj/YUWQlc/KW2RhaSNqy37Uxc3RfEcGkBJg7b2iGuy3H4E9LeLEtGa/131cY9+fVJ9rh8vQvW1w5
rjPqgJ6yxEJ+rX/8ILhA6nOoofw3K5m0oGa0MrD0melgcVg7jDzXCoxYcBEnPVFw4LNKFsfYmdZg
lyf+p6XCg6cyzNzQ8PEulgDpkSkfJCnBb49DFXHBnuycKpGmpvhPJBSgAZzRhMp8ziUajY5f3gYL
9ffVDA6FPrQrj3mYwEo4bu2kovnP2uo1IhuZUcQik0HU2RwVOBvgDVqXJb3FE1aeKhLjT9BwCTgK
iG1pKFxP8uLXnI6TKbiGbpLjDjSWjP6futH08Ot3T+aV1O+rJj1IjXuI5zK8YB/9ri+PrfU5WDfR
8EMkw87q3SonwQkm+5PItXSTkR6Dzyl5uB/J8Jgxv1TZ5CzSBU4WbkyVaXEf/v0fh0GS+/wpQWej
kxQdVs2ug1ctVTdlDYRv9ouxeIO15Brg3NbAJDHM/D1flELP1Kim4oH7SjZ88yDMaiky8fIEYj8V
9GeLZJuomYF/A/51/MJboNd9ndHcpJfm1To2C61tgx27wUUIt5NEZY+T/qQDArZi27pF1tB7s90y
1LLsqfbK31XaopT758ljkaoOuCYgoOZ5F8GfvVqW9cuPC6XuromDByAd7Xdj8WT58OoVx5SxL98R
UR5kPAWQyNtAX30iVx0o5Ohwf+NRGyHNlm8dySfLQ1GqtCDYFX74D5BQ0ju1FHgaH55g5eXH9xZM
LPiHLcXXUSVT0xrIReUkgoO6CPAScZXWxlA+wPjauFXHwK7z0QiQjMmgst2WlwTTJZvd7BXSyjQt
mAQ1PWJM8o+nrYDl3Ul9g9cK/soTqBaQ7wOUmXQtKCnhHrNrE7hODexpx7tGgPchfcP13fHMkrQt
zg+adyJuhNE1n63EYUc4s9cvZgQmvcP24eLTCWqAeJA3XQ2kaF00FLeueCDNuDi5f40taGZ8VUwl
4OVD9oUtMc6d79chYSGqbW2bqxOnc4aa5P4MjgCzuWT8yMwXX4+mathM4uf/ywnVokSKkHPs0/eu
rkBpIyf82VnUvflDPBuoskgOlg5jhHUGBCw3bHYgY826FB1Vnrx/tBUqxaLIkC8Nhm4FrPB19AZC
CVWGFZ35IG0p8tadw69kAmW6j5w9vWbX5lyxX0n3sOh+t6eWOpuXOCUyCGpjeR1IwTu8QkYYHB94
GSFsSzNoRAmDRgteMNvMZLManBCfTETjsoN6ny7Y8qsFs9JLA35a4D1bkMBh09jILuEW4GVZXf59
CeufFUbmRcY+Sblr1lXMLeVAQq+xzgmCgk2tv4jV25h9LIywbMiTr9aCjO3MReMBHJq06mk99MNp
5Gkj9sQueOQua0eL/9mnnO3y1ZeF+YKvhNCXz8oHiO6HaTc/QwZ7Gfosq8iM6nkfOtIHb2ZlfpNf
I/EZHJaOsuv3nRo82+br/OUfUwrOve/2+rfrBAGaWInz1czsVQb6Dt5WDlAV5wdcQHOdoLVggzX8
staGPfZOSpc/4ZemCnCpb8dFr8PH8dZQ/ujc4gOun8WO0IVaOOgyPi8iHqnYGasOITqBm9r9hbqN
Ezg/i4el2RV/OGqc8ZcQNjSFnEFdMl2hq60D9zhqujl1fRgbIo8sp0thdiJp3LFSC9h4dzIopR8m
iUidpIIte0ec1WRDEB1zYibCnPQCWUT3BJf3+bFnQww7yu7pyGDp2YZtm4yavoGUNK3h9iyJ0X+C
gvZg0trJnguNPxTvFTbh5Du6g3orFqkGHzYClnEaEiyFiJSEIM3z3Sco1fH8d+zzQvnDKOkOBQd/
/3pV+2VO0UW/Qv+wmHjQ4YUUvIhglEc/dov91ENxxk1jw4SaOv7x7i6ZNx9udoQp/UUidICcUm5w
GliW8/aqQS85vQTrW1DoPxM4InMXjqFmU3gtZlbiVK5Dwt2Kdu0ZX62rou0XJqNk7d+GHJip/bXX
xOBT1rLwBh4mQpUbwBZspVh0rrP0ONOxwiAUhJUIertbfKdFnGXDJBAKfNBNljVzefSeujaNZBVL
7A770ofyyjiRbYrSnGDEkeEqEr86clE8r4xB32ExgFKsoaPWSn6MfDMDyba90wo8HxNl/J6QRt2L
VS4KG0OOSu3W6VCMjTHQbcUnTcwuQ9ea8pF7tFAGbXPhgxXppQj1panepUwiqzWaiQBLzrJzAsLb
io+1tgLLVdIv2NC48T9wCzoiUMGV5s9oQAMUNDaca413Xqoy2/3wojN2D8gt5Ep935xEyu2bsPo2
fPe1oinJzY5KsYAeWPHIEd0K6JeoqkG1hJrVuZPNSKFYZv4yEKz1qZImvKVgjk5C/seuUf5iIhhM
fozgj489XTlQKEaNknH72md/EKvR47MXi/zxOpA0K6Se14BDNC/1++zFnAjtB5rpwCQ8cRtxmJER
S6pP2hMeEitUGT41qO5CRuJao41PBZ4q+1vQOm5z/eotZ7FuJRAsma2DY7WnoEdTwp3T8q/3Xym5
T7KfUyqhh5eE6//ovz2+SMkBkhubkHl4JsmmwuXYf5qgvNeGEXKDUYIta24qylAGeMxYZdgQEqgz
7f2nxK2UeUZLSrPIBiK7DxnhQ267r/s8XldedSQjsisL6y3QDRSOrfXcrYZqfDaSjeST88t7uYwl
LLHu+V/wdKZ+unndpBgeuOHPbG7di9vLRQ5BLd0QWQIJ8jNUT0qdbHTysENZ+ZfE/ugVkRVIq7zd
usNzkpU2OtCnzxHjeRMYXTdxy2XrEfhwUZOPBuI/a0kQHJ6XbbbF/YbYg2DxmEIW86nYBvX3hkWt
D254UDuO5MaRYvKMulczc2aZJSSOleJkFh8A8LETPT9/UDqloQU/U3/HfKfSYfu/i6O7Bpy0zohx
rVJBkEnPHoIPB9cUvPu/UlAH7juye40DvLSl5vYSBMSfTe9GXjnbKEfsTavBpSP+gVwk7DBhJPgS
ksUb2SKLlj/6yq5jkg1yGDGTCuh82o2UAmPZmyr9BD96Yh3a4oJFNU3Mk/b15Sgkhihkb32s42Uh
YGCbdmtMTvl/jiBA6lb9TPw0sT31GJMpzdtD5yiAFEkLR763wZLv7bRBjdspMwWfRfYlJIuxv6Ms
xq2l4VrM0jPrvI0z0z/pEniSXH54B614L1qK5n31hBDHCtFkp4d/akJqaDsUx0pXwHycHt7iLUeG
zAntgLFZ9N3eSVdTyOIPs0i8ByCncwUEgiWWqSiNFMAVtW5RmFmOek9qGrk5Enjq88fMi+QGqLOr
MVNJiRfBZdBbDxudKYkPAiKnZFx0W+A7C26/bxuh3iEwQ8jdcmCCaC3lyvhlUZPl6kNUoqnX7SRv
4/oDRPfCnodHAxk0Z6EZLhEQz5OBJoH2yBhg81XeQCgL4lG8Kn6H5aqA2UghNqsKr6uCynVtYlta
PkW9K05eHInjnAG46SASvgNodJV8NpCLW5WeDPQGedt9vurAV4BkjOwGJNE6gweoMiZ3Im1nBViG
NGPwbP9r2EcLRSE6KgDcso9kVDa9HXzuXk4PFzLbhxiUUOywQQ+Alko0gQm98O0wgeIUwjC3ANv7
ddT6T36LhNmshwv7GVzynu6KYRLWcoWO9qAtF1/UoZ+Un9v+3355TDRouaiS9vwV3dMZS1hYxhaP
afdT62reqKHLS81+t4ahu5uaZp3JeEkKMQMRrR1IqmROkrqbv5AqZX/rjnM8JLus44UIit0jHlwE
j8vw1detO0mjeMdfFnZDGA99T9eBLG65QQeLz3Bd68xfoK/gcNG9g7cf7Jw/dHmPauFumChTieAj
i4WXkfjPKxBcyZpDeUAi2SVSaOcxM31l9ml8pD20PAimxYDrsivmWueadsL0sU6sN/IwSoyuDAno
gPFKS7ZYNxN0KUXBWjs45GxXy9g7TiAJfW4IfCSOLH8Y7sxSk9W5jLhFokwHPT74wsaqBXsZ7oRW
PHGfnm5ucjtHL/FOtQfdIIoSbntRhlB1wH+i1x77CW5yhzJtxWkDazXYfpc7B4F6uyxMZhGv45j/
W48gU6BRrG6zTH/IhXxASQ9xqLoWsPJAi0dIq3htz3zFaLEgvXvevo5XNWcIbhXjj6n8olhWv90c
bMn7xysN9EDaJ5diZTokerobE2+SUB6C8rOm189fS5PkQU6QtDfjr6/7y89AHYnCCmW69o/1A1g/
lUL+xTraUh2rJbWD9eW4HzJT/ybzw/6CmyhuWCyDiKqxU4Tedynw314S4YZDH9PwtKpBmqn8PXWU
3PeKmROf7ddBfQof5ha3bqtxgxTbSZfVZ+4fklALMXpIWb6Cw/NVoD1L/mbrfSfpSAJ5hc5oiwUt
HgjPHTRbrWXYHWp/otzC82VwcBTp/T2ToaRkEDsJaxvrv6pKqVwfTz0H0TimhEm5M0PKnpJFalI3
nzVPn66JfltO1S9NfA57rlXeY2D8WSRkRA91tKY/Il7jMl5hkAQWAerhIuaIKbhmXyAm5vopflhn
2aytNberGbjTH/wjlBxG31DNTC+6ThVW8uzECJHVPsVEr6Cs2j2w+6nq3JZEmFsYu5UC5ztsCmXU
fPoDd2yqVeCQagdMh3+/RY6sdJqtf4jIkLcRc58iJXq5EotFwSxqGhzukcZX7Nzvp3UNuopAlz8e
qfu+EE+CDcq0Djw+mA7M5khhEsUQjacKn6CVLZG8bRv4roCuk6ezQWMHua9rfEXm6d9CGyjxncYo
eN9TLQe/stXHmaWXEpHUcv39afZEjq9ad/RM0qDaUMJtn3XcYiymYr8xeIrwwN6nPFRU5SuQbryO
q6pFkSIMlgvseGsfDLqp15QKLjHVagxCl/XA7qO5aV+hLRWObqNWexZsUjjgzflTLJ6VV7kRI8/E
uiCElPmXkGwZVpQPJyzfEkh3k/JHhdw9BI7KEPagA7BzbL9p27AwglrvV3vh/uvaMCM1zLkldNfD
9GBFRqU4eNUDdYZ0htNaUoX2D2AWUG8Ta510mLbGDL6t8qB5HGxt9gFqdCQ7apc6kH7t/Bs4z1OG
Rp+UCO/32BzG+tTn5V0+4iwVxBejRKI8Y7K3OV8b8X33WRmM/wM0q4/MOAWWEl90L2jvel2dJ1xK
66CLc7OD4a/4OuZvTrE45ZLug1yscBqjrB+uRe41EFZQ1uSgmYA38MndNvHlk6fMJQuwhN5t8XKF
JCNUS7H3If8mO6xDJDth4SEu9+Z19w9uLcOfTTFIcFJwGkLM/+edE1crothrh8kz6eBZ6cq49c+A
rrcq9EKw1xPXAKY1BGWKWDBjy/BUtHxV1zNU7UIgL5k/WCyXA19ANRWbdtu23QXobYdbaDqiyJFy
8w7j2Tqy27S7SSUqImQbMMEOG0BG3gVk4GJAhLoK2tvhU9sM1tei1l/DbGwKsKxtRammIsoHwxZL
0bVIffO3uDu7xC2oktwIqbbvAoaOY4/X1pmoc7OvrNVE0hTaQEtBClBELUrqdIuLFlDuZNOIqTm5
jOlso1sXSvhPFEe/8sfOuIkdOkU2cKBHrr8o07LFVQNh/I5hS+VZpLeMJveSqCVnt+QixsPHglz6
0oFcY6TjMJ4y3EHK44ZDC1L1pHNZZu4/Ion179n0pGuREeh6Tfoh6t7f8RnY/M5rrtUcIG73gNbS
tQdhRyE4hO2oHfnsKdrxf80AXYy0Grc9FBj0jtPssH5SidfUIeHzwnOzk/EX9pkqN5Dq/LcfK/4L
Nv/qSF9AX3UXDLa0e8itJ1dIWunRUTVGe0kpYfMvUT6vwRBXyexWNZSX0vCwure7VotI5zVqE08F
MJBEvisbrxv1DEo8+9jcggZqeYi7gHY6HpFi/DQpMk6XPeKIVCgCK0wqIh4ZQca+9MyitaW6EoPB
vxnyY/1n2/8l1HwGpJyikv2woAb7YjiWPoxucvMCZVDA6OZxdDyomOsNJ9DWPYq3NKh2RtTdppOn
Ro2UngNwCg3Y56HNPLXVKt16zYSWR7AZQndB09M5xKEKIhv4qFOqAC1u1ovZ37WJka836LZusc8x
xfN+S3hfjvZMhVopfndHC5AV0+bHq9yGz2MJqKkarVk15F613N+bmndmSnJhu51ppENDPql6KaeV
5UaKbBePWh7gRVnYU1PEG9cKMMIh5se/3Ub3nstlBX6vmk5rx0y6jcedOjQOYEUgZweK+VrWH9Y8
ZGDzy2NR4M+LZ5XVt4AWoabS75jKFAfUl63fhB5xi9j02geczs0ib6Wi0B/baLPxvbynaU01en/z
1K+Cthj+obX8mwBUNm3t1+o42mzEVpF3tCZVh4fPq1GQ42uo6qtVlMvP7SkKr8GlwurXVWH5EAwa
IPuUXCPCAx+ywXfj3syl40n7uTW65rfjWzb/tC2TZ4P558JgXATthZ5O1PaNHqpeVOeWNosWJihf
wrxpWtxuSZzZsnJogwWePMnM59RLWNpUGxjS6K2j0eC8hp17VI/4pdhKzEfD4dRzpaAQRbGfqK3Y
oov7Jm3+uc53PvQvueTnZigjJohXufek3nnsvjwPksVEVODIbXGNPx9VZRLB99JLuR039yCriY1N
n0xyS0VkmF28Pe4sf1hzOhM8Oy29Vp5yJbvMFfthPr9sPwF76Zoh1FYfYgts0JRZdOi4J2g2EBfm
qUW7JIvRKjxkbGVBAlwqjw8QbMe46Caw6LGKpPJal7VVgXrtFLH+6IEYGznIXhE6G9b5FTSpbLfd
j9vGD3KSEp9oh0AyRqpcts60ZM5l4zZnOIdiZd8Ii4yjE3v7aCO242rBLiLkkgGANhktsU+0P+AP
8XRJW2r+gIOsQZbdXIpPwdJZ/+WhfLGp7iQW7cLFgk59MsXIc5oECOsiqYVo/R7CbcYyMy3+Clr1
D+/Vue79QuAhw9Smq9cC2gJIaM45LSbs0ZHmgMr2DNhTq79JHokwDTIp7SLegg4qZMY5Yy+ZSQMY
lusV9R5L37mWzoDb3oaeYmN4f04dmTLOjKpSkSzB8M/1BjEes+XfsoJbYKPq9/ZZdnGwtAyh8vjp
u7cOk9tNU4Pu634Rd5C4JiH2HW2YPYUgfDvu8eJOqamkZr9SSXo6uyekmPJR4RO3YtsJyS0P030a
KD8OZnYCSxokKhPC58KdhDzNLiI9uEkSUHhZxcxfuqud3EP9/+4PXbEVICWJVNpx5oG6a03kfGhA
KCPmvTW/OpPcqO9jx10HH5sosWjSl8V6I2HvRDaCqPHHLWpS7n8R44545XI6vTy1LAx7dgvgVNLu
mmVMRYGxIqY31W6lkqiNBFXpDqdc/83tMykD+g9xE039xtBDwCeq7AiI9r4q2d9LkF/nFBtPeb1N
19pzal/0iXBvmg0wzx0CQhdRiHlkGnHb/py3l9pFBsmgYhK5DrzLX8PmiHxpLSoKnDxW6BDILMN+
Rte77TavxXnjSnNyJTNCL/j5DtTEbt6IVLBPVTQHe9LVwmNDYeqo5uw+QwrXnppiNO2pW8VON7Ec
xLxw6IK30I9EZonEl61iu4bZb+7qja8QhjyT5JOe/33hM1LkGakbXdKKt7xPynk1a9YsDXck9JLO
tVURwxdHtkZTKsNRn+QD5iFYI/LLP/IPCr7dhsEFOsNh+rBsTIDtJ2KHNVKvcOC/bB9cXYQa28Zh
cBdCN5gVIJxCkVP0Fvm5P28NgIc/6NQewME1ogGLfaXxoIIsaaYnG2LFvb4hTQQT2Ckq7wOZyGwE
UnYGFUzDrIdPeYWvBkDnLxLYSlgjHrXmm+FjkqA8lhfNDp/VjP3X2CxBuTbJ87xEsR7dAvVb6eLL
4wNRoVBa4pvJTVqAdbx9yNj3Ime+MsI9mt1I5ZHKSo/KeZN0lELWY96kyg6WElvWlWxv7qREc8uE
ui8NhgNzr4TsvvqDdAVQYHjb52hV/ASiXrdq8HVUA0pLp2GYXtrve9x6wFfRkfDtAihHAhdHnq2j
KazloplrdNkPytZ6DyeEVuUWOiLdaY0wxBht4OP5dw9D2r+frXQ/vEO7wrWnyY2l1B21gHBY4upj
FpfUhRkWwe2MbeX5POTxPUM0TSaaEIIGqsx+HIsn6wRCMAz/x6MIhDlrMqWRlljCBU6ymKnfsRWD
E7q93sWfJuAGp6ZNE0IUY5lxniUyFickGTLg5Lnh9HiLI2pvshC/mIKNAZiIQrR7f3ZcbOusDLuH
vU0U73Fo2y9TIvgv3lDNTtuuu8zx+9GVdzYWVCO/5R5ZCpwI6nnovQv96QcWEBGObQrkOca2d3zf
Zb16Tuu8GWNeradYG1cNJSGxGffgtB2gK0F+tCgyWgjTYuxgEScH7l2eW7jthTNfdOdk6Zt0XkxV
tIEbPBt6Meb7SLsohWLXOoY5FEhTWwj0W8Uk4YOBjoJ9dhzQJ3tc8Wftht84doaCnzcG2zS7HU/7
vktiI4kUjuxEORPPF8k/D4LuXAslkQmNrBaSTSG8lUUpnjEOpVkteylZj5XWSaYhcOXTZtbhUd4U
uiVB+apJPI54sMvbpq3hql7u7pk4v7g5gOjWBw5eLiegGteZ9iiFpWdirZg/8m+weCylX+NnubMW
iaPaIvn5K6NMGbJVendvOtmx9OjTwQiubTcRtpmqFy0GFr/nKBhrXHCHz0X2tmCIfXTTu50JBSuJ
aEg5w9RMVwRcrjkI+Nmyraxjw9OMGWP18vJgAcVvqYpsKu4Z9fOBq3rWBswR9yBJV4Yy3ciL7CHb
IdOwyDGmgs//qeXHMuvdgPENXw+pAIlAqEL4prYY3oSgViEBJoUejHW91dxietQFQ5jo015B0RY9
uiMRLJwnHX+1RhqGVrWsLOWvWQtentzDnQ2N484jHfEuzkZvgntDpEi9xXPDB1ir9U4ygWfG9PZq
s54aEAn2lypeH31IeVU0E7mrZuzXK2Ke+haHmNkakdo41tYT8lcSSPwFYcEkHdpotABgXiFoSaAu
wRA2RxkuZXn2rBpKEN1yQbsr8H2xmlnNu+X2auL06Jl6NcWapQVQdxSCQ99QFRX0eCoiD+tD9Pjj
x6xmuUX8anITJkwUasplPwjR4euLVYtQd5qEDn1F2RLVESUp+MtIAVM4eQSeDHW/eQQExQ+WGlTI
sAsahUHQQHEfvXcE7c2ehVv1wyyPB8zNH86TW93CJOa9RBM/blgCo3hQO4ya8K0VZm5vGvQL7gdV
RZAkWnFXcJj6lrtVgrAZ8udUgu65CiBdqq8C2G479hJGZxYP95mYpOtpuvJff9ZrEAQNo92jLEcu
iAMut1K1XsNM4DPxiVjGE3RgnWDk2kiFS2kRhhAW1LBvg6iYz7B9YYDTGEkGJpmcm/M4+Fa7KHsV
ckzvFiuKrp2Xw9e0jnuhipbwf80i/9y1GaeLAH61m/J1vJbVnhjK3BNRbUKIFQartQfVdkb5vGVf
HrREFOqKoIETS91n2UV8sgZNEy6/AoU32wq15r+MhrP1a7p5amwweelfO97mnMCG7F+0UzOCEdtd
QSC2Wvkxjnb878KRwzaeDzrLXD4HkPAB42ED1hEssXMGJfgaO0DhbrLKN02+b87tuBOWR+7wWkhG
CL/xot2Px/lJG2KLyxSRzErwN/gBj6+hhAf9e7037tN7PSGkLO7CqWKxrHU4yhcJ+/RS99ZPAPNn
W8iPdOdjGeZt9WVqjqbx6Wea2NzbqEgqrHO3teLwlMEMZirilJpEGfv7cIgx4gQRORt40oj22Q5y
+Pwj7tMGiC1+dQPXgazvsddzbJrXkrIcNIsOgIx//TBbTHpaU6EJEMlSxvjtWXRO84VvIq1k18le
8aOSdOtD3MzjEqf2OQk4oMrzPrj5n2q37Hrs+0UonkPlElUIrYis5rHkMQcyxMiXXRdhL6146IJj
By2olWlPeAre+F1LLMTDhMn7OYOEqD/Z72quxBgaeA09eB8OnVvm78VPbU3qfpL2x1UA1BP6AE+X
41NwwLZRs683vZOfCNB5SZzdx8LmkeyDRTQ2K2BLrPWS9wk0ha6RBI/Q800UXKQLmWVm9UEodesB
6PljVs/b4tnYC70RrTWf5et1ZTUdOBBadq/KDWS/P0F6S0I/Sgtsvj8OXU5rVAeCutjGWycPFJ9w
P2pm8VwGjdRd/6v4f7n8m/7zk7jY8x3udWLRnFp6k68UKTfMLQHGcjRK432wrRqHjZyADGeWe0IV
d1i+FWSQ/oQyMGV1BnMqxdydsSXV3CbI28FTMwqV7QqZWYgG+D8fBOscxLYquwoLzQzKShLamQrd
Z65JoM1uNT5bIkwsmpsY7YTxF36jjy9zPWkogw1ZR3ikAL1kmfNvRjQkFjwbqwRF6seDiNihJzs2
78OZU6wdfzXZJmUavmnqNBExyHTmP6f0jFzmZr4fWxdOvSIe2leg1b3BddCxb+ai4jk5A3sFMpp+
rsMe99Os3nGR/LLS2C2xcSY2rREanGxI7UOITJYIoELzAOpZKzsln2tsG1yRgN/EPobgrva+bSIE
Xor4jKRyHEz2NMM3Zxa7fmE1gBbSOPKpbfGRJLab6HSgGQ3pg0ZoodytB1YK9FnS3H/o8VPO+23T
rj3TOoirN+kJXdUJW9AoiATa//67nQy2JR1ItN9pdPTzVhZMnBX3XbjqDYJFrLDOJ3BkP9coufzY
sLpt/70SFFX9RsN4b1eFdRF7qhRd+6U4T2BGPqYbG9IT3XKNZoDR57V5Z+i/f3K70YWs76Lv9X1G
Vk5wcRzDqVnAKMmzYO3xRsTw7CdznkWtt5Hj+VA2WKM9HtYtLGb7YCoJzldI9WmhyydyacXwfm5A
QBVtGn/60InwoHZnutfqQo6b4DNpgLhV9I+87+Z6jRx39Y7a1AMbfQC7DJtljKn6LkjvT5PtgCVK
XESNwx+bxXYpje1i7ZFYeALweSXoXoP4WsubHj7/3DvHopozA1sSuXMjdyI+oVtvcXzhruJyGOry
7J5W1IPeEH9rJzxMdbCjenZ78vma+KzRO4luhicZ6QLTY4ngdmy/kCwGKoVfyc5mlG8+X3ipYnLC
er3moLqyZT6DDhHLT0YEdAe3CVtCTdUf+JViCdpwC+witfa8n0HYRWNkUheosg3thmVOuvK8HJ20
D+xVDPjmV+5niWxI30i0leZ/JiXylns8mf+zhg5SPpwQpJR000vPxMb0grtg3rgNYDPVDrKVuV6F
W2u9dlg9PD+FMxonK/foGJ67yX63Otfgqtx+Aaef1Ax4tZv5K5M5WlwtWumgs4j1iCMaFvXaEuVl
geQWTQc7bgR9veAkpTFz/HFMv+drfu288DpMBWzkoJeOGvji55pVQ5ZeSAOf6b+M0jKttbVxLCU8
BTAD1L2AwizVNkPd7euV8pdFaKWQ6PwbAOVvFD2pZKcGojZFSZB3oL8BhvvXOWowVZtj+w1YCi2p
r+YTkbxraFAkgNIN4FWcntTOJi3txbT1osTL6KjwwmWrbVi0P17mP6kjyQNRP66wDW6ev5eLChvG
r578EBVUxYy0qqAJJ6QxiFNmUys5/1TWGM8VIAOgzc5poJJqVDsp+/JVo42HrDQQuzg89nswzpNW
1lul1F+/fOjZc0vDtv/yk/tZ53J+MD2t2FFXm5Z1qDonneBXPLUZNsXEDQzY8K97OeszA3JsJmih
D81M5Yw97xy63HDGmyFQ3o6rM14UJIGFF0H/N0UFHVH4h+NqPCFdK8AhBvklBGdwtysiMA2f03iL
lel5fCtcQRHRsOmkVSWKvyya7KAUh6WcFMj9Hf6iLT+KbeTaC8tquxtej2X5AcgZFsp+YabO4k7q
thCIp4bdyBqWDM/wsCi2T4bCr63Z+b+tCx/HIlnZLrC14Ycg/rxDHbvBMZ+i2Xx/XXEWqvW1Lyj4
6xgrLKHH33OEIx/ZwS29pPwoeQUoWTzlcbONl2P6WZ7oFENTMS6T8yM/vtTGUyWIUBwyB+Zo/IhM
DeGwodUTOTg0LG24CNMiCs5qtB8rFjtX1YjS+SfjxvOz2faoXkZdLQUsVdlNdEBCPe2V3Q76jBz6
4p5rjF5iURIUPKFkSpN36GFAJIi7ozfr/wRChCbGUf/nEnT7O+jsV5ZI59RuPIxez9r1PEI7Ldds
gWrOpKg8q215LlaWE0GNQxGlbBpPdAQ8N18OaINyGbU9i8ZguannwwFbXQGVzavWsKZVbkabb5XE
WF+Md5jsNpbRfyHvLXF26yJpPIioEYX90p6dEhjSLb2hhi3ZxYXQGRavXy9iLNXgtMHEvjYg7OJr
uS9aat68OSbA0LRkj4I3s1EboTHnGnqQ5tkF26qhqzDNjf3iWuFxM/k28FtSKISjNWdRg4h7zK9d
MDkgfHZwMEcPacwgCtsKBYe1ej2wroUYK4aDerMh/hLCCLotK7FqJA52X4ZMTtmNoz9OQKeDTMyh
z/S/gn82ehbsGmigArHZ9wUGzREsw6SjRJ5nPlwvAEuIrjNSxBFLDFGEjSA7AF00NrMb1/1nBpDd
rjMX42edivTKYcUZ0EtftHjYz4zybj2snrQ8gJFJt8+k0WobI4YF648mtG0ih4T09yF288F2dKpi
F6P/ZkX5QJ1dWBCaApJyXqWQsjAbyJ0aa5abxKjS9FeBHfwZmLqg7q8r5+OkFPLFdf7FSKyKAOdL
OW1pd0MphrplfVnAKwjCfPi9kirEKK2J3zonGSNKjPufTAgofvvfYkhxV6NhCO3JOqwP6efuL2ir
ORl/MxJrQPBQ5t8KPu8LmcI7/ipz7bTuzr/E3LfLWqgT0QDpf8nvfmuEbPOi1G7NLrhqC06/jEDD
GHMnCUdXXCVC+HjgTLvNt9aGzba6MUyrnS+hfaqVf3VaJyMvju2ljOiomaTvpB4dMB+mxPMgt/lB
+9k3e2cJbEoLTIp0reGyuNkU0AEBIJLk75BjTLLTKeKFQUzpMVGFG39aGtLnMl1erFL7Sp/Lb6gZ
BBkuuDy+xlTaje15BkvXV0Nn3itExw61YXrgJZw74a0I+xNm8UHwVT5ZeM+bxwPwZGLkizPzpCFM
O0s3xr2IQt8P8Z6OIMJil8sXHa+Ie+iKIoE3ruqWOkKxGlz/3gBTwKfeSQ21LgijF2U386FQ+RUh
AeAXRQWWXcTQDTIz3J3er4xMNIf60kzhZzPtCghlh7lLHQRM25D2O1hyIZYXAEFeljvilfUNvS4x
5CHa2GCZTvdgd1ZyBTcOMOfnmQ+bFiM6DtjMIS55ljs0POeUhPEAVU4gtvsqyioxrV5hGEmaNcMi
uvw5SaCU5ERBdhYl87uKN/ABuU5F4zzU01AiI3pprijzHn4JGV7NN5N74h0DAlDtYVDFc5Bj9m5f
fjJv+Hgsc/Jm2kinncDsO+vp+nxffKF9Sjld/8LOU5MjpnZLrN3DVNKBXG5yW7glwLKgNCqsngzX
K1b7uj57cXK6OqHK8GHlSksMZJtxwa/AkfHVadNQP4vekHJDtNFIzfeB4a8d7r7eSasLLnPiwfaZ
plwaGMr6p/RQbwUB/AxVC1HwU7kQ3xLvPmwOnc8OjzBS/ahxJFGhNiuUv1qP7z3s6pn0OeWCAyf8
ZVdUjfVA5mQqi7gDfdzp7f4xqXkwOuo8BFHsLsg0n9b2zjFfTXuIrxDPdzSkVGAayF3Jg3uGCoBt
SFlgV6ojGq6IcVCAK8uVYTk+ylx75wB0YohlBfumKuIG7QQwP7aOIo6QRZlRoHrHkCd075puZ6On
27OTcu6ABOoYXEyVgxfFDbcQW4xLRhshWwu5/A6X7faOaFv/wvGncq9t8msPo0i5+r6tlBMgg9q+
60swL8vxFcun+fuFPDTAtQLdNAbxpVkq3x6OWxs8GOGz+miNFvQdUMbaeJKzIFn3S4TTYMsANnsh
Qs2mw/GExCdZYKxOWyHo66pYrIB90njUmUzMXclSMMLAPZzADh14ytrKiye9kQ5SqzHLXlSP/31G
Cd2t6XMYGfrfOedc9T2cZ1pMZyEk15Qeujaz0AZnv3OfykZTOOLg/9JjvNHV6vBcUEm81bkeMcpZ
Lr4+DHQ7FMB9n0uAp/0f/4b2okvmfmjcA60HxBG5I5HafFuUH8WBISBWp7sMOxbkikcop4qZKvqd
bsK8Sj3ayAGLoTbKgIU6x1zpAkRs5Ht+u7b6vRVDdtMweJomP/vOgYqfKsu7/JbIrDG9jA9RrK9v
FaR3s7sukdmGDU9AjXfus6erl3t1lBQPMocIV0tJMqExFiP4BYbj+CoWaBHDqvcQ3BgzrXPc3+Zp
hvyicAKUOWXE0WjObImq+7e7F+uPjJTP4m8U0ocCv7m4jR7cJT3Ft9sPgqlbeIRyg0pX9o6XK7MI
23NiAlm4yairIr4wlCB8b4XC28LwtuJYb+JhqsJejwY9QoyMywiyU9Y+6LLaOPBhFtMzaeUZIviF
x/Q9JiN64sxg4X//RKp9+ujrRaqbfu5AknPXpep82AKdZcx8bPft6H6e9qzUJ7jktPmX5v7jJJD/
y+WrbQw9mp3pjYQ5bPbqF+9POAlMbfsaPgnex2Ohyst5/7b8OfmWRbI+pH8GhlB6l1eStl7VM0k3
h6s0yZrRdgyv1DeMfUbOpW6IqQa2YYgjLqLDuubUMZbyopz5yJn5kYRZ3pmdK4B2KmWlNx0bbTuK
F+0UJd+ztgOwRbCnrYynMks7xsb+Ludqc/gCaRKRiByahd2Gzp2jBqJ923KEoFO+ZPXwNC4NvaoI
aFrIlO/WpfwDDKHx74yAwNGgJ6jDGeptPoXGgsNpglZdIt42JuZ+jgc0JLNUawTxNq81jP23pudM
LGQljc2CFrtVr+jdKlqndPwXuc8wVYPsyRccsUjFckLpuDRGwV2FnBxoLqpe0zEegcfRK3flBVnP
Nuo0gZNogqKjabWpr0myzOP/JUUhDiWLRzn5qCs1cRqF+YElEtJEvOnLg2Btupi+uysPaHupC3Oj
8AzUBC2FErPhR+Yo9xePAIi5CMUhPRo43g00I9dBQl2C2vKTqsOorPWr2J3WUEPZb0/aiyGddSfI
fybOFSB3c3KKZq8PV4PtDyYt321kaetXVy3Z8LK3BdxO6qhbdJKrZAMJcHIs/VaUxOhtJ4/UzzdP
qt+fCb4D6j14IJ0tOjGEtXaSDDeLG/b3mNfbF345MyB6QeTAODdK7+pqbOZ3wF5uTntgjLRrY86N
BWWLogYa0xnmZ6MCZvhe4wlMth+3Lkc50GdKBLa4ijP5/zicEjPBLp7tRRnGheyRjBlK08Af5Daz
/ZIBWCtNL+KKTTWgn7S7RA5k2T3QCb4ouXY8c+NLy6Zb/g/2ES7TvC+vyRiiHprlZf964tbf4BwC
BLTiU3xLjByWeQkL/e+v9qq+0rGqMFRWCgd9p1GViZ/Ukyzkm4W18+srT2gCQXQqXq5ddjO7+54d
8Hmto7JRgtt5/YQz1cWTZrIsYVo8NQEN0xDtN+NTYavPs23lJ8/qQKHkA3zGlBEUVouhHRtwsWeH
kTWqNH6QXMNbjwL+NzKDxhxZQFbiaSWVRjzPYnNOpCBGSmK2BPdi87v9S1CKyBT/IbWTRcwcqBEc
fqm2ek6DY/3y1iQ1SEohI/no2Nf4XBvSNjqyUaHWeiJEhnDlf2j8DOz8Lt6wpFtV8WXsRslm7L9B
iZsL9BZfPMiCDNLuJtoLHEs4PTbOjiHrPPhGKaxFm1dUZd477O6vyaAwTKI4QXOrklOCwkVSbZsP
5adWSwluMpT9ccaFGoZcjsFo2XoEdxqAye2a7Dz9PpeVxJoMytlljKQRPKt0ItdPAZOmnbxSF3CH
2rJiVTYItTDiFqnKuSCl55DUkaiWLb4hLbwk+a64neQwk4fNVGABVYdvgaiNIfVqWq1Zm1xegj8R
HXdf3NUxsVGXt2cXLGEKgD+ZrEWVASuHt03NabZKNHj3oa4GXJJuasJC4uPupqbvNfQAX6a2KaMh
WBG5sSE0lUgHmvYVcQGWjmEZFs94oq1NSdhF02vSlfyEYp7xfjbyJNfSU8Ua07Q8uHd64RJDSUX0
96k+Bk0BQ6TFrMya8TkOjIlaHf10b6Gnsy+RGXHtF9k9JTZ7Bve8Q/TeoZChvF/20rkMm/QaWEPL
MQhqra3vUlXIjk3LwEOR4Xhik89/w76vxaJT6XML7POPSPGxejYEdhja2Eyr+I3IRagxTue2A6dk
MaJWLZphx5v58OjGkaYbz8iEPKkykovf6d4yc5MbujbI+tpIwv0TBVn3T0Y4UTvyOChJLILE7hWn
jtaN3wc+090UqQvr6dwx1DHskZq9TOYcwoWuXgULIB2aMKO4O+Q7CZjOmGJTyNR0zo7rdvJQvnW/
E2i+n+GI+G5CLPyb2MjCybcJA2lG4/XjQQYgeAvqv7rhj3r7tRD2vZlCbGtgAYLYjVDRlX3ZhSdT
+YbwwxEdQj1sMvkAZ88gwn6wIJA7HMJM2G0kE/KsFNw3ME9/R62E6Fs5laNgU7K1zj7EJWXZQ53D
bNNbreNU9KeqEkID1vzCQhwy4Cs5x3YOzjcqtb15Ra2PFNT5d0B6CnvkhStxHma5Att35vR3E7sE
uWk+SD+VuH84331mQ4wp3FjyrT/md1OUPf4Ukh+7SdjYN7lEHwHkoonH1gbJiuGSMRJG8bJNj2vx
XDEvM85kJQqt4E6leh6rqTOvfYFvUQvSAPCJMSOfkV3uq7Oy4B3nLvwZ2NJvKEg4NrMC5dR+PFh+
8v+SYwwQQ3DjM1I5vvJJ/Um9xxsvPd2qFddCOmMwa4FyLOEhwfy48N2xJJ2UZ7C8QLX5fpq4Dxpv
TYsm58grmecWkXPWjp193Nww6HORLJo/QR3yKQ55/n5M0zOw28YJ77UkDX3aIqnKeX6Ryd2YDD8z
lqgSK1myoBNjtgdU30LyYpYe/bWvGn0eNFgh6Ws7wn8Vy4AP+/ghVfibBWin1VgQdUVaWA/A6qdk
CZhT9q0dBmtSJP8RisGaA4v22xV3lZ/EQW3JtRAfLKyI2ndnMypjur2/N//eD/h3U3IHxd1rMWgd
CGmdHD7NDNR+KGruJE6yfywyeIVB3+lUx59yNQ+XSsu/bNENRAkeRFYIkx1AdJOvxxVceINRpois
2/F9xlH4W+Nr55T+L8eadY22e2lBuYZa1/7ziWNBrccDd9bWWfQbp+twaQv+BuZa5KUuLQWlz4IX
8vbNzOqfedV3wVLEhLrAMU2/t5xdJqDn4bmoKN8qRfbEkgPBZ+hiEcODK6b7N/RjODMAoZA/Yh7j
xjb7Ym776n4m5JJGOq6NJQ60zCCHPRsjY0vLTrt0M5VMuMy/MQwkSI0BIocWb7ZYWMWQxcrmUW1N
PTG0Qf3Lr+JutTebTNYozR7BJywmzVQadCiwns6lSR/R3dYtlklWHMkwBKc31Xc9A3nOGqYvahlK
u26MsPSNXCVB6po2alOXw1htxE/a8LlK4LoqkhXgvdi6wr6RaegxI9ti+Oj4WBDZYj0YiXh5N8YK
VeAlGA/iGXQPtlV85ZxFWrC66gjUQydYg2khhUakXdYhOEYGUKRaUz+qgvdASezV/f3qXjkOxp6M
ZXbRsaH31ezWHc7tg6z9rcnU0xl7roqg7sjrUIsglWOIAyDW4+PEY4gA/9B8RsqUs6oKq/fxMaIb
1nCKTXEaZbDTxqrlHvezByGlu8LZvFWGVmsc9K344FC91GaP893GxLIu2EAxI4ffx4cTDgrwO3ri
3aY7T6KuIl7Kee5c6sIQW+w62axeKPsOPcKcXR4Fm+k/JZw8K83CkSx/Xr5y6Xj31JMY3/bfeVYf
4U7WUugvQUlHtufVcAFx+t2ShfMSomDLkBee834SYEnmK9ZHWXIupN4DPfWEvgzdfknsG+lAlGsA
AWWxOfZ0efoKCMj/Dzk5IgNOj1vLQLs0xY0U96SMbAnn1um+jwoNCwSSy6HqY+x/1t2XlgOIBvL4
wmS7A3EbYFBuuMVrXsCREsv2w1oKyeoWw97iIOqpA53LeD034dNC5VWk7j0wQgAyffSdRny2rAyI
V3oFGiraxmNMdTYKutUpxmgUChiJfB/pTnvWTTNidPkJHMuFzZeqMfLBQboB8j/gj9nVJnABBFdK
ZLmslFkEy+B2zUrvrun+Ace5ifnym6su75Y6getewUiZ2//gvTBMXbMqaoqrOK+Taet+uy0l3D3W
aUMuu9wiO//FzV+W1Lotrtgs7BXsY/w23YN7TZMvBfOicmZETN0YfVQbs1qW38ZdK0GSbji/cfB+
w6cAtT9PQZ5MbmGgIz2e3Pwt8BklS0KHPpIVT8PDMpI6eMXmIZNzNQNvZVgIeSnyK1oVB38elYcG
s9lhfmjIm6R7ONKWI9PRgZ12onOw84gcQRV2r1fTpVi67qQDnKgLhEPSNJvCiw71xgCR85EfOfUc
X6HmbaHSWIAz/BRQ45wGrUc3HHczzvfxLh0rVTtbfvm8qMeagivH4gTDx453RFNI1yh2D7mYVD9F
I9dwI+QTBV0NmnXCfhxxrjOeL93lV+9+/OgwjhxHfkKDFtc9SaveUTsZumAKsETr1l7Q9spkqXwX
Ma2/DNUK19hGaERFdf4iR1eEKsPYehv8RyssCtllu/3g6ZxK5OIbxwXWkgpvrkQuU33a8By8POmz
f6tNlWhJ3q/VnTwYy+h5Iq8xceeMo8UItOpyrCyK0Y3O8OB2dHSEljyRYkGsvSQJ8OSNcUUkOzZz
gtqOTW6EIeR8cD64IuVDRgrLoBxUabgHnKJ7qorKQEnyAy0Y1C9S5x7Tl/fjm8Sbpdr+8Z4wrKrK
WdlCOSTKOY2SScF3a2O2bhQSw+o3BCI4llVgzpJBrHBNyvRB1xWb4gU/w2ATr44e7Visc+P1tMyb
BLdgeRnVLiYx7SgfYW3T2GZJkbkh8UK5nsnfQmx42HHmjeeijDagyhpWNXHRv7L4KdKH/mTEE6C3
b6FGXV6dDtpfIGBJNE7QMvIj99i+SiN3ly114xlmNBB1kiYSgXga+E/VX+1AwvqwUg37uxRxvtFH
iZJtpAmFdiYcXRVd3iMQm/8YRmBCuwdkK1ZuWvufalGwVvOQ5wr3cV+3RyowaRULGSEY+hdxjgHv
VD1mlnSUwQIYfEYZyhV6KQy4sw9pCgVW9RAYL+KzkWX8AZgnPBlEZ1QVyKPguQo5wFm40YHJIKDc
16rFvyXfx5uANMn3xnbWm8BYvcTWGK9Nl4lC9lihiCNMlh69Ig96Gc9ugLo27n7bGWxiiuuXyZ4h
zBvHlRcWWQNdYGmd82PWJPZngBlArSedqB+dOX+CBmx13zzZ5XKKiEKMJOJHbRn+Kjt23tZLNfD+
dV9L9n+E9gUeJQ8HhaV46K/17q3ItNhxd/z2JBp2Ja7m9vXHuI1GqJEY5Gl+h/VGIHVNb4OoZ1GT
xwJDB9r1FbJw1wrK/bCIxL4ujIdutXQLtb3I2KQlXixnwoDfkBAgB1DGI5O/dQEmOvDNdKMLeLui
1gTjopoyKmmWNumzhmQTWx8LrxAAMCDuh5yZgC68/bZdUM4ozNU4NQO6ncCYBDxME5f7j6m3Yxrw
Ln5bPYhpxFmKwh0hpWNO+YdoADPgSZuD15Etl4qQSexicnlovNeRzGmJ/KYTrH0XVNIGr2UQhW4o
ZLoC55YXQhjIk8VtXUNtoIscaHQe5DZvDD0at5/OCt+uaVpdsQU7kxmW6FLuhit2t9wXi3XZM08k
UyAX159cx7drBk2iuV4q5qzpRmqyEaU0htEVb5jS8iWDgDawFwVm+lhxQiCrQWe3pTC3hWCHadpM
HEvGRxp50+mObfiD4gb7fgSnyOL9poRSOjpGT3K5iqBNOj/L91U1Q6OtOKdVusn43+jgg6UO3i4l
fKC+aqTgUeTo9KBToSu1F5VGbPjfEY02WCXe2+yDusvMOtGT/f5t9/mFetcBrqQERGg9JrwLqTMo
SaPKWsJbwWfllbGOIWs/rpqt8EW3DgkYvXe1mwfOY8RX+5C4W/tU2TJ0KCI62SjiB/LVKAzpn72a
gjSnfTwg3paV8IAJ+5IWs46LCIE/gSi0BqHBdCfAK5k+hfQoEc9td4+e6gTV6wRxiMRCBUdDT/00
koxdIh7nvK6L933dryA+r9I2CEaV9FIr51zDfuLJTcZ8GDCjPjs7yQ/IPxkdWQdD3EK6iyQ4gw1n
HJI8w3FtLVjpWfLSao2NRn9KEBNubbX319bSh0wmNVre2kxQ8DqSFlHgv89F87r+N1DxNI+sN8uA
1+oOWB0IdFvsqB12zk9mmAXEgv5bF0anpPrRwNokFRxvWXItAUNKLvR3m4yVrv+TYJds6pE/xKwC
zurh7Lk+QIlL5cTKCm1RcO9KjQh2M8feOeOBiwo3cu55EjCRCo7B68g6HVT/nLOyOzTQMxfrzme8
X+ZwQaknSka23ZME2NV4JEqRGZyngEgT5Slvf9On5hRPDe45P5GO1kTkA/ZjCAsCqEk0G9E/4Umh
fRzhyNqTamOa6Wgs7S1bnlCulpZFooaLOq/FJ/7yobFXULG0XjvSUnSSxaI8v0nKeujh4Pn+pNJR
oT5LYisXfocWg51qtPfwS0Z+IkCj1UMDbwY8tHpQWMAk2hE0AY517eyr7sVUy8O3f7lkkv/vFGDb
ZDw1JcUMgfQEu/ocRifYQtY41oTN7Q9de9pkXe2XC/wqz4I2jiSc7A0kXMu/EjjbVHQWLkALyKAg
CtBAgztUe4JefxcgHtEQywqggnJDWuk+FNZkXZXl9dcTNDzBzT0pyPXMKUCj6L7/slj4pnHsYwr0
zt9Jh+4HfJ3M2IhZG0KHBa+5+6D/By7DjscfzWdaDl8T3DT//Dei0so0CLPmB57aIUJJZzQ7V9/7
fq5ok4+DZzzhHtzSQzH+2+oB9wH6ShPgz41J1hn5BGaTnwozDC9n2rpzpSTzNLr1hSApWH4t4GTk
29R7DTgWSU2JG+RGACT5iAHM0ui1VhyvheLfKm6CR+h/88acpX+LaoCo0voWP9tswOnVbXc/w06z
l96MAcVxNBog6JmpuP20XL9fQCiQno0wbwJ+rDKBMWeAebOzPrYP/KaqwiJymRCDCxxPdLAGAgPW
7wGUhRX++4fPqg2if6bg7f7cQ88NBW5hmN+Zu8LR6AXAqEuMkJq3WsiNvHZzE5ZA8SnQooj1MwZb
NT6nU4by7oiycwYIVNxuPMo2RNfHZdy/4G4HRM2BVAB9RaQYBy9QGNVRrKg0L/jAhArAa6pDuwb4
ORKuS3SFjpUSXHkD6OUG/Y7YdNmtQ/ldECceiR/d7yk4fxPGFTMttKKlwMnOsc5vUs3dlFeblP4F
V8nr4PK1ZNOClJQvEqqrg531sU4cQ4Sdm10/uhormArsmMfZCO5sGdOKaJNRuIKidoAPxhXQPB6w
6stll9LoNbXMNihNmQMiiVr7sX8j4juNVihiGAMrZiVZBAh4JZk3C+t8+aq2D4FdWlZrOkmADTVh
DOx8jdJHSrdMqgh5IDXUWqypeuKD0p/ACA/CmVYbMFMuDDGYcJCrtMxcSuLftWVQJB7gw99tKqyS
vkKGSqpoP5bA/Rc7gS9/zphTU75XWdSJQG7c9X37+5m2uqKxofnsPI+X+kKKEkiPOCo7V16g7gE1
bkX1BT5SMSvymCOraSe/9jT0gfVUPNMgk5Ehmfj6RDaEhNqMLkMCNeWn6b/+ezsXSAKv4GtqUges
hDRtdKEzxzLS6hQ1YFktqvQOBw9XXsRAf7ClX/r+AEktqBld6KteChRNcyrymcrnHV440PL+f/sd
e1T0l7AXHidOmSAoRRmwZQm973lhApxiR7rraYjrmONLw0zi7ZljOl8Y96gIW4rtF97hX6QaPneA
w+w080M9dC9ewSPu5k3fuyJYjBCP4s3aSidccfRQLIrwT/EndSt7l6aLuP6g9clFEfvXCjfRktL3
459Zthi0Oo+Cu1NNfoq+pbKl61z8Nl+IaisG8bbhAtJLT1I9L4nFEaj/upFGfc4hQDIAsdEYCcoW
rXZ93g5qayHTMmLd2Cqew2FQvLxeLz9KbXlNGDpsaVwUSEEMvE5UOcn7sQtKpFVhd8F+KW8W2Qcc
kPbDehpTPNiev7BKXo1sS/MIC7J1r8IrHXzAk/UPGi1qCZ3DExGjtNkaBXUyGpIhBktOrYMM7uik
BfQAMIYeMopVMCYPmkIVveztzfibj9zSl7fL2mj5aGSYbuv2nsJFr5J9gXw7f/J8T6byTRvHAgFu
UwKh1V60Rw9zn1rxwb61KYhjcBYc2LXGsC1zIVrg3wS+92onwb8oy9hU45pysR1VafORrg5gcWb6
QDPsYlmfyi7bFBunRsM1AZj2c0b9O7YTFP0C2xJkCdfbGxRFNJpc4qhS4RUpnB/xpn1cd+OLa0ML
LnOhd0opmq7nKM65bi1W4X8u2L1rUy10UYRjsE25FjyOZwJBgrI/TVwBK979muO4wDLX2KEOFZ/C
2Zsv49B+qJLSoG2bZYX8boR6AOGwgRWt23R1hIbqzPamuBwBzWIX8R4nP683sd4Hbf8koECP5lJU
h1RBgZYjnSTpCA6EKgOo688Jtsp/x4HSe3Q3D7ajU7bczpsS+DZSbToHiFLGXxsHq8yAEwMXNOfJ
XiRzjoAUrhkNbDTcNhZe55wyy5DYuSfV3X+6zMfYvJ5K7Ej8JjAMuz6jZgYAGJD/mKLXCWKWZ8Na
x4E9yALGzQ+JwJblFVPIBzxf5dCFZ2Idhhj8fvXckMiCuioynMFEbmbLoOxASs+tRcasBq7TJkrN
KbcPQebmMxBMuy/8vLhc5YoUMyWdzCqZ8ZGYK5cOyG3Dwrv1suo/2s176wd6v2Dqs/kGruHILAvh
+hlI04+SFePzzCyOyf8rCLEjaQNCnOozvbQgL3DSPzK9Al95iRj4kf3d+PHEdv8DvbFWW61LoTWy
ndpez96CEP9VbD9YSV89xhtnLPxrGAIOtFOjOIoJ5GkUZmhhQJtTSleCfIBxq6aZ2c/QdshENv7C
iq1tuM13AqQUeEJ/3ngb75mGlW24dRPM5i0189gr4j8X29rq3e69eWfB2nus3iRXQgovitCqzDJx
DdIaEv31vhQfwpIHwugegM64C93l0zRHDzLdohP+xmUG3tbn3u/O7FkiGwBfOp2LQLxaQcnYSkk6
dR8ALL100ddJ3zbod0aoZD5BgB5p9NhQ9K3tRemTAw4QvtlPAN0e7vx1iDQCqLLGKqVWfrSX/Dvf
IVW9Jlid+3+ptS+n0hSv88DHLPDbRpwP1VG+7UrFZt6GC1c10eHh5gT6kuwUdjkF2L2GW/9klxPP
/XmK3eHcepPDNDjFnG1yzMjYkMQKKjmeKXqgg1Fg4Ll2r5eXVrcP4/RQmAk064nVRn9oRd9K8xHl
+Ws/b2oX5OVEiJiyrdecHm4ESXzZdRKYYFFnWQXsHLAZqCzx3iMpgJt9L6zsbosZlG4l3w2a8JzX
k9S31GYxi5xMduDa/TY4y9jMx5rHncruNCw1PC7cm3Hnu45UcwEjxVL0qELeL+VmKPEKp4ZP3O+W
2YXoDdYm6iDgLBqDqMzx1NLFA2zPQLuAPJcO7v04Tt/CMohwRlaukVUutuvVo3Rjpy/GzPYYL6mU
RWauceXFIX07fizCYWhVjhS1tHHaOHTqwSpdV8wke4QTXS05pqnnnNYt/44HIi4sY9w/PnrfN/AF
n/ulDAIBSDR4JnC9SUboW9B51DmaDalPT0wg7IKx/UusweCCGO1IoGoPEOoJaECM2YX0YAVepl2b
/5OnGIF3lwArbMfhSVNRn7RxNR1dmt1YKuZpY7ht6+vY3fCJ2uyvJ0o606Hm4S7EEFIS84HaD5X+
ZCA5WlxiH3PtyhBV3L4KE8vZiA7+vCSqKgyCfwM6htzdxv93HiUfOrs/Cl3n/zyROeYEOxd67K7i
FX1j4XrKBgG62WhFRTojp4TVfoIGAfMCQbqi9QKNGdKewpTVpgadv7T5D5N8+H02gA6esxjTx8PZ
8j4R6Evvt38O0gts8/xDkE/THwBoA2JV0Tg/kx9iSi8S4KOd8dNuqLcPI860XoPcZ4MPPRRoSCrY
WF3SGIdsDxdHcJoIwtUz/oQT0CpwfmxBMKr01MGUekmwBL07eartA2FA0M/8R48Z+E1m3RSDSNOd
WXe0Z2Tr5CMht7MjAWO2ryf/wL685mpdPRTyAeUnSvP1u3UX0DmQ4a+JsBKuKRuTKPGSFy8/i9O2
IHSWav5UdVsLfJSZkIspneAykCbH8VZK17T0z6dVfI2y0VDo4z5q9VWBsdV2Z/UJFCobW4rJaQrx
MIbq/LLJUthTLWOo0cRg5nMOUK5JLXZWbzMu7+HfR9VtkOMCG0v0rTUND5RoH5sdBzJNKCYAV0yg
L7WOwpnclghZhkX0zZJOlESNA93K4sm3OmTQGIy53z6D4d5BGjwRCRVWcfc63yoA9a1jh+xhEn04
oGW4QeyxWsVW2yeflWFyJ3uwTMaXFbYxjMMilP7h1CqJMmpzBua4as7Ug1RdzZqbyEcro2Xrhuz6
DpdYw0vjQnzeMuH/ZxrKdQxfWZoWaN8/+uLJDVz1TJ5HcM/fHgqEwdJuxykGT/wIpnaqmZm9b+HR
jy7VNXBN/UH6ta+OXmyWa5sfWupx3VVs8z5Yp6GnX9B98IKbk9C6ByuqDaeRPtoj5tNxlVTHAE6E
6bZQ242Goq1qSOViW6NsOyRBi3TfbY4Dda3yahRNdF+/aV+NxRFwT2CRaiG2Nb+fZr5M5ml4YjFn
l/RK/teFPQRfdCHrPV4QvDrUvd0NSoF2cCOhXLaY0mdv1c2i++krY6zInwHOby4XkIFbHTWqdwLa
HGHqP9NDxkCaXE4+263XcBrdpaONneMc2ank37ukRAT7JcMnfsHpHqXSLNk3oP87yrkKtrvHTIpW
CHDYGajo0CD5yW0QDrrgyqNWYLvBtK989BJIKDPhETZN+ferr2z9NVtgZhREFbQu/8RzizYvZIoF
igfUaYK7IM2JQ+xrpSOGWUI8K6Q4e5D1SQRUin0LF7fURIEEEVgqLi1NmA9U3kAXiorh5WO5+y5x
vr3xaoPYL4lXzkU5P+v9jzbqp3QE17wcHecDb0XZP2cSk4p6nnVFuWok3ZFea7naUNYHbXqj5ebl
N0FqLhZVTOfCQiGveQMRtfFZZElDmpqY7DONB48ENrO6mvJ6g6rtTUrc2g4VJGdpa9/wbyDUobkH
hh9RsvPB7SfZ7OT7SF/y4IOe2+QwxbJPSwpXppmhwF3xXz43IIIaWNp0mV2a6YRZ5f/Lmue9nRsc
LYQvGhefj60b+hGNGtN30MZew94Cl/ZLtSSc87gZ0FzKef9aWQHYyWZ/VpMNft3aoBMdt5HoYA3k
soSsqbAcEA0RZMkfFgKjN8GBxtOwDgdGlKlgG6hMj6V1m114vkfH44+yulqLF8ZjjKRYKaCNkPFW
a434+HQTMTNY17IJtAuqY8JYeExRBK4E7/nk7dUpNgJwbGu/YGFyLGRKKXLj+sFkC8cisB/2hWgR
8xz/qqqj0Rc31obC64S2scOEmYMo1nFcRv58lLx7RVuU3j19oKEBVm+3VysOovKA6jDEDaO/6hoZ
Mp30N0fYEZfQjjCAPjrl5KzDs1DcMA80zj3vFHyEyTHALM0JBCEJeiKMdKm7SBsMlRbIeoRd+iyA
AUM/I8a4UfE/epWwpfRxvnB0hqy/HsvqrAYvcoh5DE+7TfQLk2ouKm4ZgFP6x+yQgtVYxqf/EEwl
Ut7ljZNN29dOeADR7LX1KlbC3K4uLBK0c0YZXrXhNMJJMarbC9eh/4YwaRaAuPdgr7xEMrE+losi
p1w2kYFUVGIbGR7hCLFXZFPJibVWcWBpmDC7QcazJcc29TgFjUT/iF7swOX8FZJ4k6ghqSOFqcff
IH7xaQIRZtmnzorxjBB8XXok9Yd7tLF2c1h6DKBwvKxNIar/cXkdcNv4FxusHxUon08z4ipK6KcN
uzWaw/zApkWyheC92d2Xzd2VsuADXLJwTrgZXkE5xgTI1P/EwSstOkGJYzLfnBnbWBgmfcBdGh2x
9LuA4G9TJHcBxu//lNXo9LGbkswZK2YdDt+DhoUJKT7qbMegMUv70iSGmX7baUoP7tSOvqoRzH+b
xF2cgMpjt4JlONw1Apv+TqCn4bLcEtq3wvomgiqe/bRl2ImJZzFwBBE9TdtWyY6ADmpOOgLWr64T
/YE6jIBbFN4W5fZ8N1GIwLNtj9Tk5Y+9itYAcutDXvBIxkwBHDBBPpv9oqO7nMVlZTLhjDhfKpdZ
oVMHSLxiBnw7XCG1X4vafNc7vBNdQthu7XS0pSBo/3h3AObhPF4WE5bVGPXliGUQVzgkPr0Eb9NV
5yNoF0exJBbnzS4NVWu+usAYKX3LV+SFvYqFMmftW0PEW1SznLX7aQl5lv7UKV9norjhfHOfY5HJ
ZtTwugwPxt/4ms3wQ2zvJ4POkffk98CYVQ+Z1Az00HiAyCLsD2d38gaZVe0JzCB7t6KCE1VKGUHt
CZDFtgPBr9EAXp0W6iSFqSyueBHOhVru5VOW9PS63el5WXFclTwZ3v74W/i7mc4mQ8k+oM2oBwu0
thF7dY9HpOnqrgAHLoOHb32zNJGaWzwk2Skyi4fxAIYwO7JvhtXCXtnBxI1kwRAqzZdGOPCsSpVe
mam/umWudBxD9QKJKYbOkSH7Ja6UqkuH6DZ4CjEnbCz/Nq62Kuot5ckslJbUcWhsBwp9yjf2JSJP
IJt45YzqBIpxKTO49NfGrqaK9pXK2iDJPvh9mh0ACQUFiTD/Ob3s+abOQl5k1Qul/iKsZBdeMjX1
3f/ddfYPKJ9Hi6i43Xppo41sffTOKG1CN1ksI5s/RxmTeDUa3ckFOV8oAtTTqbVxWMZKzop6xc1s
1qyhpCEM0Q6BrDzjxiUcN4uVpanffDy++/Jkw65I3cWipZpcqensm3kiw8cMuSY+m+GqGvfIXgxr
yRxnCE6SycNwGnzHa5amqPNSeosNwWjJSNj/FOxLCnZrMqCb+kvyUodhhFnddE7btJycx5B15MbR
fQ6bE+n1FcDmaiGJLNFehLi7WPALZrlLm6ZbwYkG3Ql/q+Hiw9NYbB6l//nNRnjCiYfhGtOx33CU
kRq6deZhQ652HZ9K2GWaIM64PIlcC+q+eRfz0QRLmapjyTYV/mYXt/ll8yLRR2vUoUYzN/REYOwi
1twO6Pw1SxQAfZM9nd0ZG8yYhmcK5wV29V5hEsvb6aTGpGpNVXwbfsSLl5AM7M1AKGlO2aBIkapr
XDavaQnWKt7wi5b4xeLzwhysso8vu9eoNSO816SLa8HR3KVatWEOOZEgkg+tfs6+bLdTqVneY6+A
QTTWRF1uUBNRYpITYSTqENzWxVbAh9pxGwnFwoD2h3kXANKtX3PEJfGajaHsapkKAJYUAA9PCMKM
sRUrnZluxyN3QTipDuK/yFmX1xfG3NUKJvmkiDyyxbBHdBXitiFzolNKe1B+zZlYbID0LOZ0R89w
uVBcZlajyEYYk4+eEt0FVRwYPZ8M0UR9tmOUJgEWuVy5ALht00INLDS/dzLz03eAzriS9snJ/oI4
Lzs5mC/QU98WNcEOVGHTInbEgL32fX975jhYQsHba/36HGACgpICTcTALh5DhWNLXO7dnBJSVS6k
hu/N6uDMWmDGhBSTjO0gk6UOCayBLVnXeAE+4anlCazbNKfxVzMzG+xZfwh1lfIbRz9eyaFgskRA
6xmBtzjGIInoJ9I+bXGqxxpt4Ka7yJBMLmaBzZK5zFqKG+0W8LWMPXEE5dMXDFHn4mEO5UKgkUuZ
HE/tiyL8VAiGuG4vpyicmyOWWwlGbiZO57otVDLMIimG9gZI9T2/hDr5U8yf1092NzfkTilwBsFG
c5jAjZ6VWMFI1HBbzmFyY++sWwyASKAs76mn8QR6Olt+Bv7THAYeUYuTwU28vHSJCfB447U/oQIX
8i3O8W7RD7sQYc0hm0FZUb1dVXLGfnmCGupFvV26F1VdfM4gen1uHo9uo4gzKuqB/hh1ULWjfVXK
cc2RF2MLXS0nmJDPqiNgIBsH5Ryck3pGX5wxIL7IA7jhaq2egTTTj/kzDXZwA4jEwndzjoD8gXRG
XBgFe14bEfwuKOUkKG4mHOBEiXaYZvY4meAD+c8sD/RVj4DbMCdbito9w1hLM8OPw0pIqjQrp4lL
Tn9nVB5wyzbr6+hkOIlnnBw5/eSL8LSKymScrud/TBZBIV8SrJHgmPmqdiFycS+3Z++XF0Ro5tV+
2YcLRBJRwnFaPlxG0ToGv4kpAGM+ckXZe/0ftscB0epjH5yPg3nH8InJL1b1nGP1Q/fNpOHNaqB7
eCTMVTRo357g49foV0FardVATs3dnrbm747c5GkR14aX0ixYZMpbDcHcDRAG4/G23QIZOPVNlh25
9E5tzaHgNAmdsuiEd3j1sufsNfDMOQpg+VFrz2wllZT+bLeHDjKS480chaiFFhwCL4hitLYeLWY9
Aljfudu0ayE4c77pNUFa1CS7Cs7uK0JNL/9EXZsmzsCgQnT5LzlIzEYllg690fi647pElLw12RC7
BgOvKOSDJqfM2OUK9Ckxus25FUP/PWiYQB/ulmOwVc+XDIt/gkyVLPX9L17LHwECOrMDdg2N0buo
QXkchkbUHr5L6tiF7pL2b5MQOpDMbuN5id3NaE0dcvLQJNYuBKB7WTs8BAbngHvy/oJ3iSTb8O0d
ZdvnrasdjiyrqG1aa8oNL4V31F+uxfQcR/Zqi2PXibbd1elGC53QGuTnJCTdzBIKU75b2s/bqQYj
UAqciUiSezYsOP8CrA9r1kHfWlOoGvJ6hXGdaCTyPt/ylvfAuf1pw5eMy+gB2KxBOkzFxHxTQ2HI
7DS21scl5WsoCVIFW/qcbwQdnKEOtAgOanw3ieJJ6CbQxAwjh/LSJpXmmlpp+pWdaxETssgBBkrx
gTVWt1JfhjQ4nDW5cwJu8kWA0RKGjXTvsAyI525/2ohOrmPVaTAM1mBa/Ze0u4t4qh+BdIZx8L2S
0S5YoUmmvBUaRv2Jo831rnl7wCokzmaGNfaQ8Ik402k4y1lLMc53LFmwHMS9nDss+PPypXkzCWP1
hiAj2yUMWsuLp1AxzbhahOWkkqa2dtkYcdX4t1t4XZwuhKirFQaZGnckshbf7EXVzppqYoPVUjHE
SAD8WbrGLzZEJ93mpkXeb7UQkau3K1RnKSV8O4c4gPWhHWl/1+Hr7V/PSiSmxFq+Y5CezUpax+S6
pBPbYi37zIgyJKDHH7XM6EFyhfWCb3XUFmtuZBuuYWtRRq7z5TxpR2HWj0oOXu8bUZe7u7ra6o1Z
eBr3f3uMCkHDVNNLTdd4lR9xEvFEhrQgzZoz30MFl0Ss6w28ufDlYoWYHvl5ULOo29dxksQs4QUK
qYYkSa9TK6ge/HyBC5E+9RaNLegnON5umCHUsMobPyP9KXPFlg30HjcUL1AIXSydeIo3WU30mYRY
HrN5WPd9ef8M5tkNHkmNVUNVtmi1fzSzyyovf9Ntdp94zZfDXVQ0n9fWt5n+2HfZ1mLSvrPJyoHm
pIRHAouecTGqRoBjoSFN/svHEJ8CRnd0MlGHkde79yb3xlFl+u2NA7dvy0aEy2nDhWzj+xYhKSfi
BeSmUwmPc/DLsvAmGZOpZXE2VqUufxutVJLz0qfNZrf6+5d8c7TL7dpwaN9IWP2dyMikFFeNjfvg
WaK1dWhPwGB6zgbRumk/3QEUq0JXBpHAvjmiFrAWHYgBvPjGWzTDFotE+GjQXerHy2P0gLENUqpr
EXJ+gEQ8huskifOdDxU3+NzKQJWtY3xZkwovtuPo6DNB+d5+No6DIotVujbtE/iskOZD7YHMvFaV
ur+UM5q48OwMs/ANOEuQfCusspCmXYnwJXP3+f2yT3vHOACPoNOl5G7dUpHykGVb1vvB8usCxvTO
DShBiB2PTC3bHChXkZ5pJDR7tmlcmJwOrDUMlgLRAFuZqQNnQ61YgG7dLviEY0hFREijhzrJuXr2
O68VkGjkoMvdHZ2NtZKjENYhRbMLy5/ez2bml6lzeT0qIy2okTrqUqM22aUaCdqJ8momBBNFRILf
fycLIpUiLvBYGQhW3vQTdDxEQedsvDv0re7f4K8RbFfq+ESdM5dMhAcZytLIzTqz1MfUVYg/cKtz
CC7taqLWQOwY3C+MqylYShGvhgaInUv5vnnfsw0WQMnKxrZj06wirn+lI0c+utsx4pFrT3/bYkhw
PhaA0ym+qcIL5dGsFXdbIYZyA85XrR98dyB3mt98ieLa9FVbvLJARr4dl33B8ZQHN3z3XErpO7Lx
/TFrPvmw6J+Az2qnM75XXMgCs9YQp5Hsiupcn1Tq265jibKM5OWeuR2P7Z9fg/mdXz8hNmFC7pZo
Ui2nohbmZ/tgjla6h5vB6dMPT+pehz2yFbuTpaqurXLqbAZ6G+YzV9lxszF++hks1LO2wOBjzfSV
jLC5NO4wgfbQxR3v8Rv+a0ANv8rnGUmrH8ntEkAU7oTymlX4xW0qjMVMTtcJGnuHnP8fGMonANUz
LdiZipVud9yWrZdx/TjrxOhBU3R53xo0VnQkf66/DiTnxjI1jnV92+ncq4MncAebNY9g6h5kVtep
P+qsFXx2zBc7eAX4MILIuh1z5ef2rCE0ax2s5cfkYbUY69Z7gqI4V6E9sY1efDP7iSafp6UHSmLE
lMgRmozNVHWthW5i//Txg+pDsrknZzMYYLZtQRGzWcwmlRIHer54qPIT8IJR5X4tqwZU39X/gWet
LElOOySf/20wMRZ5o2Pys3yYrz6luOQdrjcd8S24HW/HmedZCSaY6KQ10D8alIkstFjQKFUjZbkg
cuXGdBORS+VY8QP3gmthc/rXv3/CqEUPI2ne12Cpi7FEMhcInv1ylEC+hSMVQYxlXAzZoz6v5QU1
Yp8BqnZNnzbDfORT2KF4ogtlMsLf0j0H0Q4iRz1pRf7Y/CavKYPBffGlNAUHO3rfUxhM5q0Mbbvl
zeHZzGX9pLrKxM/YnfsxLmVIs5jeElYgiNwa/3ZKM6Gg/z4I4rX1wlUUWrO+kZ8taAvKJ1DfXe+6
7+ibzfdkpnDDiOPcdV4g47fxbIWmanJaQIZre/+4rxeaxHlrhdQLvTvH54cCAv5T5en1fRxS4fhf
Y8WEAa/02v9oVc041UHKz6Ofn+OGPIzCJvu7BVxEHSkUJ5JKEV9FEZblTUXqKy/EIBnH48X5TORW
QfbLqKCK7F7RCkHl4gxkUabx1mjWcsO3ZY3D17tBvEEAeqp5ciWvE2dxN+UnzmVFrwuMgsENM9qf
Dxq6renfaJQgwCv1BX60JySaU12qm0oV52W0qEqg24UIq4+d2MTrQ2+uL5RLVdaM8EClHE3I8ZyM
2fTOgItTDMw0dCeDWdHkN8xQ3ohK7fAXZWpY4obTeKnFUhNGj/kejD7XwggKaqvK7lUEedKQ90BJ
x9KO8GHLZM5u16i+NKzUWkO4NCjq0yADDmAdgqNUK8QG57utmVEb33gOx1rEOfqoFz742cN/fMHo
duea0aQfwNEQp++orj6JINv8gS6TkNlpMV+go4phht9WcVXxNPyqyJQys7auqku8ago6XGbY/WZh
dlPEUQaWjYs0WNjQA5IL5yW1ZfOCQICOJjnm+zDwRhCqVk8tBYNaJfGbOtoLSwsarb1Yxde5d2EH
IKt9MT/uKts/H1itXqoVxY/E6trgHexwSDVo9WDEX1qjeAiKl2SBq6pykGhM9+dxEI5tgtfEZIPg
OjZBohegHSPAdURpdYdVBiuK05Zj4GXXb1Pz8UBPXikRbKtDsPeO9V3TOAewaawWDkdcKpjMEn4e
78Vvebsw9PvFSH1AgTmBwud3kQFerfk8x0MNqr/35wKmWtR9bUZera9W/5GLY7RB8BiIWcT+wY1b
9PR1RVaOqzE4rneEv1+rwtSODcowE0BI4OOsGkSZHiPavcj9NMrbBjK5UKHxkrHxM8LP0Ou91Yyg
DyKHyTfgYTTknD3pjKD4p8upRqKDoVZ7zVWd2UVgksnbeJhihEKQ7gZyRDqhw6rZ+nckBWB+HpTn
nydwXSYTjmMdDIq59OEqTisahzkn0W0WizSEx3dm1bwtUBP1O3LjerMeASEixKPYvCMgI/5Darn4
IA/nqD0BkkR8MHjAE/Yc5Y6CZXlfRFQ5CFUBJTmWRBeOy4yiXOLof5DLfFkVMIqv5lWeCeGGVy1+
FohVevs+ramNDScH1fMmIyRQOEWeQOMEweNavciDfKiIZKzqBgc4WPVnWUReSUDrPXtgsAh89XMZ
7eciTUYpNQhhhpBc7HW0wDEDXc1/b9r26YWhbNGU2ZxhJcL553D13xglpRDLakKZdfBtkb7YGnyY
+EhCHE8wiBLkdv8xmBuQFIxxp4WuqZeBTEtdMb9eER/XSJKbc/09xFHT19ZJaWvSHdxLRk7rpPka
St3d6cTWLMFS0nzUj+2H48OlgrX5aP3dXw2Fv+PK0sDDgtY2jsEX3C8d4Kgfb6MBbofYujuY3y69
Fb2qPJaB8rYtfm8QB9VqbWB56L/PAA2XpCfSs8ggtqQTy29Kio/OZ++cxEzWG/hojv+azaMDswEI
DjUnNujot3qRtEaQ//wEKHeVlO6janH9kZNQPijmpck1M/Gy/gS2D+15a6b3r7fIda12w67Viv8A
7ruIWP/e/V1s9bexkQPev+RGoKe0jyR3/wmilDWMqesRRfMbaP5bKKp8kQErSnvnlzMuCirPn9Nk
dJ+NTshxFRW6TLsMM9xXK0ubQzoug2kMuT0jI0ST3M50hTDNZMKkWv9JffY/PvOoETi+sDyu1ge2
bphqz1ZKYfX42LpMswJXnJwRLH+xNAO1TVamvirbkrywOaqTn3h0ZXQ9s4nDKNtnILb5+v7xgXvi
8GDq0D6KO99lgOe3IIODeQ43p8WFSM9wT8WGHCdm4QnmwTdzddeV3Cc1UforAEIusKtVeik2h5QP
eqHV1YdJN5GuPK8YO9Q0xefxuMiSYGxA6ag/8irtEVha6OTvUezsVhR+Qo8xbXj/+0k6PGO1eJrQ
kMzTyEaZ+Ifsz/id4jOpu7+8KXwySjc77FP2jD1yr00iUI7zJWMH9qKLWa7YjgtzZLk3pCUnbHqS
bl3J5OXplFzsVnmcUXA0MiSbof4AWHgHuc9w2WjXHFAfSiKxsP31QBeSYbgGPaDBpmx0NqO4h8IB
oXPKgmBGnNb3X0wmIW14O+gRfM/yiRU4BlKChCFoYQ4QswxTHuijSGfYHHv6iSnmb9mAQ8Dzuwa+
hRlYAMmni7qp6oxwFPgzYdBfNSjX1Ue/fMctwKxIqnY4RA2Dexm991jmshEuaPc4hqVnFPuOzVyJ
V172BLbi2piVE+bOUdtspHMv63PIP1j5stbAcY4nI02IXh5T6IkdFLHfqT59JKjJS5iYA0Pr/EXk
BvhdRyp82vRUmbJUq5Z/p3VggiapZoCu2be90YKgxF+LKZ2KKA2+gBlROKfHalnPZRD507ofWefI
fQQcLU41Hp6+YeYQB2KQCERstEtMsDEJcYunUrE+kzcd0HNps6523QTmrdqyvVGa4BOMKqlxrFrx
aVNyNH4liS+Ejq2zr26ihc6920xyA2HQmuziUQLqsebOj8h/obXWKo+IbGbsD7BbMrvnu3nVQN50
0T2qi5gVuBIIwrSmARU7TrHNFtYxyVJ9Xd/qy9srmTcJD0gg8P9dUwoKIgLHql7T+mB+gpcla8Ma
K68YwfK8wJIurG0xCos03/rjsIYt/I+eHgetLYaqEJ4Cs3DyzoplFnGmpdhxvzWJEf6ibxZKXPUb
NXZDF0HHfM/0xEm7yuhJWXBJFOA2Qf11beoX5pkwtJk9hcMnt330WjfajVHAqk5Y+GATdT/AZXoH
cyjZtGtjuSFGUqD659NGv9V39k5xm7JkA1DctUXYF7UbAafjjV6/QQSaDmawSMQWph+gYfJ0sKW4
iiFiRYioQbw4bmz8SR5Xx+aQtL/VtbaYD0TeyHG3KI8ikhvXfFLciuO0OL9Q36nNxpIXb/fSsO+h
51R8vtiHjvL04fi2Fp1APdG5ACqydXh0vhhRaeBnMtoUMdKMakYDCeyZ/a00b73hb876cGZIlfrB
vf0tBCnsC9eI39vgdsAiNDQw1l6E6giNOiWsHRQ99poKKkYaS+ucvsf9Jed0HJQj/mfF4OPsOMOf
FxF7q5pb9gxKvIS9YVI5Nr0XLinVBD4dUBTHXpms/r/CEM8Zh79i/ewWMKvXhItKd6vRusaeot6t
9MXtfiCtezmeVJf05Y0dP7grccihIvl1IIzrXEgpDkVxGf8A7mOQGH/XCFxy1QDTtvEB2v/GQuVH
n9DBe5HbeCXwRSsGDgxAf7fp4J16QnHjf9pZH/bACwMHHoo+kFtkRIDGdvhhq0HUyZZjyDnCnd/g
pu98E/WYzDi91Pmts4jpW6DfAH05H7ctwgPTv7AQnANndXuBqDdHTUFg7cQZURc0tIqAWUgYNxHA
prhPZwOS5Pxtz/0Uvl9MUeKY14+0Z3jH7t8MfWWmX2uiaNpQ5PDoC6YUZbE3S+Aoau6+MskgGWgt
PZk8CijOQ1S82OsyOPsHAHVEHOx8VFhh0PTn00CEeuFfaZT9ZUBPsLv+OmjgEtuPpH5kC6QYGczN
J6KSsZaIAa+BDUQxlLk+mlXJjpcfhtxRWRQNuveuBm1vrYp/8645zAtP2SpOOVpKXXmy3WP9qOpS
7ReyJtFijaTg54IPN6ebSQkr6oPJudAL3eKYRyosdhA4sVWGkc7G9niyQ0Px2Cb16NfuVDj6eg3a
P5JJC38qBumayAN5n2CBq07K1x2QetMA6qC5hnSm+mv2bI2yTSfc3nbMLKGfAlHFlDvetBQOEKov
2aCtCLUMVooidh2YSG/Od0AvhtBCfP2L/efAjLAL0CnNd6lmqtpxa5JVOICwhcVcMUJCtwTOvlyq
IPomERvKuERI5GUUS2wu4SmbFzWNc4fYNeKR8lG/V9IcpMLJAMcPmovPtinMhLoUmfedy/RBWDxt
iEsTJQju+W+2ijTLs1DdDI85IRu3kVwC4jduOH2OCZNBKZgiBOgjjzAYHLb0MeHhKUR4e9ktIcJt
VUQ+yCZ2DnWbjAl1FuyqjFV1UA9XIJlpNRMeEHBpsFmRotTSNBALJhCmkiGq8WPNTH0UHo2L7Vuv
EvHktlQ1G7HKdnc2PNi9iPEFvylheeNEI5PnZGOIBdO0LA0xAqKsF8DBc87BBht8kZCOe+NQIAOE
ZlDas+yvQ5TTcZLCVLzs1r0C3jsrZZbDMLtW+qL7qkiQmZWBiUBBmzWnokxZU1bAJgYKb2ETiNVK
qTEpgmW5pyDJQnKr/VbcAo3b9BNo1+hpv0xoVyg+bkyBbw30vbaJPwtRFOSi3Aouc/9VaDc6N8bV
Jn3Ja7bO3gw/9ix2aitHI2Bk2tKioMD6wGczXWVG6W3dPVHAuhDDDUWWFN6mVsA7HzIBB81csUNv
omhcwImWpE8bBaBQHXvWDPE+s+EXUQb1aYsSeZDCQFP8Ee8we2gGObdkUpgEAVpfqnaZmTB4dPug
VIe1ibngy/iFUKj8fCSaOCUPV6jTesfWyfQU6ZG3XbV3caMZ3v7CmPmRdCuuP7zhcSkKTvAONiXj
fkfu37uU5oG4v0y3M9IZOYiKxbiZt7Egonc0s55UOWIYh0L65sg1QDkfX60vWeFGyZ8RP0wcHjwI
fGL+NAPZykEAeaKPj5emiGxC9fq7fIRWVWvXrZGBX1bRdQZpiJoQHk9yOFFTaZUrzIv7BSirW7Q+
u2lv/jK78qdsY9FLfJK/FRfKP0EGS8/uq4rNFCRQ2tepd5z/98nrN3rH2PdZsHg5Icph29PhPUgg
8NjCpkPEiXGd3oBes+Lyl2sjnxTUXwM4PKNjhmGXQZi2vcNg27hRxAhCOwFF+SAD4s4umg0HOqS8
+Rab5mGF4j1RVPfvqUMEeddIlibOAvJC/0PVYr1450ckxEeUFbs8gh20nAFBLweDUH6G0T3Kwgdg
QcJCCW5Y9qmh0OVHunyTE8PKS3xkxZx3eUCVR75WoXG53dln403gV8ocCnwEw5X74Kc+sM+x/vHN
jR4cGqjJPVZ6Vc87p7AizTdnE3JvVsmu8tgzrFR3ivMT0vfjJRTh0YFIUtP1MsbianaYKrgH6USC
6j8WcZnqAhKX8LJTMswXDMiW3z69fRwiTs2cF1wrFp5qbTEjjxk6oPin8irlLu8t7mg5eddh0VQ0
kDQKceSenXnTt9x8muUKdGv2Jy+Jgy1xos1EodIAEcjP1xo/P4QmyAICKHu0X1PZKTTlodeAO/BC
IcjIfY3ewI6vy6XG0UBQPOQBB6/d35ToMbIPPJAUeA5nbfl3wbSlLh8zf0q3gijZdxpLLVien8H4
9CUDiVyMzSuxuez1LumGRRjxm2Tcpr5C5GBfoiBB3X/RciDH1tl6MO65l0JNBivQu/Zm4yXf1PqQ
mtw2jOjM132YZqCXaM17cW7E0wN9dj8/dVrQPR1wNgE35HpSt+us1TNEsZt2zuEEuX2WtHrr+3Rv
/Eouz0febAtR1PuIpGHjmH392l0xbJ1Le6yB7O4PjmAea8nvwr0gmifMERwlYJ1LP2RJKgAJF9Pv
w8mWiIzUd3soIz0YYVlyNYKL5z142XALE3wHIyPUqMYG/zo7pPmNveTtD2YT0656hmRnTAjUYGP7
OmFyyuarHBb+supJ/Yy8trlrwWyYabOmodcok1uw4uW21qdLEKwMomEC825RvoEbDRMXoWqw5c8v
tnOc9VlLBK3GX4wf8lnVRqb4Tz+ohceK3aPxWe7+fpZMpXSHz2yZUCzIfvQn8zajU7gC9+oNas+O
lx78pjBMB+KWD+V42f5bUuykJ+DdTkESscWj/Kv56X7q5qAXT243qs4zPBqsjfU/SBOhW8O7zdGC
WVzLpyxPn+kpVFXyzRkV6ZoEPX+p2q9Qim9sC4MJvfX+l2c0wJ9S585VByCr1nD+sqNuWVrWx6bS
cCwZgX9F6DUzBuqtWnFiIrvxtA3e2VRmohbRzINgsDq1xNelSP746r3e0MpX38wtbntAygKovYvt
oy8b6R3ejrXE+cKgx8YueGyBIvZYp9e9fnRaHFoEt1uGdYjFWa7fimJQAnl5wVm8LustjtLveIh5
mJj7spEjVirqLQMuOQn5kSKtNNI7GX97yyzEhD1GQ0ezMlKsgGWVWMvMIGLpoM4vKX7Ut2J7iuuV
GY3moWCktKP94HV67tg5xnUrjZe2dbWurCZSC0923gysF5qFQtNl47ygTiYOe3nl6AMKy87sOBWD
oZ1xSV5xaFuRCUOZpalWhHnnOQV7lXmsVmffDdLjStlDhONGOwuICGmQqo6YjjO+pgKwX+cs2Eqw
/65SJbR9FI5qQPx4wUPfEhgoY99rVLwshCPGW3FBKBXnkDyK2dHsvx+LQsu5WkqfrJqzjk6MxCDR
QJWp2xKacDWM1QmyQH6/bAjyB76F1wqw5c3P2Wuu3+w1cfMqb0gn9eqiQmUiCioS0s8wzM7G/l7j
pwWksYBQpc7Cck7S0XJKdsmb8Sd9SqdEIsgNRtHo901QKtFw4m/8u9kmluLKCy1N8QNkiNsDOoQS
A9+z+3LLsLlOdrSg3/kxn1m17U2bxtdts4KTR5UCcNCbJQXoNdAggWspbptQ1DD98N6ClcWWBvq7
1257zoWmPP/rG5RHCJIn1t1FxKXv5prb6IP6RlOYdMO1nCfFPT852tACB7Rj1UydO+UV0zfK7lSe
MBNm5scrIqDNuccb1BXx91+bFoXmG6yEIf6ekqXUpNsy++BtYyTuuGB6BBKJvCFxs/+3CM5yGUfa
VATYrdN+e7mZkC1mNF82e0ag3swzk9dZYTFW3GKOfLXh/KVkC+mGZW/X7zN9n+P+RbgvZGWc+Yfp
HY878zu/K1CMRpk1Dcx+e2Ncy0Fs9K98To62Up0u9r1lovlJrMmgOhzw1TeTPMGZOXxihMwigFgG
UejzLjZlMGE4Jk2xmcFLb3j4hcmytc5A7iFAJ6LtNa45YcsGUzx1wvS2C9LpZ/PQToeIH0FQ9RT+
vGeGFgRf281+TZzDXo2iX76ePgmhSgIDmX2AAWM4agq0ZKMFoUX9g7g2Jeu9eRmILgNnsrZ0viI0
ltPWmWuIUSI+fG5poaIzKW57H49VXNrNZAwPBgHPQmSC/m5dOfAo+bptckr1y7mKv8aXkopoI/Uq
3SRDmyoQKqRoo5qMQyqaMoGSmedLdhqu1sB2b/rzTiyJVePOYWwCj2SYV43gciHKb6H4bMBLN2gb
MFoaPhmaBhqKP4PoRItbIoxvtkWiVhmi4lrkJJTy5xODTW76aZ3RgDrgluQUP8jLyphaRm39xzh1
RvbLZ9IRe5hZYjcyrbl59LMFgwZQ893rMfyJEU2gOFjk4UzBjz16LsznwcWox+m/yssuYwkiprI9
EL7YlEpaQY/QWE9CUI2/eQ1MI4RzWXD4teFv7zWm6xmeowSSke+Gj7Y8Iwa5fL3BueLdJDML8SeV
P+j+usx084iiWCaueATD05JoTj/RJ8tswAK9ZJh5fvtRxfR5iEHDaPCCbN/g4aHn4QQ7xojIn0Me
grJrlGdUSqIwRXoxvSBndyNsBSmpcyEOUn9Vk8dgbPP43EYa6LMkzjOot9Q7bOqm2rI6F0QPKBzp
VxdGR4UxSlL95fakoP5kyAw6zV8JJxiwBLSphOT7z4MNHiCV/eHds8bZNx6DOlUf93VEuUbH93Ee
E27xUF5PZCJ8mZdXtEZ95HiyzY14U5KIdtXZeY/W8UrIieXbQ61mvNTz1aDdkWGhf3SqsOV12eYn
hnsZTYKgk1cuOAMq9Y59nw5gr1OWF9LUwtZTuEb5BrnFHP8rh1q+bNDu5c5K4ZSxgncs0EqtF/qm
RAhdrxZM/BfR8h5/EqgMm4VX27P7ydexTGsLEYc1LEyd8jMbAO6wJKmfuuZ7nXJQU5SFOznsf+2l
Lro0fQ5WOfy8//2HL7UETDQmMnpuhUUJXQki9+ke9xeW7/sif1+V2wBjf8oEUFHO2xc1kUffwEcf
MR5iXtdgFemXq6sCnNUfA4ZSR46GqLpY+6JPgC0SAUmaREIZC0jdFEgQyH9x9f0tc5nqaTOGAgWu
Cf2Jw76igxeAMkFJiyCQgkWv17hTO4EjmUbFSokpgFENdjtT0tGiG0nTcrEHg67Ljy4iJDpo2HrG
oBMHW0FnYeut1NA7CrLTtRpEj01P+Wnf8I8dZoMFH1u14Z0U8eaAGEi33mPDg1pMLLUnVxcyIKtj
IkKkCzWR916S14tTFrdZmOSJNJpU59mzA7zPoJn69ZF10uNuuUYuAgj9bi4LknlR3sqEXbwIn6im
zjQKTVrnCNGwOtfLp73puKLdIveXATVI7TAzIO7y6Cg7ZX+N7TwoPn3i8GVdA6fS9K54P8skPhf3
uC6Q0DArCdAqZo8J7htbWihu7+ytf+V2FTw6uCoruoyIQSlr8mUlX0QbsRSI3LSscibza7pKpqA9
MVhowhl1/fmIJJLOI/7jqH9LOW4CsM3BVqEOS4XH8Z4igBYDzGTfyGU4xZmWIqbyxgL8B3qNG7dm
1jbh3Fo7AfBYcbNh3OUg7wKwqIftrmad016T+b0o5lRrWStYZen2i764iJakg69Mx/G7h8I9FZiH
dU/pwshuyIRVgsPiX+MfOfrQs4ENMHvNgqsNRd7XR/eiYzpun3qO87aw1gXyQWPkSMC1ZspPUwUC
YWec2hwEXL9287shuBrZhiWjXMpROXftZ6ZvWL6x1e6Mye9nUaqB69R9VJYOdZyk2fd0H9kmyUaD
dIQfLVSzoSzU32f8X81ooKxZZG/vosBNX2sm1etS7O7l0aBBYJ2XykIrsjelNL/yzYpp/xir6esD
BckfK5wFvRb+tpsYmBFv88UpGxSmUE6B5WtXSz7rLZRI31roO8W9O28vK/ESQJccOQjRmQfdtcSE
0u75dJmQ+lFih5VeYNixFv1MDw3PiSGHmOsC5jIO/vlLY3KqA9jRE5sqo4Cgl5Fo8dUW6AVpRKfN
VDmkJ2tvzEIOhQKcDzxPSLKk6T0ZPHZ6VGkWNUejxqEqqSWDY4nt3USzg00OMJEEeh6r5IvzTJ3i
Q1LjHJEM/SvjVkT+Qoyjz7iYbe7Vb4E2O6J09O0AHH24sMRZFOAEtJ7uEeI9apAK8CBKQqsxLL2C
iONmlElSUJMJONAwByUyzH7zX0GYHIHS3c+kKTlMLck9LCfm4tMthixIZ7riG2pfGKZJYosEusVj
3PLXmQNdb0eKSizusY2Vby4R1fmsWUTTBL2jR6+NSr+E0hzMW9CrY28B3Z1iRKDM0d5ZV1urojkb
CIxS2jScSOSV0SMiI+oGe7JLxkTlfSPQQdbutjLrEhx0x89wy9/Gv3/lHCvkUcl7WTWTJt43tRaP
3PtPis1EK/4NOkVAoYAewu//Af0dfgnureL3JcP99yrklMyWMCY+PYN8DLbyuTdVhKyAS0vF/UJn
sIz1vGcy+iqw5RsTR/pltKKpjZCB9m3Ebi8VBK0PELZi1q/tGGjXUmwoFpW3e7SHS/njDQGqIBVj
Pk3IRMRna6vmBG0sTMVaiIYJxjMyBFTOd7KBlfuCmF6+5sq8LYhoTYGWh9YBCdGg4cwZf5TbKwq5
J1RNGDtDUGNjQhERdP9rkfxk9BbmEwLffpfaNqWfF2EXi3eQbKA8c9B9fAvn1+t6074QYpNP7oyA
K0mj3c9KJKrhPiqLovEkqvwhpa9isUWHKdXS78oBQCauE93+pOfd7aCxnJ2QYDjanfi6o9yNq+hm
0TPtbswEYsiOqWE6PJIMC9DBVEb7YxiGeZ1uwU9BbH9C3P8hLSsLk/Oo7QX7/eA9C0tLR6Z3aSJe
i+MUA1kEzYV2h6U+WVY/GL9oD50pjm9nfOYCCVmWYnL3jPQo8ecLztprgItyTfinqWtquBOVsYZO
qPv/unBeOkwcrjJ0Vic7WPjxcyXA8bQlx/ia60Uyolenn6r4K0nmCRSfQiUR8wBLDvz/1x+fI364
dqmbHf/gerJP3K8TbSGMwNv856YdwsWXxOOOodyiaXIeFttl5T1D5ETy6wkYX0Ek7t2I18N5if+t
IoW+xkpyhyf0r/QFG1xYhpq9Q6eJ6anGEqt0jV2IkySfCv/if0V+WUVDtG3D5QhZ9jykGqRC4t+R
P3uRYrBBUESjPlKHCU/yAE6ETXRe8FlhSREFqQSRnuiK89RS2I+OeViKX2ik7NfgpMBdMXXFNQ/6
tCsWpmIgvrPg2Dqnfd41+R52lTKgO+vPriUnMfacufMJ0+FyiqQluyWdzmaA17GjjEq0O9neaASW
Ta9GjuxSwdHrfKtfKSr16m3CdBmYJpFdEG1pKzqGSN/CARSEdSLl81VZqJd5r9JBHinEhgA/915Q
14HB8L8QjhS8QNtG3XB2L/qZ/kVbXcc/Zg8PU6ii1iA9LqOAiV1hbtPdMYoFo8ysZKReb7/xLAGM
MKJpj/ZEvWS0wLvWEaPrX1kwF+MAc1Q0ASWzFOOBxqq15gnMvn5UFOdb2EBdo2aWsJ/btLx3rjdP
Ovz47RA0uQFG5v5vLCQXbQY+Ro8Wv2Ex1uZ4g4Y2+DI1wUM5bKJ/K7DMbHq4/AO/4zk7LnXq2xSc
sA0aKDvHPAG7u2xs4Dk3c0Vro02HhG+SxpnOLWAmeEmAdbqd9EUOgySHPldz/NlYKO2OfkUwm/me
dijA3we3D7RvbxStQLPnPr29QA23yrPMcWBFoRA/R3dgbxYHtwQ6S3k2+Uxk8EF2V2GiVMh76FpL
x/2EkM2VmeZBDRk5L636KP+lAzbAREAJdv5ynwQrDyHoxHkijgHJwE/6csNlSSdXi5zjgkP/rWy7
ZKiHqo12lFL2/i1rHVYxyUQY01rpDJyWWzAvjOzN/Pe1aJ2Zt3vZJh1PLqV0qW158PSYNYCqpmmA
j6qDrjISR62rjsabObDsue59tnO+5GLgZtZ86VHzPSwgRWWpPPFBc+FQklVyBQy7A+fQYuo3AA6/
tInaLVbRgbLfp7z+dN49Vfy1ojhRKV5GZ3riLOIu/OcS+c+GfTwCTTt7l7CisfpXumXhn+wtZypL
KL0wLc4bJme5v2o486n92u23rL8NqEHv4Iz8JRuv5IhTQC8QCqCOPUFGFyceMqgIE1hGnLZsui7t
8EQEevhXs5cAykV3GrbStnnrqBdAnlQ//hcE8WcBiJEluXzeNcG+UKtSsStQsHHTrI5jRgdyqiO9
sJwUDL/WrEHRuG1BvdfFa7gyHi90xQzyCJYySs6UvdTXvRTyBZosABScEilCxQX855DKM2l2yR44
4UBp71bWPO0Y3Z2PBxbo1xZ7CgX+hFnsLT8ZzsZ0L1RL/URiBCwmCRhJNLIi4zUmPs9Ge3ka+tZQ
Xnvhh5kl4AfnO6nk2Wg+3mnqnW+Uk+7q/TrrjgNQ7hCKMK9XsS1H/U+kP8vqAocblJJ4WXRdEDGX
dZVxe7Vp252CnF3bA54L8fIzgbkITk1bR/4XEj2ZnWRfebq6mp8BtLSZzV0HPkwjX+SKvwb0xu2H
Y142I3431ER5omWQs12a+j90OTkRz4a1Lsw325P4apucL7Xio8BrflPLbcDmP/VLN8PPvi2CKsuP
lPQZaNgKB38Gb5KNg78B3K8wvTPzRQMpRrfIU5D0eHHvuyS3t2OpGraMfkrcdRS3Z9CgE5PhMeT6
WicQ5vHRg97jvwZQZFJ79p3am4DS7Ue8NgLNOrRwkZW9KCDdNlrxQrZur6wCVmWTTZN6B9QAe4ct
Rel9ejlXNxX1fU30syfHEMG9ls1j+ob69Olf9XGCne90NAUj/IyVQ9FIXYtg6hnwlWtO2FsgbSE7
ABuWdjahg0i/X9tV3IB7whjt2hM17lYIYFpXkjjf87XeZgGQRhgQ3O/Bp8BZri8DGD8Z7KdsHeji
8UtXHtrXGMwtln6My0yKX22HhDd1AA+VV4WkuH407llNeOnfeB+KQi1SUNS/LOhrXjxAqe5vUbsp
rOY4cW50Pn2vstThp95kuEXwNrpGad0cCLKFvhEZnGD3kfZPIwcRyv3BOoc6rsrnyhTAEFpaJ9Fo
YikpvvxI3gDNwxtZWLE+D/bDmtFjvshWhCWyISKfOemM0F3tyRrLIfwU24V/z0FQyn31eylRcjES
SEYINEWAVY7SHZEfCTlewUuA3NnyjO4RsE+EHL866x046lKl0QmLtS7kPMPHpxmzXYv8wW35u2yq
1QASfutWSz90Sa5mQrV0O8wDlbo95uWx34+Xp7zzd+nrcwgvX+KG6nNry7HNDbO6dSE1TJYceFqf
HO36ulxOIXuvMA5wRW/vjE9sih4+11CUT1JOsYNALBLdZ0WnbkDWiaZNzjI9o8NihGKNIRQKZrVl
qTffl6PVDKQq41/IenR7UjdIsT++DF0jN6xrhnjWCE61MYQbvR3j2A4QmH69eedCwAeH+k21Sf63
XRS+CdeBitNGtWXln5rWV3ecQoLGmVtu1djSXXJpPwIwl8ImZhSJWNSdQc9tlDwkCVupp1qXJfGH
LWeXKZd8Np9h8d+tkGaPqDA0iYTe0QT2+n+u0/N+6zKh5UPK6DOVaRxYiBuupZnwq7wmq8Vwjwga
cBgs0O1cld/THwbyo1IczBizIi8Wlb00oTzFaelQHRioV0/F+2yG664fI4WMih/GWWxcnOQ5K98I
Jb5aivGDhNDxW8ypEIB9g9V8qncSuG5/g1MrNsHnWfx8KA81REbpRFGDs6LW5U/oXj1jNDJRit7q
qVVvWzHusNPFc6vZ43R3c/q3SUayjixbhS9ekihwaehcF+iWfcIKfa/lR57dMvV7QHQrCwOxad3d
3/5F+fQEnyiblk0EcODv9zv+IiUhJHSt0jb6mORJDfxAXTPtbc3XMsOYAW/qW9tnow4/KYa28WJj
GiqVUvaDtK8JYTW1PN4LuFVL9Aw2tM4HzWuVtTrYQpRLgAvEAI0oxvMYP+oUYQ/e2al1J1eP3V+s
OgxF0OP8Z2gpL6xiZruRRuNAnOJXMAzIv9ZsBvm7AG3AJ+8YMDcq9nXa4s13Vpj9Ew/pCiXcv1Nu
bCRoy60kmETnKCKA1zkkk9YUxPFW7U1okBS3ujjQ2Q8HCVpKuyJFdAOpa0ps2itcZLuv62LodAmg
Uhofkjk9yg3ziK96XPUuH6nF9Wfd0K585xDs66PEpD2hhh27Dkm0r/bo8n7hSkpNjgwhwkkiXZoy
660OcuObnjKS/vtaqOyzsvesSE6Ved0QhXhtMnrPowM/nnXItoGdq758ePrjNRls3tXcAmsJ2gxi
a6F1tWCVsHM2hrmj/Q+3wEf0t3YpzWOd3moOqiPfWgvR6TARp3e4t4JzBy+yTzRCzpNMyZ2uufMX
b2EKuMJz/AODVE+iPN7DKZt0XztbdqopwhgJjMaPTwy6RRV4UTF2THujNSv4CDDg+cKvSlV/Ts9B
zenj0iDDT12ucVcNghz6A7YK/282VrM3kJtdZSOWAESACBUoKjV2vBZporYSQeWgmmtqrBpXiVNC
rTLUvjPQvgsEfy0V0UxCszIdiDG8RtqEdidK+WbdZcPbEOLT8g6DOj04OyNzVFNpcbrFJ0ItvDuI
a0HJA8ZOB+DVkRlcCoA7Pr/5qNrwYvVkKNOQcIFRgB4XxQNRX9e+qpb4Rs2s88nGqZ2YhmGg3KRu
MDoxn6Vonjsk3Mz86jtMh/LPok+qTXL2LB8MIQylOM+MtjIZpfh5WeGKL/R26RORcaJXTF4scOm5
DBYil6DBp4I3yZ2pLa+ZMh6nAbvvFHEyWU9Bm/ns55wcZNdbaC7BpxY4s5JH45okcAEdM1d/LCz8
60FiXV4YK4JR+iYOLZ6nxizmNyQ1Z2ufjWKqAFcN6zawO01sin3Ks+097mTY8ynGvNmEaeW6mmXc
ZI5Uzw5pYo6YUVrfd7oiEK8FoT2X5nxtj4a0eudY4M59JQLpIhUxR0GVp1ZJqMvaw4UxOFg5wXUe
RUlxKqlcIdqLpjRR+KG/MR37ZEJo+ibvr1GcAIj311YK6ULYGJsUlN6T33rtfPm7nL+FsVHJ/FI4
c7aj949InFBVFuRNbaYnR6Kv7W7d0RLH0n71OMQH2X8O9FtG904BnzonhJ4syyOuicF8K9RMxlXt
JRVImsRYaATYyWStZ9JWtukkh5vET2abxJlpAGW4bhuipixfMGrg8WAzAq8Sp74V6v2nAVlnJ/EF
Gxf1WRE+Mq4zGH5C0kHiArXVU6SJ71ABlZoozMeAZgOB/lWyyFZEi0ZpGSvkKwzT//EWycrFDllY
vESxg7W8e/MWBHfyGTkkO7299npSAeF0P281z6p+4z6fSvTt5VTdnwFTEBehXzsNFdWAbxiMfCuE
4BioV2qLObY5N52GV+4q41bZyUNY9B3YvSayMUxRUuuNerMWphaCtAN4fCdzVv1pHkQ+/wqvJyJg
Fp0sQPWx952yT5tmC3spPK/r+GVED65lv1VaOLZOphNwtS5tyzdqozbILm5JGcbGaO97aYbPfybr
yKghPvcgs0LlxfJsV6r1cONWuTbZtoS+5Xdh+dIJqGBf7sJcAXtBJw+0uwk4Dcx4FHT9T+a7fWx+
sqpWbnqeu+NfwpIgoNrBNBaFJyr6zIRTdLBEfGmXQHmpa/iMHUjFtMk0FIa7A2e+15Opc4tCtdrp
TVVdj4MLMOrYGdhyoo64/ovn7VQiNbsYqF3BHHDkHli28Zb63LDPLwIuCpnUJanIPtKPqw2Rp9Ue
S+X3ph+SRQ3HgAbrRZtz0HpDnlgZ5ioT2m2578w8AptEqBBneqHviaPot1LgvY+yoAQysVvo+xqM
V75TLWqUY/m0Bc8L4odUyg2QclDzqoISN7GuB74Mkz0a4MF3FD0m5YDyuo+OlWGIxpBUwvVRg0NZ
sToo4uQ0+iDUpy9C5+v5kj0ZLb9ICF2VHlUZGbsiVDSvI73F6BcKol2Wy6VN7hk2xweLyB69H+1V
hoeUe8j3G20vp2neR6N99LfKaJyS/bvfw425A+CJT2vA9ug+SjgEUzB0IV/+vZ5xpteuGzFSKczI
XEvBuNef+DnX9khSfkwikgSq1ex/3SnL8AKexsm+xT3Xbzfiajo4kkyp5vKATzTcomd+/f8Ab4Lu
YjKvNJJdeg+rRkNxwRkWNq6Z8dxY7hDRXraVcJg1BTzA+VnBJDcw6VzeqP4av2YIRsmXDJR9zjf4
PJPHcbZMwhWCydFhOHxQquzCtblEzATfhhahQ09R6+2vlUJIIzl4R/SA9R9Ky/DdbTFuY2vcL3w3
IKAZrq4Bn2UAHxoMaJUHj6P292b8epSRa5qKmx8+RlNm3YiXD36+Jl58TqJnTCqGU7VH9c3D5FQ6
irf4ayUGFCaO7PL8V+o8w3+R4iS5tX6P/yHpzqsqYtNnthOPczHTFvw1XcTnJJDlnxwziwIYCiGb
JJ7zKw6VTWzlIHA9c1eleRX81YZ4EpR55763pi800UviPyPJWEJb0cWT7Nd1dTBqQMGMuduDvGdG
DYP06fe4Gh3s04vfNV+Rre2ULsi3547hRe5cmw/ERlBuGVfxIg7/10P0qei5QHWokQOFW/GJ1nFw
hW4lYjGQAlqvHPH5Yc51xGVQHFkYjOqnRtR9UhdhMUXKGcC73EX4+gcqM3LQUvcK/3WkdeeWKXPI
Se0Vr1HqbTFeZNkTftED8zUKd1LE1EbeVkIuKDPQ2RE8MLBSx3LxvcTItP7LIUD39G41EWTiTpK1
wuKzwqGZqE1VBMLtKJ9mZa5SYaTLI1TRibaIti1vVVEN1aH3qjS2pvvjUyoHJ7KpcSQyWYHtJa3O
w9oX1wrOV/ux/aT3VfPlZtGobkeSwfdlgXBSoiIjBCq4zdPtkPztL0VpksyW5mHHVv+9d1nc5l4q
d/0CjGfStk6QnVvvQo+fjFNlcCDkcApmQb0ZNovdpMpyLqGKpoBjSaCp72pC0Jj+DO3ZBOHUyyqs
RyW9LcD4Uh70gTnNjdqKRopaiO7tkJuImq+a0aZsreuAcIzp3be9mI6RTg+/0vf6+1IMHO4ZVhVZ
XBTQjR6qnaxDX8h6yMwJcqDJr/aTveE1+bU8l7GpAlhpFWE99w7rrJSCVau7c4qiXGr2MReKi/o/
teOIq+h4ecyXdqJn5Q2+FrmBcAku1Q32ccr+GaDj4ALA7YzeVK7tf7R3akiMff2erABR+pZUgrcA
pXKwrEpH0RtblOk8lcLj8QcoZjC7Nyq/uxgeQvyjzgw12mIeHe2f8l4Gvrd3fTNgEj1IiF58ctWR
rSZfx6rMAdc19yS/bt99JppBPdtf7ed4qoqRXi1RIXavYEaNXmeF44RDyeyS91+/7z2QYTpHC10z
p+TgzVpYe7DqyoSFFQwhIK53G2+J4bHS5CH9LBVUQVE00Ok4bpmj2D+EmQE4lrL2ZCOttXsQf84o
0QYmJAGHGGJNsuAskSDctFoKCqCCxHjEFPjTnsRbv55TaWeY33CDaSjiRx7Jhelce4pTK/K7YdFQ
7+74l9iM+TO3ddQXNT1pWqzQ7z6x0eH6TQhDhH1BuEPtjImUU3U7wm+jT6Y3uctigzqhxIrn1NgU
YmRnPNXHPWIrgUT4nrJUpyrXIhix3C0xF5z7ZU5YJQfDTePDlQnvUcWwdLQ/jEdlZe+cSfVKpW0X
RKIJWnbh0nmkezo0pgvlVc9mCxTryNsxmuaq05fVE8V0E0b+ml2MOeAkVQTNHHkDjlPuKCpLFAah
RYSeQyqrzdougFF0fBPXMC5UvYFs+6AvsHm9SQDiMT2ZOo5veTt8vdotgZUpwWBAolq/W3Eq94eU
lk2GlHw3r/ub8Zwn+2YEVKjfMpI8/xMjfASBgJ4NfMaz6nR9Hn0deukjw8L0t3GmbX4WM9qTbhip
m1wiJg+J/sBc+M5oNWrgnMkILWnwRp/kZbBFgpXNm06K9Xd1SD4VULrqxz4EnTqY9w/FeBlHhU9P
cYlwBtDYLwPwlzQdiIBkiHpcNKH3o5VOeXJktSRAoPKb205ZpN/icphh92F2sxohkBv4P/LxVU7u
uN1LqmSOvhyuvkSOhtvIMXk8v+To8Wyb7GmIoUT/cI5SmQ3IY8mQJuGWxMaP+xFhwjC9zCsG2GUi
7na+Cr7RyCm7ytT49DY/cBORYNxGGlzOde8VdPBg3qb66VCEOdftBs2cOVuICqprtheEP7dPzu6H
TolgE0pfEj15xhTYQUkiSPpL5RASFmGXuXZPADIM3fmosWzjIaaizHGfLc/X8ax8uDHZM0T4Fqxu
AsOREcvPupTDcppFL7TkH1I5FfWGLoZKQiAJYTeXxHaX0q95cfqzsQxcWiRpLBNgBIYbzWR3c4eU
ZH9mhh+JGocxLi+AcKXC8kqDX5+lDYXO3Ov4nKwVMSKWl7yqXUWWm1w9vFAyls29cbCCKiZtp3yJ
uC3sC9+1A0m+qLPKCSqeDDE85qX6DwNw+mJfWN1wUL7SnH5AjgcPVXt2dlC76BbypBCcSHZyBLuH
R0dIdERrtqBDWmeZxb1XmjbsKQU8JSr0ep8eOYZMoylY35+/5WfuQyD8ENE5JZiZw2mw3W+lU8Al
k/bPDdQtOwm/BKT4KiCMeTl7MDa2X3gj52H0enslnx3k5IyMQ+4rSuF75QX5DG+T4vmcgbS90gMp
HAVgvwvkCwu9b1VC+vbyaE/QwXTJmjDidxk5KIaIJVsT7pFhEvyBZMvCh9jWZUDoyJUwK9JPvfR4
97nmseRr1fSJH/4E2eCU/m0Ny9TiZntB9S+J9BoR5x0eQSGIwitlpfzK9dSzaOERX2YTgp8J7WZB
JRCHe2T9+3oBGDe12r6+urJ+CF1EnrM0FXF72nGL9s7SsBNgTH1xKVTcNH5beECX5Kf620rxyESF
O8Im1wUZSNqp8rOsM88pOFiUPxKKBnRIXx9ghXyZr+rkip+VOKwj8u5DKvELtA+bxx7vZiQmoX4r
pLq/HyfVXS7CMI8Au1a80DtS25DVlT+NLUVFJe9ZBWdi+UR4ltJeSY1lCFVHn4rKuojjKa9MbKHl
mcCn+Igm4nHrRUOkPxetEcZOJExaMUiSrC3dM3Bb/g+ewXGd0/AJvi+SQOPW+91H7Mi65v/LBy2k
XtL590jnJe4cUTbVjG7tqPGhuPEKnvij4xngHgHcGNfdSDCb6gstsvThaC//zAbAdmDlzo1AwuAV
3zonjTNPm+zSIhtQPi4fbwUJkrtbNmaQ9bzwaNc8WoL+I4sLQv1y/28T9NfU2vSTGqqaX3vOtnoQ
E7fHaP8oYgBUj7Jio4RQilICEaenoGyHCXujcCPC6DNCGdPHMRR9dfULBqVuogsPfLPo0tdgqtS/
YMmtaJcR4ovQ3m8J2pjg5+qhjftTMLJY+wicDo0Qr1r6YqoNY4YN3PX7fun/ZhnIgZ8BhEKkZLSK
Fb5v8ooEBWpQRIntABYtwyIz7zTSCtc9GkOn8nIQ4kTztH29wdlSIVj3WGMTGaU/LyzhhV/jrUwl
uYnYRD4hJzUbAfPIcqty83esRarsLeW8ON5LBWT1N8COT44P09U6UL4GnzWspZGyddgdZeQoleeq
jLKNg0zbv92wHBn0BgGghZtq9BQ5QN10f/dqha8YdIVNv/0ZV2avhisnlcWMAGUNB9NNrTXsj3/T
Z73l0c7I5PMVHwQ8rl6Dj+ZqLi0/e5R2yYozHqYm8gsjuMK+RPnA2vMZKehNd60euGgKGV4IJ68z
zws4Pt9HWf+N+W7E4z02AF/JbGK/EUHZm9mK4pWMxM6rvHJ2umoqoRnCWJ4spZh5MzntKJ9AWVyg
mEeEdRsXUPbfoytpSAUhcbUsgQQwLvX8idwGLN9baRk936RvWFjbuQrvWBf28PESPMB/zGRLmQlV
U9ZbQIndjnyfWToWx+3qXUxGBw+J57AacT0AvDoBouTJGH9stz7t2rpVzq9oul/bGTAIIUY8spgi
NVtAZlWgp024MuxsVpq9Lcjbea7a9LIjHAkRVB0mPZbkdiU9+PvBcPkEdfvLbdzbGRhCD5lHv3Ab
Phz/TXAZjzRBpLKYp2EHOgwRgw74xSeA3Qp0qZSwpWMeiH+4aLu53kiwqgC2mzupAHOZyFvbqTFq
5oy23giXpCUcaabRF7tzTQqaBEJwLF9n2H4z1fmWuqFJZcZxLsqeF9oW4viOUYXPI4Vxm4mvm3f+
FCjtBfEZeQoQ2KEZhzxlg4kB2uHYbo1ltMV9Ze25uGmeAUTtgjrA6j7fA/mAh4nYHC++sa1RK0v9
1CTQIBlMq9by2zDosFTHV9CXcBhTf3JMVDbhtz1r3t2LJ+pQlqprOQ1RfNxEUt0K36XHVEvqJQKP
azzcMAZSHkRvRzH3zjmqvoRa+P4tE9UklN3rBqDMq/Z3wgkQz+v+pxmbMOnfme/hRkXuGGSK5bgs
i5Dr20YoZ+ckQkqdFcp+U3yAG6X1yZHbEb9mf/Lw0Dopis+l3GCOb8qzXUGKnf3Xu0OnR0B1zopK
p5czUWHUhGF4BAr8tMljnBE27/x/kcdF13P02rtUyDXxPseLRJ8S84N7FNH2nmVTOnqfpBQRe6Vk
s5EGrmQ29EASvPqbX0GEWQkkJWTYgGiORiH9yz6qSNW0EJ85Sj+IJYerZpZLgueX4YxXE+op8qIH
Q6DWhVV2Ap9nAovSmnMA34dPjo82MfsT/VRruAYT42Q74E2UcpazSzfsD5pvSoMNErxQmen0c4ec
m9AyJ0E7kEcKpVei/zUI8ABJ/ufrHjgE2fMRyv9kDuIwL+lgEtrWNcmco5w31kJ+irMaXpVoWADu
lqHOiUaj9iRde+0SKb1pegU1d6gWZfaHiI1YewvXI/dPuUYrD70Cpod/0Rw8xjO2EbuAr5SfLOXM
2OJowtxKhOg+1smez7dP5bMW1nNEieWqBRP41SRWGu35pJaq1XAsm64ZRwLaZtqWjQeUsr82mIjA
tI7GjYBh6dsZiCrm+MItp4YPj99IcMfyP0N/mta3STTcjwkJNj3Te5W9Pzl5VEL3tDGTf+d4sn39
YZE6GdEjDWQBycMa8+FCuANSpgXeQl+Ss5FpsRIjfeHM4+hEsGxehAfIP3QYexdB4rSAwMIBiO4G
Js3hZtLqI4wN8Jnx3Ng6lx4YjYsX1p/lrGrkAyj4Vt5EX8naFZoguRHk5gcj7yX8wkEwokoPlnNX
jANhajMwuymb1ogq8G5eGTWCNuAOhwbqhEPOiF09w5H8MQT9T+Rf3rlQ6z0oR/72ffSaaEri2QqI
rT5suwqGhydXlAC+F0h7RVjbfFIXQtUpjVAHrYfUB+cH3FSTqnpLvtibG2l3I5jkfigMmWpvU07R
rWEPalsO15Ofph5tnXgcbIbrzmMh2Z9l7rCJzmqjEbncLUEVMan/Z9ECG/tXKPBFWG4/gRS70HRh
Z/PI2WAOxWduEjSOCWF3NDtq5SP67WfTyt/7OhLhgcopJhjfvp93kHy3GkE+3QNLVFPp/ezuRqk6
H9y/JZrx9Sem959TPQtqMkk8UK30SBSoNzztHOMf1nSvBykEOWJjsTtSKd8WNYrMyPZZHMpmKp/8
MChSHXittCBSQzWxH6Y15fVosjVEKd7HtSEb+87e7WgFVZISafCMKh/6rffIDq3mpLDIDYRebw0z
Xs1k0ennBmhXu3lv8B5m5iBg0XPKwTGilDHGj0QRjgHZmm/p6EnRGkCgwe9Ph4cX3kkr5aXuDbwL
Y34VV2Ay07izDwyChZBEuXFDqD6GiCWhPgW0WpKoS37M+8zVSzPUzn0AQULSqQOSMJjvblTurXqc
Bf+Y5CfR/zgb4iGSmSDdShPJfz2SIJ/AbjcslgZo0UVw0R/mhhvbeEdxgFymZDf7VPPYUSklXjv1
smzMxC2BHWOFncd59xRkOekNvqFJKZ5EFGQ0G5pljQFV8gGnpEA26DqPU7FHzIOoqP4qCt6/+jKV
I4lXo/+u4bpEQ2S7kEc6Y5icMJk9m/Z2Pq4OCQLpP3tQuDPQTrfifALo9YZ0kGVx2m2V1M9TE6ET
aoqA0uL2V6bJAvtWoYXmeoyWI9SRg+NN5VXC0hQnEb/1ZO6kYcmdAuSLygmK2eGjPvqHg7wqMOUH
a4gtHwueDEFvTqqVEgN8Q0/nlfoyYGxUT4sg0yN0MMBqHP68PFIQ+aelnmtQn7+wk5yO2MjoxIaK
mJ5Ey8v8uiPeHTlMtha2ydsGf4RLAPm8L2M8Sgt422y4Iz2P4AZyjWZlVhfyg62G5/3kZUkH7V6p
m7tdpzV1vhs3prKj3rElxE3qTBoBeObdNwqTka4nB3Xvc07QghB4Ue70M+SBZzeQH6uBh0Dsk8To
bfWI1BBMFK8pJ2fxR96TDnLFM8aN05h4LOD2Quhk4LnBqWtir5rLrmNWEoM6fxd298hfwX4PCq5G
lF+PKlJ3OHtAWMKCzdM9inH1WPSICYG5x0060kQvAePyfjb/Z/sn54TDF8qEKjgfhlmbcIKi10R4
eBEGXfagiiqoTEwIqjaL6U2JWmwyk4vtSGF0daq4bj3VvpOW9jGyrxqHhaaCi81me0dDbfgNHLw9
hzzuhDRKUi/CSAUy3lp1wcJpbyxL3WKqxkhuimtgcTg/+5xor9jSscxajWATgNH+tZ7GIiuSijui
U/jzYbZloVfXSTGTPhu6H64E0O/tSPTd1agDR12AqHdw4GNelqyGQYyUn+bEPluDk05k/I4NDcCi
cl4nAsSGBEDO5GhUuqQXjlcx1TzNtSYXYPPcyN9KD7pTjCjra2ChKdxExmYspDnbq2tgjL67s4Tn
yrYh8qbbwYrDYasQfoccZorXT4rB6JfY+nv56t4C0X7XH2HswKdHrT90Z5sDJNoiXgtVpyYdLhy6
68albxqKCxRypGXhULjCNtuVSSynQWcYvhfqiW0/LZbFb4l8zemO90yuRRn85umiL6QeV3whJ/SE
qRe3+hxtmdzf1Y0nC9vWqJxbxopBfMr/Io+anSio6nF07vYF9PfqAqYTeF41n5uiArHTk9K3gGCG
ME9VjKhfF8QjNth/QHFMuj6jro+vzZQ8m9JqJvzuDDET5X9wJkL12wSeh6bMV0x0rjM4ODbfM0sL
Xlb1fFEOYhBPvFFKYxz22iGRxO3n9/LjjSAmKOjFLw6Uf2bdNTiPZPrOqWVH9wpbBnD53E4FdE66
5/DJB1FYoY/ajAq6s9D0NB0QgjA7pS4E/mG6T20H00KPDbLwZmelHb2bbq6GQ8YsYfBI+2JuqOPY
0aujazL31JWNtaLiv0Cta2QFcYNF+1CBy+viP7l0/dXtbBC1HeKD1n+P1BpkHcC4T5yQ10FfRGDw
Btui6wGD9E44z5FF7ibe4wMexBSf1Ukc8wxNczodaNZIk6S3wRy6JkzYghsRziZWWAsbfXA51Bzj
MWCufvAv5wGW3aqTjUavGAWv/L6Z5cVRQVtvoL3Gtf2d9xCR6SXiLvXvDzVql+eOYHyHOdu4qT7z
eEEXuNgrZqUOkcVUOp1KppMnYvl+CvVZqmBpW770idEvcFEAB4ugZ6Rm5445d3qhD3oUCcbfce85
pQzS+t9/tRM/8pQ/HoO3/ajfSEvMXZ94rdFRZNtZAkhvN3ZAgoEJ3ypbMiifBY1opjiWvcplG4uu
USo4WjbI2iUglYdlX+QjyJfFNiQUIBTTno6Oiezm0RxlJjI2YtdYfiYZ5kNb0+wH58shJEB0fGk7
s20bAy2hb3U93L9Zrx6FriWzr2HeimBxzm8bm+Tb6bwJ+zcRW4N9SFhE4kb9HKBp4VfxPVafjJ3C
n97Out7pqGynRFkROPl0RZviRvPhYAghsq4JLC6EhinGEJAq0INGMr5AR9tgPlExNoxxg6FIj/J9
I8c7nIGzRA3K9yd6l0Wz7YZ4FY9pKUWJ52ab39wJpumqIdh/6l9ksD/64mOJKui1jKEq3ev0gKFB
2RTBmKo0N/AVhMKSld+Otz368sbarRwfzvIc1/vrTEv6i+o1SP0nZJbnVljnEkaPSVrEjENX+k2O
gz5yZqtFuOfw7tjKp4XGLe+PyNkyq7tTnxK+8fqJ4X0Uz+AZjGk8HTjqke85BM0VRsKG0GsCNBBd
J5JTYIT1FV6LDeHN3T4KowKBTjZFOv1dbZO6QAUDSyX253iAJDyxdxJsgbCifmBHzZlaYBYJppvY
8c+8nYxwW5zq8GMO49pkVaXKkop++gfLVnZ1T0vRFeuLJKHxhs8rWOvcSUjYlVbkLMPG4+6D8CYZ
j5EmkXwh/CpU41Wf6PCAUwBKCbiMIsAVvzuOjINnebiXVCHHD5/5ure/6V3IugpTFzvLMkw1ARlv
bwp4B/3MPGU8JGGbVv0diZUhOle9Bi8uc/UZHQWeqsoXeBwfG0onhurAknzZPoR7PDn4qtHYwgKP
odAiJh4NnLsjDab61dbdXOxHVuFqXnMDdUZ9BMjB7Xk0JBjPBs7o3EFOlDb/QjCKYaRjcJOkqEav
F9JfAoyvpWCWhHnXPgKB69462nTkunFqkNszuuiJ63RCXYUISwKJSl03awzlNjO/hxwp7QK7kEQ5
OIlJb3WjKmDBckJqWdt0UgxWJANh2BMSjog9VRlvQjZD3H8lEysyWZdXs/YGboFLIDw9XorPJktt
3oxCwFegDB0odGvFM1C6iBvcX5TtAgE9iPUANlZ2l56NoaHzSKH7DMLFCKRRdbEW/fyZ7LVQrFiI
84KbkBSHdzbik7i7l0wy+OnrgeC1xI02qphxYmVyoPwRCXteVqDqujIrtYwClyaZ4Kvo3QSdm4vr
awzKEB5L1TvJfeIZIVlOEjtHdQ1CAZc37fNON5LOLv6DUhVVfsiXZDfEle7lOpZNMgO674AlUaXx
r0FQfvBEGtaf/CW58KYZla1lnAXzvXsLPyBBvXAxHhutlqXC1CsAvlRNic6Y/CsbIsHx2EmUFmbg
Se8uPNMkBUP9dPJv9Hn+wptvy/gLjGbp0qI71J+vq+Sm8ZoFHFJSS7zFCqZxm2h0aIUFCsE5arrE
D7ZbqTpKQAaIags79o5ZwZKHH3c0uDWjhMJoglwTQs88oQe8o8cCnO0nFxLXTjNBZF0dG991Fr+e
8bOUIMIFz6On3T5IbH9/JhWnhnF93J3kfKPVvKUabvXJv7uFfFkiNFjI+/n+US0LYrjtpN8pPXzz
ducnN4/4aZefYe42exn1AUSp1nsvRnSb8Q9HRQ1KxGkYSXBEiKxG64XTX5b4RzGfkAercZ3vF2Lf
TDLgbie4lQuPtj3G/6LsQ9c1+JHSWicZ8C6QjYLJ1YVdueq5CgWIjqUGVJWH8tnIrykqSFn3vYRf
RdeL1ip0fGFarziIIs0uw8muf0zNRZQ6eQemUbrVjQ5DqxPngP60USqwDbNnm5XCbaaBPSgVN/fV
RLC7b7I2qyjl13QG9DZuUXT6/rG8rDD0A3lJeMgstHYSANBLvS0dFhV3TADADM8Wn90esSw6oFaJ
Ap8LjK/EyLIoglqbxooQHjkdj6/9HOsilyo8/oBYzJxOxjYPW3oEbK3cyzul0OqFV7N4CJleLswx
Uq7VbwTrJ/b69fBWpleSiAGUo4bZFeizas8Y08767P8ibk40Q4njQpgfdwYteaow5tOUEH47KpcM
R8W871YhsAMvdtof7s7p3TCURzyssXKBO5S9qb737b/vv5rn8ymaoW58C1U6lbEVaAVP/LoKw+T8
8c7Cpv9vaQxfu8JQ5y0FHD4MZJztNw9wwRZJ7VAGoGxt70RLld4Gighc8PlEy/eIKvY9qBRK1PyU
U28v97U0ccPbylcKr78rVMy2V5gvYGDCq3NokDkzCIEyKwnNbaDrYee0UpRTgFMsMqiltdJge7ee
iHraD4hzUbRn1YAQZGQcGx2gG3DIUoEMD/q6v8lw/ziGLmeLxYyb00Vf0HbxJhRmNinQv7QCrmd/
yBv3hyQUtQVZxnHLDPBImmPnEeSW1s9nJav7q1rheUYU3u+kI9/LUAzpS4ICAjCFMypfkmvE4iUI
dwemC0V4TvS0br9v79pqFcZkCA7LEPiccA2xanCDuD8fSzqOSkmQkcHvymDyUiRychiltV4KcSEo
f7VWg86YNdb5TUwJWFl4z/hO9Ebjzs0LRPJaQ0EEeNuMR4p2cwVAKQJElkpE7h17RDOwCLdZswLt
Flrs4Mi6HtbMqQsaPFsFmTNc0/YUAeOMemobFHhsMxCFkS2hd33WLFU0zW/VuLavVYrUPq8MjqFV
WQop/Sgd4Qmib/IOKxmAR+8dqcolDrp/MRE6numsnij/57JcQJUk9/zkBN4S2XMCE/fxrlw5uZ9Q
+EJm1M15giryE8r/z7fPx7WRs9mdGRRJS+Lxvc0f66898m74rUlIqXT/v0ttDVadW8utTWJkPWuF
jUYyKCtk5QnA5Q+PfDvff2iMfug0FHP+/L4CbXdT+tTlb/w0WP8J4K0zJ7JETocNyghRpTbDRB3q
vyS9RWF6iJ2WKTzFSBZAE40N6gJQnwhpk7eUvEKiJJoDkN2rtTBDVODOAB/xHstTPsEMKpwhWHXa
qVWw9kZdGj+aJD9BE2+/lsTABqDR6OkD8723ZRX7ftIPtikQ/3/MMJtfZG3i73f1W7GMxaTH51CN
xTxrw31yKt9hhghLBuwZNmcy6AWOcaDnNYAfu2eTFu+6uC0cflVv+hoQth6ibINWmaqvD+hhjKqW
dS3mQj0FZukBYFYJkoIcE2l/vbRML2H2RvwCEp1eSqPJL+zGXR+Fnkiiok+NHQGypn8oSawcEo9W
cMAiz4w/AI7dadAcQOY+h3SGAoGylUP6RT8VeiaAGEdUwpZ0omu6Z1AtbESTaDNsBvadnu433OcU
i6yx4OKlCUxQVN5Rlq4URsMEJtEck1oH5VhRfOHk5AP095Q3jS5mJWRz7xDnFyGtBnixQTmyEODu
1sw9OM/pi/vCECSK+f7eSozwoPOahqxgJz+UePt7GPYebIbWbV2YJyzEvQnKmqbfP3hYLAk/zcUq
A7xF7zoxUWuvkI0TaazpNiO+C+QD4KGyaHzz9KPDbKQkTyRp8KiuT/dVcDJWydIASQ6RSNy9uyhW
t+qt8DQThLg5GS4KiWgwQaw1fsNS2H80W7ikdx93fIy50YnQ+e145ScFD235A9oLGqSUUZViSUfr
KNo6e9Kl+gkJFpf5QIiQY+qIivEXD8EGl4YGH1o37PxdntBuljoXlm+1hiiqEMLB/2rkina+Dion
GLR9/Uv3EppVLrMzbDNUp3YyXQrJXuThgvoq/DYaAQM4hcoxUYpdhlExaVWUZGFMQAXXcYYvTCcG
SCWFRVcXFNZxPodK7H/jtYHImpsJgkNEyt/Hxex/UNXCGNmtCvSWJTfaiUyAiLtGLG3dRToqKbf0
A+5euA4yeRJBNC5ZCdacAZJdu9gQMkynXkM/Wz3RBxGqezIIlW8NwNP50Cy0aCGhW0WW6pwmEDyZ
NuwOeN7Pn57ORxiO/a1+bkRue99F6PJXVTNS+hFYxRsBSnkwcHdsIBjeH2Nyj5OMoS0pfEP5x4Ey
c/j5sxvLynFoGL3wSJBevNPLVHVRog1Xrg4v1r36Zt6YfGatQVXbSduGm1Yjorqpxpgb+pTSEaQW
+/Z9qiH9RtN6L9ozbI4MW9UbOisSxmTMUXqchohp6Fz6VowhdqnxzKUBfj0sCZWlSFupHHQ6tHAA
Az9I565oAYlbdwPrLsRQMiGAssMOQ24eZcpruFGMAjgcA5z7CQNYMEnJr3Cbu0ZualtQ4EUA5CBS
IPdo5gtbnz4zSj+G6vvwajyBgog5RpcZWJgnqMoXPgAwU5mKKE69y6lEsiHNFwwjWJHWFAmE9BHq
V0tlUEZzB1Azyam7KiyshhAu8zutCIxYQbv+zy7SgtXzsSRXz7pcAsDI2wJXbRWzlFt7KExZNajS
1WGgVqYDh/nvahsxrw8OdEMxVZPDiAzHA7fkVk/Fq0pSZlm0IChiyWoaiCd0zR3gtvC2KSrENE5n
gtSaTlmuFuzgzOnfLi9bd6QxnjQowzqptA27L6poxIhL3ww1zl1KNdIIPSCc5/T/ywIZM9IQWiTK
BIUxIOVJA5KOPoAQLpXz83B5W/CCdm7Sk/LLIWYUwHtcxQcjGOqQqp2RBEX8ZuIRBQbSppPcMe4J
2L8k2wC16e5WW5W2dnErNBdmrbcQTwapD+DeOG5XHax+Af/qw17wkFPwwmSIVhft57ZxOKnAZE1v
c0ACuJOCL3JMSHqK8MjiRnOhS9w2+sY73kklsPHxHtRjjozsdLHr50+ilTPy4GxGV+Trv9AHXj5J
f3h8+nRwLRnv0prNTvCu7cWVZVr9xlWRSIdQ4Fm+G79dl81BHXLIV/Yoo1fjHXAcoYgyt4XIBBzq
M+xvBe4Bc+2qvLUUZz91jq5Yj5mkkH1ox2jR63VIGhrlyCY95q8uZNi1zw4/o92/kyQXzK3v+gdl
0RrfzEKqjUxvlOAB18EbYSoLiboKxxJAGmqHH3DOHAloUu9c0H3f8knSNwBrR98AvuUngxDl5C/n
zhCT9IUfopRieiG9K5AxK21mQHuPTS4ax3WjsASgAMFTTV33SUpkUFXC7795uQsLl9bjeL9LeZwx
LEHvEfBlZ7fZ6EYHH87fM+42z7Vivs7LUXaA75dehIpflF+Mn8o8GBogwJaD21zdUqZjhPwozyVq
ieLtCUjuifPBRfZhmqemeDpwceGz5K3hhXxnjwNksDL5KhkrkSjJ0GHzwBoQ4Y5DHr3/nUPjE2VM
mjl8/W7JU0GuLVFmETZNz0iYZWG5E33viuWBteApXlLTkOBJsG9QYfjOXuqCpO/Fhh2cL5lIFQcg
kna7698IED4tnJoDrXMXdlhPkVUB2crzLMX1wlPWPQfFnteQeMRyqfKWsk178aR34R/ulVuif3VG
JPCd1HJU8EKB9ptcHyQW7tH44hTU6vNob6y1ctnU62jsD9fJi2v5qJ4mf9sJedYzKKSmapcC7p/1
x9jVIDiJeyi2Q/Wg6c1cls+wWX1wAwIro5HZRcrWsg2mGGx+1NNqSevGGUlEx8eP5L+d9ekTZ8r/
sO9p/dGkvz0MLdFsmmOjxsKTDZ+6GO24Ouy87fo7JGl08gjBfIBFIH9emiJE5RQm+GtlidL71a6K
TdVx3nwpanYXgzkp/+5fvzTvZGpiHayqi2MOKDg13a1PUlUMWmlPqidUxSRYqkglo1Q36k3zZir7
E7V0inM7bw7OGYXoXALYYis3cm1ZMgeJjHR3LYD6iaP3EvE58OBhrtLygEgBgwskexxS4M++ZErz
+p5xUqZUUncR1eBFmDcaVPqNBo63bGSTueEYYU2zN1BuphlBNC9xTmkL2nReHm6UtvaIexzZ/tRy
ifqIPOmbKCnpJZ0u2ZVTdNAvSWJ/mMum2CuZumlIY2uW8xSajXGSz4lQZ9gAcptKW3c+JaDHhLBT
2Zvzr63Wi+5XYY6VG9DzKDD1qOVDS1/dCCx58lfNB6xWMcCVutrqf72zfFh1H88fZvGDhR2JD2wQ
vMkMB8qAGtpMIIp4qeRa4rGj7jBTGFGCbRQbopBdvrCAgVTGWSan4P3hTktqHzS8QLz2Rq/Suu1l
RgYzxvIQ1j9N4XVM82jmskfHIEjOQcvs/JGxYUwwSr59t/nMgHtCgskjBktNMnsKabX1Goc/8PmZ
pkmIRlxt5+JoUcAOzokUEAZUjsPY1iUcBkXGocNjKfhLEdYqsJJjqaGx9fi3nJruhqR8Ice3QE8C
q4p7Tlt7YnfSZHUzaX5fb45xedysWnnu1eZCkAfiho07D1K5g+0wAAClmZB+PYErScJ/qP7FFKA5
k6OEIo+mUCZUQrASbhvfzOo5q5VH8Ow5V/QZDl9EZamjl2gNukOxh1JCTaur2KPMIC+Ig2HhGT6L
J2ihDIrtjY9vT15nK6Vo/nsfnNBZt/XSiXjFqPIQ1s8+pYIPLGpQjKkMQ5XR0bwW4Cm/fjZdz2S2
T8iKSwjhUMSKjVW7wTp35JP4szSmljfHmKqta70roJUrt7o0LOBJL4SFfObLSDIbRegDakyuQrLS
Cu8fp3nNt+LI85HQN/AaTrjzo1eTLbgvRYGrYUM0KOsvBX9vRqaKXjE+7UmgYjwkxnwj2F474m4d
O0diAc1y4ssZ4iPyel6AY+kiXZBAM/NZL8b4wn8fAJM4nejk1kuaX4ZwxogcSGnG4sMDx/lawzwd
v5Cpdh/Tv2JegoNIFkUGwNYncpzyM56OQzTLTLyunc0DTmBQ2yGUKs4gZtW5u3SwD4b/qc8FpM+m
V7NwgjGJxxBZ1+XV3mTYb5hWmOsLmA4qtYOJIWsjo/0F/QWCHXDaXyLjdFD4bNywhvCAkGl64oCi
cpASf63Us73wjG5j5hDbGFO1sTebve3J6EHE4iE1ZpnBNYiBAkCp8HmxqnlPWZFt5vTENx/3WpdO
dO1RVNXD8IR9oAHowzv9h/0L69jBenm/CnWigkah3crKE0AXLHHQ5XTyBBj57+jVNfhIxEkbIGdE
UZrxFwawHOwJUoOqn7j6KiySHSNCN2rq4KvM1LqWLWgeqg/0roVIX2rZb/4pLCpz7vxVWZ+hxMG3
JK6TdbApIdyOWqIDGL75f+ACh4g5n9hVe8q3c+0RXYP1eXIomzr22g7muCOqn2S7zYQt623ZGh/k
1TnNeVsmBv5ThoYiXsdbtlIW/59aXR7lDxCSTV+7dO1WgnZdwgr5y7zckQtxF/fdXPuHHpIH8q7I
uaIjgW61V4Di7c17dWlwmg1FMNx7wl4eKUJRZ+0LQpSaV7wK9pBl3eDluIECvnpcllHrYApUQW1o
fPC8j6EDbUMax3kFJS8SgFiBWBNue5kzyPD7O2nwtwhCiXgMWG72ISZx+dCS7sQlbfVLXFcgHWZP
VwM79G5lM6lIvSEX+5AiulE73kfsj/0VRbp5lQ1ykYiCUw5o/9tQC0fVawAseeOaCXwcA9bNvYvT
IWPFEOrot65VMfxFj9Z6wfy0JVtg1JqchcWlSSq93yO+fLW9rF/k7Hl7fUWKKuNUBaxA0qH8TkbU
Tj8V7H55RzeHQikWrjE2YdZQgxUKg+tjDTnwyh82S6CQqwdYFOS+ezfeT6prYHWFNszZnFh2q1bO
8uf9f2/38km+njQvn3wzWD/4DWBYOthRSRHgrBTJ8TRwev5qPYDYIj92jCYjmY30Auo1TaJ/aagx
Dd6IvvlWKqtV6nugQlb9/C1hE/WXiNDAncQZF7kVZLgvPm+NGAvPIkkhSW1wxb0m6+yjwz9whKej
yvcrXG3DwhYNtdLOHzqb02Vi3/o3YiS6PKZJ0FNtYhR/imogZbEEOzEVwM+wK/7YcXR8kMmxXJYn
cD5HYUapoHHsKLs4tVYwxocTfyUm29iY1OjlblschIEGEFDgMLLLDeKbX8oVgpW4hHBXVlWUOz4z
UivLcKKtbWChF6R/bt9YWaRjzeVZA2wm95mZV9Mf+Qf663JMoJ3wk1dHh/R3DicqBBJ6UzeY+0u9
wXgk2qKqsocq1gcDiYcVGCEQji/Tg6LoSIdNXYSCooc1CZh2jSvTZTpPqKLa6NqRLR7bDanm0TPv
MFSz6GeaBD0BQxKd9mFuEXLjMnWX0MJB76X+FgblsfKKd9OuUEitSgtsFvCBtm510wlXhMuO63VE
bQG0FLgDQrC+R9DMuAogCUdjCJquVDwJk/ZPzK1nFJtxk/EpZt+N1+QyiN8zRCPCiTAvctHRBkDx
WZKI0dLGg+9kTduM7yqjF7WH4S7AYEhucXb5rPE9pfSfjK/ZEn2iFofYs/SMaRYv1njRE6Hewvz3
MWC0OUte5wS4t5zlSMVU/pKG7Sf4VvayizMHTU3cwYkvRwO5g4JVMrie0NNxxNOLxFxnDXgDO0Oy
ooPgb1vbijLA5x6XS1LuEboaCCXTSVg9XoSUhBE7b+zjNl9krz35kJyURcmf8m6ctcRSGxi+UZ4R
vOVQjBxzPk9Qq0ojq9e+jNEkOZqiOPuA2XCPkWLOBHrkknAHWfFfViK3JWpDBZkENnKAmFzxNvlW
c+iZreAJbhbOq5oOLHv37PzHaPsOinbV3MFoBVfhnVPAkuv17vRaLn4gQegqig5PxQ9rz9XmaRTD
UZv3nnZcf/FRAzeUDpqGI/oOJieysPLnXq+0kOYDBfCAHgLnys8QII557H7EuJeKobZh6Duonk1c
C6oCUsrr9ZS1Pj5zWfwg/+CTXC239+tIqPkGjLd1H9059qu5z2EHc+7e1NOFyXBYvp+8g2vD9VMi
s5YA+hKghR1olCTgdvv0xUOZSdQu6zyNeUzSW9TjwHNdT7JjMrJf0dl++CW6mzTa/2/6WCqTRvri
4KM8R0FdqgE0b1rhfAZ7kVDPXyL9IHjmgIUgWh03oQthVThW9lDdaQxFZhoj6OfsKWSwUBG/jZEe
q+vIZODqE3j0ZAwgf5abiP6W6Pb19WgLhl8181DuAGoJWo1nR/AKH1FspOOqbgVwcD2mbypBcOOe
yDfL3Go66oFRY7+84qQtZzx/PWLAuciqqBHO1EJcx/oYmW89XnT1wzdxDJAWN3bp1cJnJmgNLduC
VFCpuT8CpRZWSHX++09wr8VNDSa82c+g9QVw2r7LTG37VeKRrouUupTn9HAqXixtFRH4ELUHjXSA
0ssfMjyHUIw3vNmKkj5G2CPehbNPo5JfYDH0l+m7eHFBjKZVH0d/fJtuPQUKD++iF7A7E/l0QYNr
0K3E7VwPbMfOIAqoLPptz8OV/OlnZa5nvfHtxIh4VULV0j0Qu/qvLUSMo5qnjITWQ7+33n3IXqkV
MrhLoGcLijw9auLQcH5gTYhgzAT/eCBCxED31fQpQgcEr36C+B8Q/8A3U5eGWiIyWDf9cR+m4kC2
zj4MrkftO46a72O0zVYgi4Y6S635PwRar14kEeOer6GMa26XnupnnEu/fUcFlA3Esi2K/F7ebWBx
OkmjGhAoMZlybAEiiVKvFyaX2q0KL95QvYmnaOu4Wr9AbDQMZilNGLleFW7dJ/GGRk0ASlAoNWDu
9KMunkJXQP9YahuHAiqEhSGG+3uIoeFvQVGHL6P9N1xAiFPfJsN1qZ+h/HhPTkZDUj2IjSSShcvi
Ozkdx3y+29NB5+tA3OGFz0qmC5q2bmAZYa5K9sl05sEqk6svv3XtMLuhfbDvxST0Gdwq+L/+vqiw
6YZHXGzM/a+Vo/fd4rXQaU+jGKsrs7DiMGPOghQAdk/79kgA8YY/e08LpXRof77siH5QsXmiiZ7Y
z+wEuDSNAeCkUpbGNDufwCIdQAzapSgvQNw9OiohijBgpfPKaWyl35uw48Xo331Gsqq3Ald5KAkv
yRUhZUKq+o/ktUByvWel7Xo/JksfZQlD1QxpT5frv53SgibUUZJN51Pca6zclVre+FC8e0hejCHm
2PH7K72Vlj1QFK99Uiawb9bW9tqRTZ3O0dViT/NnusNuReDOa9pp0d7DF4nZz31EbbYnZwEqVzFF
hZIMXOFD1jE7G8NwOYrM6MQSYH7y9G8zXPWbICmhlMIrKxkBWdCYrKfX8fncm2NR2bC7U4sLQ3WN
Z59tsj6x05FCAkcFGDi6ZJ+/vZT/IjzVQTXYuqI4LpjlPtp0p25FCW7NedvK4yzonzpbdwGhPJx1
lLj+g1YeBE272fqITjs0G8SBRK6uvvYp6MgBc9FMe/yihNLoR3T76r5+KIbPeYRX2zOMNNjE34en
TgkWdxAnlM5gvXkedZ0ZiNYMh1EgQB5qpqT/ZTvL3XpihqeZnNpb4/U+rV1akDHeiFbxlSkG2+sC
MdYnqlgdeXjlaWtRmj5MgIe+mTy/+2HyZwOvA+cFXT4RF/rij56BMD+ZaLbYDBFEijGy+jD/oLjd
5sH5XEn8P3qCEiDE2Kj90Wzs0+JgPgX+ZHuiSCDpzB1fQNlBRgpdLHorVbDBZrPklHx6ob27fLJm
EsWfxHsKEG64gMqAU2sTApHOxAhT/ItbbgD3y2zAg1L7fSPKDJLhj8vY1fs4CiDLJgrqPPk75t1r
0fpU1nUXqmQFd8nRmydMrQPfw4B4e7ja71qqo1pdEN4DHXclOxE8gNdQYI3DxzdpT5G5HpCQ4XEN
OJ5rD86bVqhmt+HducMQt0mvXr0oJczEpBWgdAu1YNAuBo78SAqyh9542Nyo57QpVia6p8qX17w+
KhWedbnFP/f4eouSixDwjavU4y4IRlBUzoMWW4/bT/7cPPy6oEBC1WVYZpU3+TOacefv5GA9ZXoq
kfysRULwAvUfeocWng8DiiFgNuz6XGyVGfzmYsTJ07gT6hbvtxVCI2fqHahNVW1x3VGHdZKNOzZ3
kd2K0dZ1YsBqwfS1AfkGSsE2hzLvVuxPZhuqCj+XeXfHIsNE5WMVPvfxvfkjvcg+hjnyqBOgEs+4
VztAhQOE37LDcrz00CZtpjdCXzbvEHj7bAJHQi3DVKsFaSxgIZfyZOZjKi6RF/0JoI3+cNOiA53j
SMC/I2hp9DHi9z4m/PbxdNcQsEa6e183J/T335GvpC9FlfJ4jNBtBzN6h12uvwV5hLv+6WVdxdoK
Ma34ti7j2UIzHK8qfXBegREfse+LgrE4kv/E80EvMnrjkcZwsc7ZOLAZky6tWJXaUs2zbIF8vRoa
b1iCu0UiqBFGOfdEDbkqg81bbNsP3wj5V+u5YoYd0/s50LrIjqH1mrlBVh9k3dL/oWavVPamFUe1
Ky/AtP54i85Vk7+15zFcJahomSlgdgF4gv+MvtfAASXGhlrKhrkc9aZ1MjEpbnps/DS0W7kmABy1
sofL9nqZ5C+tcz43m9ZGVPLzN2pJnT/740x6+RXqlm8Pq0Ye8kjl8AKwCIW5Z24qZUQ3Cl//Ssy1
svLezSLC6a1sVijnsq0eQ4fO3gM4atkE3bOUiFqFWLWTOvT+FwEp4dmNDwUvyhzDzZv6BfxMJt29
+XqPx2/hwlJg4PxrHFcXolh0Cemjd+xiEt4C5nxq+ZzceHHn1Iqmsd8zCFeldktIH5fjVpDSmZQG
WgDgmaK7L+U8N+fa2H85ACunEn/awf1TMb4jAgRtyr82dn1lIjlMP64G9cXktpCqpF1k/2f/dAoQ
cK2dyNT87cyyApufF01kTUqeMTYJw27zr/eRhj55oU78TiH3OeThIjl2hE4smf1z/4pMSmAyNwnA
Zk3+TfkjHLKk5kG/oLqs8PLxDFLDrPijlCF25gW9PC8tx8lIZZZyuS+YClI/X3GOzJHxTEZpAVUM
+A85++SW3VTdYyR/dpuVXDuN3/ka1q+F+Qh894d7so6WlKoiSsN7Nxb4OroGxpnFyb0qNV3gnm+t
3o5VxpCdQrhET4V4vPFAt1S4mwyWPaxw6rE7sZEIYF7lPnRlcV023Xlicp+1+W0Dm7ZIVVWC7+Iu
9UKQocDVWaTdOVbCALqOdDdA3vgbg5brXhT0jnUnqCF/htF1UhPdz02Wp2n+yaoBSX9NpzRczr/s
u0FIHkdZfMm6T4cRAxZX+RHwJmKJOD/CLT2ax/ru/1JMJhrh+HW4uBR6uhYAJlDJBaIEaO/5yiOO
09Fx/8szK69tpjFtOF/28MEN13WrgWS3b8N5mbbJvyhgln9P5UQQjcfkXDOTiHX7+ydAc24QOgjb
kTiMp/nFE86UmTMx82i+pI4cgBEokHypJAcJnUgZjh/JrRrOKOodTEBzp3ZnMMf9bVTbHXWw8dol
f1V9Ck0UJlqoZn/eKJuIdkgSIy1p0uImYHuO3ffv8z+yb62/sBhd8nEm8N95Q3vO+xzxRX5sIAWd
KK3hTTi5Jyng/WNLODD2lIX7nd48gBMVLxpWbrF2OEYalGFCUnm0qTyiz67zsg4BFfhk9ylhe+Le
8PdCU6pZuNiFV9HCBGjG643oCFroMVto9/ETJg2ZMrs93CcVcVcDuMqnLl/pzkwoWiegYxVjRpc4
ppxS/DCsUkcAAVDi/nk9HrUWdVbZZD5DeTD8BVWaOnmki1w0cse04w5fG16FvjDJo0xG3zc2DgqC
z3CQa8Wkvn4VBk7x4kbi4tChu+qMVuxRqxzMnUpeGcvWg8w7yvLAbpIS52veM4rNcjz9IngED+ve
66Di4ZKs6rLNio2VIpHMYsJp6E9qvkkGOUBwd9UZdOr509/hl58cEzdrn6J3o+Qbe9ZQoJFKYOq3
XVCuNCMLqLP1ZQote30washmmIPiXrs9l51V4l6ak4uicuCmQ/+olvcPe7yFc2tjv1cV8j6zFFzR
yHPgYiNsHhV5bPT8TCw8+hUJSke3l1eq4A7AZJWG6e3g3pHEl9QH6Xs/JykdOOKmKlNq6ThLhaOH
sXnp8Omh/FyzlFZBVBISMpX8P1Nk2rBUcatWH9XQSv9l0zO9QuV7zvF+QYxtg8TXbt6ZQ3/wRdCu
qaEzz51c2YFKx3IF4rl9nKiaBFIbWo33RVdTV4/ihjE/VPbjVJE4Skm72KUmot4up1Qgj24Ol/JC
SoGlwzInbxwB0GTG7Ft2CFP8MFecL/LqrB90uAusOkzgn3WqzKc5cjHuSEXrAan5HBF6Lw2Vd+32
xyPipnJq4fc2+6DkLeKxTBPtjoQO1JEBS4EWe4iVrWzLGlmEyWMw/N8+73sED+QSFyEfxRdfzxbT
Tjds/yYqYCeBzfY2hmuaZ1MlUizAU+nkQP/miZPUXAXfB+vclEEzdAR24k29lgpKmBeZGwsRLa6t
hZzFO7ULgr9tAUuryQ0zTx9HI8dvfLPtmFtsvt7FfMT6zrzCuzG9liSRHzdUF2DhbN+bi+qsLA9S
DO+SyxmLydAq4Ec6B1Wjx1mQQZczXmf4cuYwIFLT29B+i5tfzn5PwD/SImBgnrGF5RFCscBDv8jI
NQs+Wq2rEGBPtC7jK6M0g+96kdYBXB+xZYNNJlox1CsCKqEVa+njG609AdmRvwFWan4rqeV49vCv
Q5IUH4X29R/xsu15H6azuEBehwQgR0oUQxFkWIXdSt51qtbwvMbRgMhxYhkhb1WuG2H8FlI8a8r2
8LQvfEYMTfcY+Typ3uhp99xXiwsgvmIxVYL+fc9p+dhpM1MK6rRuKKdzweUHJAc8Aq8IHtlkZGh3
74EHxpuRwluj6KlThVQYZGL14xI8koWmLKLDfQyL26FupetpllfAvXruYvHQZ7yv/RmxwjzXdBX3
ejtMW/94O+l1EsG3u8BLJMwEVt8IvYk0cNmFRF6kOS0WwwAVKjsl4HT6oioWUL+5qdd+WZENDgST
2AkObEZ+aUE/FwKOiEtzadObhXVZaqFgrk4uyaArtgzeKFu6sciTHqDoeGwpb0SCbJh4OaDdfmw+
E5yeekHTge1t62z/+PXEQ/ciXcvl2VNfDLKGVOWQZ8jtKe0FOKqnN4lJ3FQs0HEBDyDpipxl1XlC
IT+L0DK4Gkirc1HO08BRyWqxB6UJhwXL9DjSYS3Y+LYz4uWfrPNdGv2s2ZbKEILav5+J7sFUMuwQ
E9+XC1VTP5EXv5oEAV1MG7G+1U+pzNwRYXxlXHGgAsGdoVhq4BUo1yrVYshJ6YVytTso9cqcNZ9W
l61B5ACaAJ3uooC7a1OA3XfisQW9oOGXdkQZ8P8s6DemBnDXF0EECv1KeNPn4RegUyKwAdFMKhvA
HIV1XxKai0WbHXEWl+lBI0bGcaP59dO+CeB1UfZUTG+k+UiCUyZAmCvDyFncwQRu5RJ9jilxEafZ
NaWz6qMl03R4bsjGO2vDgGsA13VKTd8SQ03a2fPU2R/01rjkWbMNN4CH5l2XYCXbc5SLfy/ipZff
4zVPKmy6EGPFA1FN112Q3SU1PGWIdPRcMXFqznokRjdaozZ9C+MCXWnUiqNKD96IKRK0zt+3cKVS
RsFm0phglbeeuArCuUV8QhmvqaLAz8OqJ9iYOVeUuNi2ftby2JzhefWQGT+o0rHtomWejpD3ISHD
UBMm8uDibnPpm3Dr33wF5EQvFsHTbRszXY6eUWmf0+vjLSy61uNnh0f6kjBtIdErCmjdYKKeceRb
NU3E3kkvHpq5NgVe1aapvlR9wxaZx0++nfC9v2m4vh1QOU8S/KiwN9ug/sOaYocmWJU/H/ZMdCB4
mfzCie47LtvVBeWJVZdbtY04B5X/AII/9TVzuFrVwe/icpxePok4X6X6um29f9OOCeVZzApJt2/F
n8QomAeUGQcV3lXtx5Eb5GcRDwCBvL4YcPM3XvehHP1MNFvAcysVH/mSvMRVN6P0mQULWqLzeGYg
ixgJHUjaLQ7QZv4hSwTw1iXunxlKJ2sgf9sFV0MHmQf1zFQUt8GIfmmU5UGgYC7sInYVJdbxpPCA
Cc/F/7F0jMa+snDC9X7U+hdDp6wGCeiqn3kOCEliGjHQZkpvudNsY1EWtcLEFR23nDNtmvC/3fjd
eC1FnZdEMCHtazvOwC2/iM6mZdgu+KtQRVdeG1s2egaDNWyuIvsWfw4An8I2vM6JE1ZK4TGRNe3u
FbUezC6rK5cliRqTsJjjD3LwVvEWs0fzui8axjzcSiOrMQ6GnydFyC0cKCOCLWwlpQc5mSAfEOGg
r83SSs7qWYT1epAnSQOhoUkIVIcc33SF+XJCWyPE8uGkIxwKTZgCzMHpAoclYTktNJO56ezLBauA
/fBFSPYmrcaTfJ788q5bLpGoBVcV8i19I8DwNt8xtWT1BfnLm3s2yMxK8RSMmzXR2xE7ZBzuFyTd
yW9XKOsStG5GU3w3rGaroSX8M7M5yQ77AoqDFJgZ481cj1Gn5HYF3oJtajUnotuokZo8pl5VWYUf
BBy5l+vmfimq9O+KN4yajse6Wc/olV2aH5Nvp1G4/8c5lbNpkkPM4m7fm2YoSsDY9+EeHiORSrWj
Cdj9cXEHnSEXUK1vHyocr3QU8aVLoarMfp+Ho65Gi68tBZ+w3OQJUXYIt4KP6xIa0v8YNukO9VVz
t95oWKS6SWim/jP9/EtOmKfV9d+xzOk52bG3pOsWLcYfcFX8MWJjByye+syaR8A3hrrXHGNMEJ45
tMA3blXywaEZGE8zSTMeNhoV3yUKhgmFrb31KC+csF3JAlraVU5aQFRv6N828gp70Q5xIlUm4bVW
r1k9Dgmd1kn0GPbIx6aF1bb2M0wkDWOmTjv8i9b8qB1QwqzOvLudy9/KW8cyUUiHNmZ8CLpJhMew
pi1Iexycusv/5w/IzgiroUQNOUqpBH06CHgBEnjpcv+lLuu1SGeTVoBGb3GwXnbM8hpowdORMe6J
0QzPTs+q9CebJHTZAmekCF0ysL5z0BBPi3FDU1d8T+0qIgYxL5neAeqMmJHLhLhV2SuKEBmwfkX4
bGC0rNnfxwAlP5wedWcPazzbaX9CZT6XhjsDHPXJrCAYEJCxsxaXVT8fk3ZUBrxJlR6Sgj6KrKMi
9OZ1wKnHLDiIFmjpWrQlVADFb/HzuBS1rnUZEhsC/lqHxqHHxRhaA6US4Ddg9Sp8NmaBgRH2UmOU
VtpbH3aV3nqxu1xaVD2tW5KCMA3YKzN3JHyeC3vDDx8IRrak9DAquVliDNvKHzP7ren68cCiXep3
znODk6aPS06Veqx2b8wVJf949SYB9dtYNvCWzqdWBFk16zrrR8tqVy/Dj4tHpkZbaIPkr/zUqQPn
EJeG4F6xitmmgk4uLLQLZjsEo0Yy2RUuWs23ZVbfknj1wm0wv+4kfGtUtEMGisK5DTiKY+bIuO1r
lIeOlG947eqM5tmFvdnR7UrXITTpIxETWR/cADfltUh1xa/Q9WrdbMCLGKixeBK3tXM31jbR9Svp
B4w4zrTj9xiXrg2UM6L016JfOqcpxokOIfllDCNyupG0kptKU7TZzzjOPUspPjiRo4K7Ca6rPixn
j2Lfi4VSAff35w+0MwrTbuCJt4+OUAn79xWyOSZRPlFuzQp6NeEOi7pvMjWQiByvpVudRoS6AbGI
De2Cks8KC8ipyB0MHluJjmz8Q+A8+UWrwKnhWORXCV02NFNZEbgSmG3MAr19s6JsO3efbX0GGuFC
x6uQLjDBZAL4qS32Ay+fyZNm5J9TqWQBIJV28G8RrnOTmQiOhG8F1qLJtFTsza2bVvns6TirWLlG
rPLd08z0eixacs7jJDCS8YfJVT6I/pjEUrVSILmcpBaMIbquD4YAoXU6KUP1+iHYbvpedG6z6qKu
QCv/2MEoatkwOQggrdMKzoJ1ktyTWX1+QUDBlo+CKkvI3bMYBjp7N3yh3EiUhmswVoxcytiwkcef
8RosXBcElE/3cAStb5N/GVyHb9kKUT+yRgR+1zh1X78lxkyjVSZAXPbXqTj3Ia0GFXY1s4IkCYOF
y44cxsQHkdcg6HlV1RvyOzwZOQJjvnRX3SeY1Ov1UNNH62cXV2za+TGhx0WhrPhiUBqO2WTwPfen
xewMBFsW3MhT1IQ9nlBChPhkOCMEB4TK9C8SvmFf74AWtt9FCah/JF9UR+1hwNofkG4x1tIeYkNj
KtceUXU2e4Zatcms5YyJf3M/9I9xcS6SOeb/8buIO+U3p1mDkTaRZq+F5sR1RyVVAnLC0yR1+5UO
RLL+zEqlqrPzJLeiOqRWCXld3y6Be3cQtDGT1wk03LfoJ8ZzncpcT61Aj5dbP31X0nD/adBV5uXf
NRU7CXe2irCC3QJX2koh9W64zZyito+2w2U9HB0HMIy1/iHcFEijYhFUQE0V8NzUhfA5DtmposEc
5LxBFg56dV4cCuavg7vJH1kIpeLJn7VneF+kh5p/kHKResPT2EBgg+cPt04fbw1kUEK/Hla2lF+5
dmZ/c//Kvo5jiHvDgxz4ROxFfBYuFqnV6Fnuh7ttfcWCA6mfSWdoqi+oHlrVzYrCiYlNVynw0ndQ
Kfo4JPiLmvHgYiKEKVyuaSEvXtG4EZK8J5jt3d3f6FfV/upV8aa/M3HNmCQiwgJWA/XDJqhzxP6u
+IFadQMQkXKYJYUs4A3GHdnnYXh2t6sHXRT+N6OBU1t28J83JKxr8LQHl0cVsEXGjNZcb/zTwdVq
63O/z6nXtgb2STmLGfO+T1yUXsI48ZC/rIsVGX10p0we/jii25PknR4731ekyNwTvtbkbyN0s3v7
ChErPXUzqKf+qNq++HByKYmvHyF6SEpvYNBc2eKnSgmsY2MAAFocg6i/YpAF/lLu2xh3HI9SZAyN
fyuxxbUfnMnmmDDxzam2U2ZzGuuccZrAmC/w92jpabXiHjA5myINmply6osOsFc+xgpMAIylifIM
Wt2IdJdqdomgWThj3vGOwDutLkVuEBn1usF2YTGo7aELcJPWKc391KpO3BFWDKmOuRWWGsYsPE1/
Na6MWLBd/pcMfMfSsjSTCwRwFZv8y6QK+YYFymV+t3SwD4IaMdBK07G7NlHhNcD7hxles0qbB41H
u2MhPNz0B3HnSVYadQMfdkq6EUP8PwXuQYv1/YW3dP20KmiR6CG6Cx6V/x4+9P/U2i5HqW9pkdNs
Ukctj1NZk4GSrwbGZDxAhf/tf9z3UGrygKTLe9cNScn8rk3bt2tdJq9iawzavTtSqbrApmReIkJR
jtcKPLbaREpQWWU4vq8E+rbHm3LPkg3ac81qfYHvU77V7yNWUiYytWrRZlr1qbUUejC1sEdYSCHQ
ifYkFCHX6riJU1Boxdn2LEw+cOMiE86zoKE0EjyJUoAoyvf/JCcu3r3kb9WmirWw7ONjKS3C5nFT
Zb9fnF5w+eBplOeGLEaLITg/T1GFWU+UnlB9kWJoBx1ZpzWLvscIu8xdM9lyhsqAJb+y/QXIw1hZ
+jYiEbSPgxMlJ0mDE8KdYMn2Ao3NmvrOpRgWXsoCdtRPLMg+rzEaXEDY1+VriXt2dGbwCcEkAtYX
kxoRxwNqWAncwVD/lJirXw5PuWTahCOYtCH0kClwKUrl051oHgLn7KN20zfDUdyzTkbmyD+SMFfL
zgXmQUq9t2PLrzShlwKMdPmQUmOKF0KMJTJaBUncBTG1zLLa9cJrtmI168Nak/yeLQwfqEYm/u+0
qbG1jo1hXSyk/ZIV4+s6As8yjr7VZwrwi0HQRw11WBYLVRY11SvnhJy2wDaH1Xq+eESVyE+z/LLE
dyfy1SWG9ka0TLZqKLhT3TPq0haaG+I44GOMk/HFzNRhytpBAdCo59mSBSwZVm94rZsTqk+ZAN7c
Vl4bt88KsoDNYuN8piDCUmhfCJrCweB7DXZgWEqbJDfmMVZmoTLBGbG/T4K/uAL8PZPWpy0jeoEw
8LZn5e3FSH+AFTmXCb0tLmIxaRJguo8HO9syZcMg9nxC8UjKfX+atp8bLhdf4/PH8w1vVVcO/kFI
Y0bLNmzGY63n1btJpueaq8shtykFeqZt3abL2UTNlTndp82tZKpxtuzQoEdc9v0uoFwUwXRfLTEc
E9GQRLDsL4Y4wq20SeUS57FEteCdHJI3oFSNSNAbj/uWtbGB9nq/cJds9A8b2rYtzMUF6SovMQue
ItlUouWp2XutlIOF6xDRdYWqUuoSZbs/MznoRRdmN7+JmqiS25pseHz4Qhp3cO52Z3cWrH3qMLqG
5PuQPpHEn9dcxtepi7Az1ZiCf7dgJ8u1TJT61ZcFd+vgqw3z5phhsNXpX4MmPuNcFdSbX6DdxLTw
Fiixr/eGyyazycVjQaTHzvuJ9O51bzUWLeUmTEBWHSm3Qx9efzqMWeU8K2/BAgqh6IbKazhrCypX
dKQDcD0pM0gICnmccvWPxFv982a2ZbIsSvYaMurSOdVO/jDbg6oE1t2tqWwkLu2OH1qjHdW2CAxr
HyOwrOBI03KY6x4pipbCtKAi99MT9fiLPm2ReKMW6l97Ze469sGCXin3sAPC1yRCnu3felmTBFPV
phUnVKhpu4zl73PiKP8zTLAa4UXkULQgL9JTcmkIaY1F34gteZWRP1IQvVO3aP+WCsCvom9HBMIx
YIo0BFnJHp8qKoTfsZTpGWFqgH6Q9+eX13g7sXIegaUf75l5CLG7uyBvc5x3ZlQ0Sbw6DJCsZDtw
s3NC3F22T9tKxHnhDOQHLPXh7Kdex++CGdtvxk068KN8jnwS1VxK/fUH5d0yIClQWguZaJZS41rs
mTVQMrumnUObFQkhHoB/JUmEXXUJoV1QTm+EY19ut1UVWVOwAEwCZ1kVddZ9ceklorpc8TKp6qgE
i2Y1iE4tPzeWYLxRXob88hOexdVpB4J/48Oq8xavVtrZ7StdExGSYTC6u8VkZY14sGnO2Xac/tQV
uWQFEJH1QBaf54eNUwyc3MlePh1xwRSwY5jzixWIu2zcUgBldO8GdObEhOUTbUiv5kuwwvODUiPz
4XPHeM/1MgIVswYR8f8rS0QIo14Hahvuw6cT02BGHZ16ouzt33WI5mvP1lxr+3aDkWdYrW+6aKVT
gtHr64NTI6eFONiZBLVIKmF+Xt0NsSW0z+XfLMznvlY6oA4Ic22b0gV9YlOAWcRUYK3I1uwYY2QP
rpW/0tE5zv4E8gc5rnnNRlIz2YGiC3GBByujAKeYYLq/bbd5scnd75m56t4InVjuxVGf32GrHfjM
RPPwFcxpgYpOdyS2nSkF0PG91x65si5RxLbpQG/w6CIA9SxTipJHvHlTrBRdEuTnzb7GroFKkYHG
PQ7a0UYOxhbabgGG6Sqk/zvV6c90Y6mXh86dCh1dJQY5CINAyxk9B3z9JyBcYAQljEPkB4Dabzkk
6v9NmOe1qwt9dglk5dDmqbrLu+x5K3LxzghD86zYzACwYPzAbHFJguoKTRVh6x9bnZItUiaKQ6jV
G3sASLrFdQs8QG5/i69HGZM1ZXyt4yJXpSO9xF/+jWWAAjpKKR+uKhV1FPbNN7A3ZuHFBlP3s7uY
B1l3hw8oAo12vJaCR6Tj+8XNTSihWvtJX2aNtxnaVnd2aSBURZn/k9yF+76sPErdqbWms2uwOJbl
OL2/670Y6pXeFhUVyLPfqJp6Wocjguzd9OA4jTGs2vu8vuabkG/Kq0DGj3Aw9h6vLaioWgXxzJYk
qB56mieOYQMeoRDyR3/jRYyz7l/jLwuoHkoz/YkGpMyILP9t+YGtpOHh0ahPSIOWRs4Pe0YtH107
Nune2aBwUJdv+yjPm/z+j2l+1NceK9q4veYiTkqP7MgJZqSrPsVdWsyCK2AQEVv8j+Z3Di6OMbTS
Fq+zHi2qeH+vEO42Fdq0SWH3P4Yfp4yLJIUKVKX1c1//hvPZaMWPJn6hAZijbJTlZuURUYlhUMZi
g09bwp0S15Rp/Zee+/aVUh1xjK/GbjyHhqquD+xWWxkdDuX/OtJjSYWitiiDkcuiyme+Ql16d2Kz
Jq4atvKLNh5ZcjCo/cX8ejte0KrTCgB7aEI+uSErbpxys9JMO+bdCOhts3ZEgtTnjPghGbCijSKA
49zmgNHK4gWMzJBgYdghsb/UxIAMxfV0jkRDJlxGdXX4eNsn2I3z2YxktURq4lr0QKsfekgQye3s
FrQSon1jYICHXUgXOvHp7Uky6UMqXx2yGLP3w/oCKFdPLz1j2s8+zpRvsuEZ1/B31m5b+0I3MJEY
q/YoSJC0T5Imay3GBU+OgnHiCTHmkoKedO2kRSHtMCvplBdIkdxhJh72SdSpgDUgYFvPiEPf9GER
gyXEF2J67gh9eIDuLmt86R8HFe3C53MNOVX82nawvqpEZThgXbWmC8rGLugQPb0AVh1P5bgTGXR2
hzY1ldYSmJ22bGz9/Skt2iWvIO3jNJIz3QurshuXd0kTYX/Zge3e7wuI+Dxvkynlr07cV583Lxbl
+grX2Fc84eE5Qw04ERUHAzm85m7ygIeOhSUFbLwTETAT+Pn/BKFEVrWXnYGOwFWDP9EUmUDSHqzA
I4xOe7XEnDOvB6afrXTkGIqyGUccHVledsEkeNd8pJAfNzOExvwcK42Rwq7m0ObueTKYElkavw9F
lTGpY+tOU6fYex56i6QXdMaKmV+s3nZyHSAzPlNkYAAX2+lLE70453pZLF7RKyuIY6RsQGCHtXhY
kkq7Mi5Lbm1PKJOF8nSF2yACN7DuQOvCvM267vuDCf2oSwubJJgw7rpqf8hE23YzpVDyrXDYU6Eo
xHf2QdPoRn87CTEe2rMLr0uqkSnUec4QvOetvMjcLVKWKw7AA2s+bthGwWIUS5VqL3p1G6eG/+Jl
kAkdSb2twu+eK6S6YrYW2NWjvmsjivvmvIUJFLDtsfarK1Amp5TFzrDj9Q+ku9pspY/ekyuRub0j
eK3j3+AKz48k1ENgoYZ+H+60pR62Oqsev/sV/8hEy0+BCDVZmWZgrQQh7jzECQc5GhMScp+Jdatz
LUSPFySZG8FWuj1JhlntHN84r8owmhOUZVbEuZaCbYKEcnojXW9qt3na4iO7WYtM/gt/j/nQWWFO
GY/DgJc2bjcZ3aqqgU2sVwDOmdY2V6P0BIcopBtdPSc40Q30O6zwKWibgGoLsPDmhPfZjyo2Eee2
iZeAcDYAAb7ckwJN9x9+1ev+y/Tj/BE5FU8IQBM+0YGu7kfGNnJ63F3zzgUKvCrRm7uWe2ljkvcE
IEmVHoO3nCvE76KmkCPJQS7itUQ7y5LTuAVN4LTk/EidGDrU1Y884LMb36FvH09EnEAY/TkS+uoR
yuH4mCZuAQejGf/Lrijh6wRdABbPyNqSymfBx1MhKbVypV5AXfY/hWRYHWJlwKLL/whtmKAAKD71
tuYRplO27mhLTK65nqBr8KTrjIOwH+6Ei8QkFsSBXgRQ1vjJZPvJmT/R/MDErNGhbaZXANhNQQBK
IYbxUZJ5oV/5sTBMIwBeTZLD1d8HSnLyUgcy9ly3RNtbB3HLgQ57vi80k5/359yeRphKqQ+Is6OL
ix5+99UhcrNJzH1zudy0wHYovPk7i2/qq7QqY4/k0ZubMqSqkxUpxU0esv68M9kfvfiiVtsz7OL+
eFDy5aSicd+cL3hYUgFtAPYBdgFs8xXLoF8UKITNJCFlnyjXOAyRXBMV5wWLz3/giPqdsKGFX5z7
X0ULJBeI4LLNHZWr4HYqw+IgbKwzGU6Nce/KMAfVmuuo6NS0DOx98WatH2t8p/m18KBU2FGC86oj
TNfPBnAjzszENRnD/TNhryvPkENg0/HaBiaZFSLMMluz0jVUJsfr8cLr18EnWYoD1/iNuAMZZS40
kRtLhcgVb1bq7cFhruacs9Jz2ygmkZ8glMA4AzBIgED6/yQ1KgqeIMXnnnQW6p017xLbbKN+zjwi
jcqTtAEjLWIrf2AwHnLKp8payoZBZpGJCdw1G3Nfw86Dmb0NeeLA5brXBIqyOM0ewyWGDU/u8nGb
2hOrOoNVQzWT67qndZhPa6xOYAm+WSAXsCSVBZdFDsJhU2jz649xnwp10m412QJmOVU9LQjThSuJ
U4k1GtjxvnsCeUUHN3FuKmS1hAAXzBes0k3pcaRJXMxVCP2z4SRCsvn0OzlJi1fy0rF1N61aB/Xf
pp4IIFaGnctW3VXUdAIvThcIgkNQjWM2l/Gyeu2N2zeiVvpJTFGH639mCnTCEjOtO3+DMRw/ADmj
4jHSFboQAg2T/p/B9veidXcpM8YRF/GDYI2Eyao6EluB3lgX4Wqk2j6Ho9cBIn4ZSfm4swiLpGgf
dkj5Bb1hZd4pIOU2Y9euEVrO40Rh0TlxzjkcRQGaCPr6dYQb5e3dvf3qUMJbxN2GYNZ6pPm+ikOG
ZaPG47+vk4VMAM38lb/Eh7Onbe5ZWwD3HWmKWvd0a6sf+BKGMfRW50+i8Txsefrbm7yd0PBU+o3s
UEjzJVvYiTJEIU5YB/6h3MIiaYTLKUMAEifYQ4BzYZNnt1xYMtn+Hzls4sN/YJcS+4neo0AjO5rT
y0wMszn9/9DzhwHHzAO1wRj0IFcksfH1nEsi8zy8mNMxw5X3NuByKS4ne5XALE9wke5kDCTvwUp4
QaWm6Hnt8GTkmuoRgWZ8aXjr2vSDcDhAywpQs01VAwf7N7OVM82un09lwSXd7R3tYwD3RI9wrtNR
D3m9U6i9BiRg6TooNc5qy53p/CeHYpnl4vUlG544f519RQt+dP5va7UwJYo2niAqlEG17EjhB1hp
hWN4CiEQGLHxBsCIdaZBsML+xOHD+iffUZEZhZHWX62DbyRROtvzQ/Z8sdSJSoxgUk1TRPc7I3rz
4Wo6CyOXWEfOFLiMM5ugY8ldPZBm7ndXXxIoAGoiWA/80fIY0rP8IsZrmQuQD04b6dKT2CDPSHnm
A4eQJbuc5qsFQT0Tcd6M7A6uEm25kmhJepkJinlNT9rJy/nA19xmbHNQWrcwM/l7lS3E2R1IY/Te
PW3bM523JLx+N+g+OjtPOjt2jrIPXE9KIJ2xg/pH1Fzmd531A/OCjlYCqE6E2IoB4JI2Pamy/Y4u
5UmOIe+iD3PWu+oTcpN/8AjQieTl06i5U97lwUxJuRgHn9FXXucu/waqg6IcjazzSYtc71BlsigD
VytYiPY0UarKkhwtkywDCJB2HIfo6Nvwd6vZW76mmv+WUFCp1QqGCvRLfEhStUVU3Wgj6gvZ/COa
v1ImvPB/PKsQ8Tis9C0SFlFX3GAKWtAXdNfiJoQvdf24eKXyD4FcVo+5RXZHZecInGyxpb+4RHpN
SIFW+umN+/UuBkW2ZErl4T3zQvurBpy0tiOW+NriAIZWJMnfqCsTszqRB7KXfEpnUwKSWCgGENeh
EsgxCOXm1lL+8higQneDaOp7mmUAElQwpezJ6NUWLBoycNTlZufw6AuVCPX0Vuat3PrO+VklpfMb
dMf2wh/f2h/98o/2vu8PEda7YeSUXtD80HI5M33QxN4axmoqClhb1hEqHy19/goPN1eG8gDF53BS
jAuu1NFfaM86bJHxTl4teA6gAs0LLwjQaZBcn6gmPyZ9KFqpZEwM3FcnSDxCA5tQ8FtAy/+Yubxr
xmGP9N/OV39QIYJu5baMR6FOJ/RDk0oVtiXHpUADsgmUeWt4GkkmiH2qOWnl103+NvDon5+u/OP1
Rd+Lw7fnwB6ZlRYAzToBSFICZafqSLTzjsFd+8hgjUCB+Ytm5JszFYAvyd6WkA6z4XToaD7uFhXC
ZgPtILmBqNRbVPgScou5vtpvV5tOfbJeAdVbZLsnvRNsWKdeVmfauJc6+MYNqP8pLuzjJi8EzU/Q
IYnXLKdw7oZdZPkX6cRmiLjVo1ZGVKgn1oAaLiO8+Dninl40pjDl7iGcOedV60ogVrBL5HTMFTEk
6Ngpx5F3rj3dQ78oShZP6+Ba4hodKRbK1iYdedoM/7xxaOaKywOFCsRIPzP2rOQjWyPshhNoXG5n
ZOCngOhSl7GEmnRpQcNyltA62BCKiwwOAityEL9LqGi3qWDVGHkY07WGyYAXmYOr/ytmYwzNnr6M
3yyMf0N6Vo92ekPAtEwnUDeeYbRnqebX2y2NqtuYHbHoHc9+VgL7tZbBOJf+KFAhGA2ShXJI8w1M
AhXcXBCoXNJo925V7SCebBOkQWKCp8A+VdaLOeVpiQ10E1SJDw8JyspbU90CRimgdGiV+/z44Px1
GshKvPkbbe0mZMORP5yMICo+M3iUfqtwg+DsynTVlcSdtDLG/qxnAFOvVa0mZNeMcW2ERtTzx5l2
SE2dALymNHEdgGWKVKsphcSJcf1YqSw8TfgBsm9Nryqjy1av41/ge2w0TcYF7oJ+PMZlYOZjP5cH
jDgq4EOqs/bSN5LztDPDGqf6p4MzKNbcSUkxMWUlEPev1MfSyPX/4RdU91jq86v7xt/Sm6u/QaUW
kCy6GD7xkthUGfFA66g6rhB3QKYcAZwq+9KunZellSoDDVR/RGynnBk/1HC3Ib58kIS448kLHYsT
0FIk0FUvEpkfaBzdp0tafTBrI9IsSC8fADH86SBhCOofVQKqtCK1tSeUgtZySya2HbqC+hI802sm
YNNu/dMfLf7dcMAnV9FSY0jUwToW8k75Edu59oGDdOIU+NSCJkQDUttcKcecVB1pTPWfJtUn2iBR
Rqn/q6aR8A6DOvZsGEfxdZ1ordhyKcng5Q4zIX6seqDLJxsa7LZLyvbbiUMxZ0a7ncEUfUvMDims
vKtUZgZgjuJF4WewgBjd85uC83uw9q1ZwsgZ1YFS8/kFmhx9OM1D5PduRN+OlcJwTWqZ0FUa6Wa9
HS1I5wuS32PM5mIWS+wUTqGRRLjaWsdgr5IaIpeeWs1gz/OrWLI+fjKVOeT70E+tMcTVPafuUYV+
KJtEK+p2e0hidMSRVKH8Nf27RWt5m5wloMVROKNcikAfdR0TrN1KSgMXGLf/wFBMcLskLiOLUwCx
fvoP2L696AdwL3gg8sXVXsWZZ55ly6hvShxYzmqoQupRatofAlK9Foi6eYxL/lNIjFityGw2O5r5
a+urvbldpbw1ivuV6h0bfRsN+muYg4zVHj83wmoUt/Wg6lAUP1ij6tdD2j0wGJiibNTEB5EIdRQT
n5DRVG5k1RqhHGXGBFuGsrabv5t1Xoh7ddCgQP68iaQxpxPApQzihrM0CzbycC88JqwijNd2BrcD
W+o8J5l362Uf3UR2LrWen2190+7RgB2GGSNRlbiEYGT1LT2YXBPKKwwshpKK72LCVvSY+ZR1HcW0
yRGLP1fJ6xs4lTmQGMLFCZkGEPOs6yXO0Dxb63L2ZpbgaQ9tjSZxtG+rHwyNKKfyMfFANtDAwu5I
Xuna/H62rvFxG02gzLkRN53JIou3Vai/koXEERyVF2N0P3+eTMFFTK5k/YTX0nSGg1KUNK0YvFlL
SkA4ru/kfZa+KJuORrfDVuJyf9rjt+AtES60MtTuJrFgZ+Q80ghDUF32D7e5IZ8Ed7X3XqsHhLHm
4qePiXthx9VvNMUWFYKBerLfrEkihfpzHbOU3yaIKr5eM1BZlaqRy48wz9sUWSEwuxKl6Uk2BSRx
/JLfjtHGBNlQ/PQLPTm7Q0FGspUCkUaGK/2gf6oe0L9U5s4yapM8ByvrZrlBF58khBJbBrYySeIL
Wsvee+pyeBJdHB+p96jDcWyuvDsevl0yQ6fVxDM2fnpVKrM2oYKj1RL9LB0RLn4QxhbyxRZ0yZvy
Yf79XUjD61OBPqy9AqvKtoy6rIHnHHUNh4g1L+kNYX+NMmwT9Bex6qXkb1IrxMX7AX2cVnqAs3jx
FuxPCjtHbBlmLUEnxp6ES46MexxLNm0xVwQTvgFIlxL97hAC6IpBjv9pg0uI4JE8t1HWmHWvKek4
c3665cWYTx4Cfolbf3SSo1WJ6GiqCVoFfcKB90qUKSFhZEXjVbpzddYgvtxuCh7dazQgj0+BDuWS
3NWsrY8le6TYx2/0gYgcz/LiagNzCthReSKwUJSqxxI1mLO1XjJIJ2nhSocDd363tE0W1A0WoI6p
cm2prCUeld1DNGGDwLCJVBIhdkeYAm6SMxA23//8+NrMGwSWPq2yT1v+HUkt7hnl6eTPCl7BSVeT
N0u3l4DPVdDv826/LttGjtgxhQMrzTiCjmuarHVgk8lVHHSakJWdVBQHQ87JQu+iACqGkEEDvM83
U4kuho9y5Kkv6R4pSKWZvjelGDIE6bfHDczuFgQ9UvX3DChUHC7cG9Bgqroq8U2bNCvKC9lwzYcU
Z71CAHqKDIKjxPTyK8HznLTlmJX0oGwUQzxYMfaqgEDypEs8Wgnl6S/V05RVM5BfyFJqYlqaKs7B
+W9mNztYcYcCoviV8eTXoiTljR2QMKT7zz8GT7XFi3606YQWK0eMevO3VHIMG/N3kaeq7Lv7cDJu
c1JXNyJtW1nY5ihqFQiVvgZ5cxsI5v1qWvIXI++mNRmqM33PC5yZF9gZkBIc5AHqm5ss75C+CjOq
TqXS0TXGVSVglnqyW/Lq+iDCwe+n/fNgoUNkAlsVW0Ao9U/yYkf4O1Jmy9oLCz1NsFtchHKBTmY4
3n9ilCP+ADhTqtg3TTEJQJXQRelymEqu+O2ZqSf+cgbo0rcsTKO4sdVDCc82wyC1tkFARDqWqK+k
Hcfm3+AqhRDYeHhJZLDAAq5/anywUMyeqKh1Bly/BwLybxffzI8PdaL7dk9VlBQPS+GSbsn/1R6V
henuIyiDwq0nA2X7+KOsaGDVVuP+3649zNegfsNhp9VhL4QTFPk5KJfYe4BUWpC5JCl5NzHoHgAc
BugpemIdWP5ynC661Z/6xCQa62aGCnB1POGtVx7LrHRzXRGKwdeCM908o5PXcBUlmmrbgwgbREk1
TaIQWUNjhr6D+cW+zUezB4ZEmv6s/05dvbwgRVyZqlg6SJo1NrDcCYJoYkSACL/iGlgaT8ULgegt
yPJTS+gefVlVLY/WxUycmpDeGRke+0oHhAH9SgPVazrNGAt/ggM8ptgnllzCCXyfpGyiv5DFuyKY
7Vq0v7lsKuj4nvGkCxmfy90i3/ZTFWguuT/egI6pJjj8KpTrvphS0UCX6ObswfT3/jtajvMNO0A7
QeeSxt3o/mR97E8d2PFtZm2obpsqqbSwE/VgpUy2cxB9osmurl2pzhWg/cINNCwu1RDDMplqm+2s
7NPtKIxfocrClN0Zx4K0vhwQa7S5+vlNY3YhOJP+oBAxZFsQaes0WrLEK16/x1k/r0KSFAV3PmMn
KmSOxPBvy2127PU8L861C77awMbgaicseoGih7+vd+pndKtxAnc0qpZU4NI3aVWhio9fnMyJU7z7
rRnIJ8QXksx2dMewaW4ElLYQLvNTBZCUTqkWObf3c709tXys/HIep/ghdfhJsuOes21X+U+u5pC2
ob1Kr6bpdpj+z0oqqoBNB5ST3Us6HqsmyTyK4vtahKrW3hcTxgGkP8hO94CInjFhuhOoHeK0WNQf
4jlFL5ae+maJhMu8IIJVfJHkE+7jf3cKeUd2DhQllf4h7RRqEqVwDDMRXxMhBVwxD7RKvG1mZPws
vTyPlUTPqWRGqEYUFwKDP0D5G6qksofTD/7KiEmVdVKdl/kth0/3jSS67wqLrpoOiAo5zpFx9gHx
/5M2YA2bFFqEgHYtrlk89e/Nkxic3C+rLoCSQrNZ9FLWN45n66RDbcvPCKbL1XFpbmD6lxzK9ltm
s6WH+NIwrZaTxvE9zuxMCAE9LAjE1x6IpzFhj4yrbGJdOi+3hJRpAAEVsBAk6vtKm9XgUj2yemJv
bNU1QqmHeypmZPaR++6ZYGQX8N4Qr15TVtYcjtiSbj+bzPyrEm46O05MLFeehyK5Jc8ktSm8r/zk
uVh4L7xgyy6UTIpuqU0uWJ7KErpt05ZyMqhB+lCVmcU3lpqpm1DVhRkfh0coCyRKlbr8gBgGk1mr
7Jaxqj3a5YXl+eJCIdl0N5hUTnqHjXU+xiIH8ik5MUvcRsjUotlSN+oEwJ4+/iW9lcRY7aUJNgRD
6OMO9gkIX2ks5tj8+GZRu6vrLm+XtrmKhIad0nf9o0VocjUvwLTiEMr0aytEDOLqznIAs3A7tpIx
NAWID8JPzKUcfO1PDcfCWBGnjDJXNHQnZ7SfYpUcgzoLOGFYMrTfCpSkVUcEt8oWqAFWqAWdaBI8
YLQjlaujkL1OspY9X36EykHsTxTCkQ5SIzkNbeYFWPNpQkjYiZvcFvxooQ+VsEWR4zbAXyNUwlfH
YuUp7ph0y+w6vo5bYPWfPeV7Xda5LrRp57DOlE8hIeyuL0q4IcP0iRcWnZOirRINpRHLrw1IYJ6A
/s8ORMFY0j4C+dPBbpvuEIRZO7RTN8vwTNxpuOg/QWt/6hyuduxtKKcz9mVdF6GEk45ugA41Is3O
ZCSbenMWKQ1e+XUok++4WzFuPir+pQHiOLnyXPl5mEUUFHq7AF2yFtT68i8vxM1oZbfBE5GTX2t2
AytZYLVAKgWkK6zFh69Q6U9fVF3gFxnuoMrcWBsP3TicU/efqBNokzgIZHI6H1WYDXs3d0IGQXth
naC963tMD8EVOQS8vgG9VLNWkCeaMHkXkuy5u7vQiz0U/nNhxtkmnDDWn24DxhoQc60M5aXVfbeB
yJZ4UDAJScotKJeAVoPYTZcx3wmoBhboMypn9IMANpLXYyXbPExHOsPJv3ThPRhKmkTD+7BdHb8k
A+/na2B3JU3uGn9j97jSPor9jPbb4B8JOgvd2iDfVp4qLGkNcyk2NA3J5VQnUm2M3hNXdzvObWQM
NeTWKyL9rYm3dfR7A20rxMehWKnenQFNmzowmb+OX1Ew+tAkyupIPb1tEyFkPPsdwkibEOPtbHfl
n19hzWz5T7O0TOArnS4WSQeWL0872jzs5yWu3Kkg9B0D2cOIv4E3iBdYBU1mA4J7koYYOwRpC4F2
ao79dH8gdsNv7Hv0nf3bbPnfgCgifkx5um0aaq6/L0qZMajKYZ7l6GwmKaKyvnH2erNLio5lmUjo
AJrXNcB3iUowbQ6PVGLC7wUiUKRoxJvyeYKbaRjvWXRUoASczzlxCpOYF1PO2Dnc/+hCYvjlW94P
7BRIdRdLwpzlOKrhAdYShzXANzaZbOd1Uch54Tex3tnTNu0cPxJBtXSFrUfAMUuZW43m4wAmWpjC
sQPFnPWCmCMd7d3wFP5dMOGkldU05AUO10NyfbTUMeVcaFYgmao6NNFiUGstfOdSDvtVEGmhy13U
5pq4zFFGNwWf392WoNxXjnHsUk2KCILDaElpjSROwRLkbHVIhYgAjX76DShfSVmAGq1yodZx63yq
yn82v/3B+GvIhlsBT10Ka7c/psevi935ZtFb/q71sLdrIoeJGWZJCJr8/weSgE1hssqeBVhhAJ/K
+yPlVv2s2616/XZBptZnaJCCl+ke28GWNjGTeIVPlMvgHpH/WcQcj7TBXeSrWzctRdbXUb4hekDu
Lz8qZLk7H9y+iEANvM+9ys2k7JSZ8H1eR1B3/Xa3SkxDhDSpw5y+ZZ+1FQMkSXxcJgKIdE5dsBiC
xXvYRv6jCvuPseECr4vHrWJAtXpir/pDloDTrc8YfaoeAVTq2aOaIEohFRFxpqKIVYdCgyJGcL0K
lVZ68r+nQsAtqgGOsUE3AhciMQRrDleJvzVw70x2YfydwsWUdaHpKcyZUqXm+HcI3TIlP1G82e2n
DzI5buzrDjIS1tC8a9aBtL4CfsfQ36Nyhq4+HbTyyMr340khvIqg4quwj6FpfPvjJmhw8EJZN2Tn
HDl7d9J4NOlwyughIqP0I0MxQaO3EH7JjfyoUTM/J/4SYQpq1lLZ2Al3/f6tygnQ7cijZPY4EUDJ
azFRkGimoUcMeUqHLugPM5IhUs9PTziOhOeRBpBW3Nch3+7JNdJu7cInPO1m8tb9NBfO/kXN/TgG
uvJvoOpGQBtcGi91bLwuy05NveuxAnZZv6rL5OsO6uIqZZMGjhNFIxtxY3mG2NQwv1eRyh6Xsh9K
1SlKF3CA4rmmmmA+ntK6N9mdAPYNWFvV1vWhSpcCLgtqtkjDJax5FyCCxrehM0ThtC23HchRvBK2
F2TYB1hxVwSdqeV7AsntrYKf7YxGEWRxbQQ0mVFM1t+rK3wNh/nOE6EZCusoOKVE8YTWQsBA3H8t
Z3wtbJIosS6ExDC5B74/P/gt6ttPy0Mx7VX+lMWRW9iEnMUqAwW8a7QTWL4k8NQ7bgS7g53Lp4iq
mj2bVYKzV1xarfnUHpDG6VR2MPDHcz8ZDPcGE+DbgNG0Lt6XP7WziPj+WbLgo9fQuVHWlz8OJ4/A
sYTYK0/LMNnH0d5s9hhWqBA3NBcz1qvj8oJFDr1+vxqmPe2kOmp68alyW78rtoM07YllZGzd0OP1
Jf1aAA4EXDB/xQDyrFGDg9Qw+1BJJBla9pYhJvxrjU45y/5IsXfPPjPoYd18dPkKQ4O5FVl140YG
t+aa3LqtXuuRFbuZyd5wD/WFSAmBi5ofsm4gxHj6cq9zSsjAtFtiJAW3RLyQczPS/gHKVSsbnjCf
e4A7E7rGoqcamp2ANhboLzVcYUmFAadte/ORqXwnvEixkQwkIpaq6QMxU1Bo4MjSIl7VppTkjCCQ
46/GX6a8lGS/82GXn43zVRaKZhNhgSC1QlycEu3D1h1lXSWbWjnjKxiF4fzNkCiGsjHir80YN9wK
9McVT5+yCvwtkG4A3Oy40vre4UGBKLOAGY1Sb7AjAW/tvZB6pqW58oSiRpz2D7BWDnxb9XPB990d
JFucGxuZKAs3T+PpBhGT3g9yMlXXl+d70DvP69i6u96yK6RxUxDd9j3+9Cq0W4npWooohzM8Lsz+
+9jG2HFC3npV06c5hq3fdrmp8igp8a5rP8bcmlJqqMhX5VlpO/3T6jSAaDy1qPMuLRmS85s6VkuQ
2aBwiiwEBR0PEYLIyj3Xh6t/WZE71oxHMEIozyYvX4I2XgS8CtTOKunhfBwIef0ru9bCzi1Gnh1l
LFgFoJ2dXcAGxwDuLRs6kdAlh20e7ip4RlJ/3QxleYAg+SG/DtnFOtLy2xJ4QxWAU2Cj8uk/rfne
1doZ6sCq54NHOiucf39tV9RLCF6pKZalA5d60yha1eHXCV0rLxtVbpNf01iOlAsSSl8Lx4nal9CT
SHi8E6UK+YA2NXcWK6i6iC+fQiztIzzu7J6phL6Dv+gbuM4dEov6IHcY/Gg8LvLHtfkn+GtHAMg6
XAqzeHLuDBAO5uo72Jm2mxTn2dZvqvh6yHuafl2y9WrbqyZU+/CiOT9oySRxKo4yZ8hbNOqqq9Si
c04MoyxSPuP3CnK7YgLJDmpbwNfsfO3pOa56E3IILaQRZ6tPgv7s6SqKN9eKZfL+TN5NaPVvGWGt
RP+p6U5611U9PTQgBBRbggESHsFkuLy9ejjKa+4YGlqQ6lw/nNlO7HfXwCFMgOedQ4dnDbc6jbCy
61lbodWgOM/lFicQCX89nJQtssb0lJrfs+TujsSRQSyxKKde7uYxlz7pNcxCra/f9nydHNk6CXgC
PgRPsNdN+MLuVWn5t10C7t2GAPgQ2tW+atY2gqBwW+xIbdhet6KRz9lyb66zPjVtucoOeGMLCgkb
HnLbbA5/a0h52+7kqQFKS7cd14CU7OfXSNpDanBqxNO5gehcthEPM0gSXpglz1PDHUnOmM5/gwPl
RR0epEKQZ/K7jjg+sQMt7UkXPaT/dJzAbkyNnqTk3wrhJQA98d0Q3zXtWFJjB0/BUbZteqcXtXla
v/rXhI9S+o29IxOyJcUXPZcrizkQLvuSR+EzJ2iQEbJgJhTkE12YbSvzpzZVU59BqoNJltov7c8O
7Pm6qZ7AKxANrXbCRI4ltgvl/nynErWuJDqU5X8PvWBet+HLmfaIhbuoB5XBu5Ez0YEtbJg03BmG
BZFiHGs6EbmxPpkLwJgHM9PQCRWUWZ5BAY/K8tqm+qJs1eH6lXCNIm/F1uiTk7yZj/v9jrxX0DMJ
MX/a3OTyCvqLUALolIfwEZh3h1Ut95DurU7IP5tPgQ6etkUNdC4wlfnaaWOCHXjbfxdTZICZnahH
HD9KulYnD3jhXmA6++AKVozAn2WaHt22PpjKhD4XIWkxwHQcma8Xlx0H/c3p+DANinQqZSfBA7kN
x+teNyrGmvGmKFZwq1G78+01nN9l+uco4PO9E6OtAMKrW8o3AkTPAlFzUmXmtu8aPPMY3UfoSJEK
pojZhg/7WBpDNHg1sdPNH+DYH8/i6ZRl/GBjTl0wY4FbbCA6me6PNN6aANZW0J7l2WE28FpsBWXp
/B/tWxbhXmc8/kSZWggb2QCjxXyYkXEW0HWdl6XI+QuH3ljId943zKkjz/jVfi3M3xcjPeBy4JU5
kJKgW7iKiz7S5lU4ixWpjQUwC5SAnwpcXJvET6bX3liQ0yPCkb4hqj/3fzqyd4X6Cp95DPR5pXfQ
90TvKBzx8HUuAV4qtc5o4D62rDcOyIudIF6LZu5+WzpWPsyDd67iNKfOfFfn0mrXykptq+Mf52tE
Dl4CClz1i+vEztjE/C+oEBo+5aUeJFx5L4bxgI64UKvGZ8rTywuQIrc/5sSTupiPD2sILnDoK+a+
4RsZeGNfQH4GRmvILWKSA7f1vNqn74u6Te9nyeozV5TwCRyDAyj1FsFeDO6fyMtAw9fh4nrXzBLt
F+i/JSym9THD85aCzt9AyuVOM2spleeSCkpopXh80ckN6il5EeQPi77WasZ4DW8k1LACWluwjTIQ
ZRYrpfHeh60ck5SE9QnzT9YvVw11Ew7Amkndpn7VmV1PyFdZ786X3KU67RNLR583V3CY4NSvTMBP
I/Y0x8gvZ6JInqbURDrJZPLJw16kwSxcmtbfyWMu4+N7kHYxeCGkH+1NYfU6UUkugxXPzTPDG7VN
hb+8ZdVr6QouKYQl3dFOpk3IEgEGqEj7mMsk6VZxAUBpEPRFS0TE8516K9zhmjgxcfhrdUHRbuwj
Z4QrSkuqp2O7HeOmTpv1esv5GLa8zEmESZr53k7WI2emmWDiYVZa0FWANc9a4X3wbViNE7aqJRfD
zi27qlA1PNNkZO9nLuga2cyrzlopjUqkx/dqiO63mSHKmbSR/IRP5udA071ulYo7nGVrPtGEgJmW
FgGn+whMvVfu8R9Go+kz0rRfrtUQUnXRJgMhPHWM8zwMgjVfugMt4zbhdqaLjHk3iU6mq/AgSk6J
hWuNnRDPRKwRdBv5vCBrW2le7ydgqN+jof1IXg/9RpHHQrBKxk/QdV7Ub8XzKKxAZ9NS9JAnIbhF
Nx1O05WB662znxUBSd3u/FEvQT40ILAwGnbjf4BDEbnqde2vq6DATsfLFF2DN1LitowAwDWjsxFS
Qzz0IO1P4T6T+mPTl/zZO5wNRkuC5FyR9VVOgKfd8hKhahOq0bOXdlD+jVlleT/Gfv/hIbH3gqrv
rqM6VfOC01IuMnOSnVX3lDtetpHSjjESD9rEWBJMt86rrVJcFVH3OUlz2FmMlipyHTVw1sLCBdWE
94Ouh9WklWbNyQ7zT7j95C2x7Ni97JykLkGl2bup0ysLSzARzTlCe99u/ZJT+sYnqclJ+27wFmlF
EFxfMVCrFLRHXJgzKDCCIBI4Nm3IMUMVHcDd4BMyBdys8sScnJk027Umc/auZ4gtBbON85v91jlX
Za81UHwyO6W2ZTjhL1AR9CWYmlHzetfPQxRdD7phkcqy0s26NL+CA/Qd47JFbmpQbxaWuSUCskhi
8dJttw4Rn7FXKJ5cDIw1TUbopxMQytnjFVGi0jdCekRcW8XsQtcofWeZXntck5TEXgf16MiY0BYn
Wl9Qodq67GFRtZf4Wlj/v1EUZ2g5CYP1M8Nm9QwH38V0yADFl5rEcCZHI4tqqhK2QFXW9oRp0JUq
JO59IAGo1+N7y6Vn7M3aaSUAkkEGWff7gtzMFJfWZAjkGfhupiXHhtoneijzz0Gy8Zbi+bJptZZC
psqRXVvUllS89xZDhuy8ytVdu1KlnjRwx6h0jxnPnSvncqNPU/YmIZ5m1C+Q1BHVbB7XpKYnO3rP
Xj/ZZ4GnenwROjk6dAByuyW+PLFBQNVC+IDGfgomu+PlgIrr8gJ+/lXr6kVFZWFTpbhmbiuVyTU6
Hiswvk/dD2bA6W00k8WvO61KXaIlDZACQp95GDMx132rH/O1H0mTwCzyYfHF+qLVtFd8QcF4ogyZ
eYLfA5fWJg8O290mFUe1Q4epf2pOMmvSq+A0fokogr51zM6bjGrBKHiKVcpntIRv1dRQKz+OiHkR
LF7/CYM8D73WB9e5PoH8RcbV5A7gxJ+FxEsV8hhGe3NRh/KN2OQaGEr3emZ7t0eOa0cphg6pd7qa
sMzLgZ9AGqof1zE8CV5elNDoq1muDu0p/16qwsVucN/xLn+9otpYT/t/Yt9DcRMH7+y+U8hR7gAz
fIxyGghYkYVtyWJC44LkL7i6JNrzrokjf606w+W3J7qt5z8bxB5L/bmoCVyX1eRNIUBoIgwNC6s2
K0NJ8ilPSQTsl+V0ypvpKK9U/xnEbrh8M25A+C6I9ZI2AK+i2HbyzDDdUzyTBWzU84oLRC/9R6jp
dt3ac4qWj7b85GSWcuwd2E84WhyPfhD/8FlFmhyBpCnTfSKjxbEe/dbBRW2mpn306zBV4qJm5EMw
r9t3JdatUAc+ZzJ/b/HCyjXW37ZPH6DIUXEaFVh/YLL1HaZBGNdTYWW7R4v7sdh+CwUguQ3wPq4O
gy1xErI8biVOF5Xb3rhooBTBG+z8d1pFtXytVpBRAUOZLgwYNQHB/6PXgjMPf6RR1cZe2qr1ATTu
6YKsoJOh9uMkZLEKrVe6E89M8jD7eA0m8Zjhdb4TPbSEwagKSOr9C/KzqYyv7dqZvvj9T725p4Is
HCIXiiIyURYxfOrKy2ShAiUDh82OfZk36A7ur00j1ullMgFRDQsVxYY/9S9UDH+VgbTR38DMTHqD
MWN29pB2Wh2qBk6T0XtpI5rP2UgpgSePeybKXWS2MQDW8r0LkpUhNxbnxxCjSOaizCA2olH2zFdu
sFQ5sDS9uwy/IP32fx1XNDilEnRX2+e5mllmkBCS4yherB8yxCx8Fu5zKF9YHWbYnTDgPCU19N+a
8larUu1dT9EUxeHvR91466ydT/3hhCRe1MIWr0ouYUpTk6crqPEmCuIpIND50MV30Fq6teLnY5gY
8x5U84Hl70vxSVUkOLyJnqb9ZpwIWTVb1nXXjokLLHArYeBJ8zHJ8PGKsGiUBicLsP/FcYJJInVg
IujNoH2WfbTIhrZ+do2fh4mk6UtEyWhuIYbNfumCNJTuI1m0dyY7QsPjIRAC0vAYgJQxXO1hK/GZ
/PfhjsBxwC1DJ/4TO+tTbXsD1+msRQ0lyaugCB6Pyfj6dxAp0IZQz9lVohs64pyc8MFFkDlXgv2a
vQo1E5GoJk1HTTl6QyoiaHla1VdAN3I36Qy4mrQZE0izjTecrkP/dLR7nMGVF31RYnsTrroV9Qzz
DHtSqdvUlK7L1CerDjFNEoQdg8FXizGVxyQ31KLtLmZ/1sIS3vt4jPFHCYikHmON5c78PtplrIUb
4kUjckykTXXqCa7Ry6R415XFT91tmO2xjyB0tjv1LggLNJx5HuzFCFOkfjeNH9+QC5p2usMneGcI
Ft5b922KPDDLD76BK8eDxtJJh9bXVTB7760gJ8EOhORJmRGtZh1G7A7iv6T1sBki8Zb7IpMrnplr
bPH1VTvox92S7F5dt/z4yK8xxf6H1H661mlV5GCSBQyLWez4j+9Hj+gL3Uy0g5HRYg4QaM0+2Dgr
XTRAKDKYGBO/G8B2Xixll1rOi5vInOCxLS7kuRQDmMJZOtvlF8hloZt+jGwAq85c2fire+Wk+WEh
jImTA2rnG27atvnph0u+czzXc7xymC9WZWM7Xoe6rGPh/itOIagvPPWuAhh8x45XlQRSfEheuvVi
6dsWVY8+Vk8lF449Z44pmfKBnx65G+xOiqrcsc9BIMPifezcUrZzC68mwB5EjCpIK2Kip44tsu/0
yeqDa3DpIffch2f/REwBrUdoPFzL671r6usAs5V3TMa6ybRlzrHDRbC+Pyu2Bftt42B1VYZ4dYd7
flNjA1hyDQXfcGQcKMhjV7+Rh0dfZdDQznKcW45APJRKLvE0PEDC8NDUjaunihZwjVjgyllz1lqn
Ahh5fweCwTlmIokmUV/+K8k4k3P1aCe9VR7i08zSW+fhEzM34EfFZcPgmRhGrWw4Qlg/DwIh1l65
7r9nwXME3N4TtrVZ8SCFQ+uwHDKKtRhsqC9gy18U2H8PsR6O+p5sOhCLDBJzPMDWaY2ofj2r8wS9
sVo93ixZDFbd2Mn1LPkVl4kEw13v9WdTZr5UpLslJV/EGMasV+oxwf3nY/yQ/qQprETWUWHXe10M
JJB8xXUI5YbFBAy7jLZV7XPnjXT2ypu2lwpr4BYVeF+wlmVf9p76MRYDhNXWEqyLgPR64OxPHL9d
x+DE8QLtS1bgd2Q77r0jhpd8Q2i7YN45eaZUXxl0ld/oghSgFsJTtQGpc2q0nXTKn3Uz3KN5Mcw7
PWUFCxdey8+34BjdCbwfH8Rvkvj7Lyq+7pBC+Bmj3IUN3IsfAslI1Csqjwz4f01qlk2GzlmAxMYo
Xvh3UOexXegUoUKOYqNIT3dcTJJvRs0ctL1M/c4OfkldQoQGbA64TUdJopRpesSppYi0k3cky7J1
pQod3EKfSHe8ek7RmYWUuC6DjbAPdNmaxIVMJla2v24lgmUKk5yC1k9jExl/sMydjeIl419nZ63j
w6+tqBdN+YT0YoCLZUtldJEuznZQyZ2UArfNbdvtIjIsMllsnE3BDdA5xgcJQzMJzqeVQS4ivAH7
R97xNU+9EqOXYT0eylO4wU6P3e/Wqu8zv2Vll7d5vfaK5LSd45yierhnO53k5zfpXyAvE1mljdyQ
KQzhWjdhBr/F/stt3gGz2coOKYM+JoP6P7VCi2GMfteyacn+LzTLOwvYH1vcFR6t6j0u5Zo2zV1x
scE4zpd/ndBHfG6hLkiIhJFgSxn5yq/hX9LGsG/lhK1ZV8qD0WEE519tzHOJAbaS2WIBNbS3AKM/
Yt5hfF8nS7SweSSQBtLR+syLJBrFifEASgB4JZmFQBhYdHQo5BpzbD2ma3scWd2OiO4k5CkuohhZ
7kWox8S9oFv5y21TOD0j9vjMcGb7a+etZfq96xqQQowQyXfU9jtS4EkZwg2oRZd1jO5v3p+GhTiR
mNE6rpteaK49DgFxsXVFffF/uwCBxteW5cr/pxR5VsK45rF6SN2/JwAVeblFer6K1boeTTgb5uEn
GnfSf8xV9VK7TiF2BiWcxW2nDaDnUjRiqeu+LADTDCvG9/WwqD3pIGjZ5TboJ2GRa/xKxzDZWf8G
6i0zpVnAbWohpgf83HYcxnQmO6R9IZnX78nhTdcKQ5/Ie20gCLJe7GLEutR9ieloQhEBu9+fb6jx
fBKuoJngQacOY1y57svRDmZH6PnF+Bcokz3EP+/cOGqw8y0grW3xf0JDr4rWTUhGHPQ+CpFcXoPx
b0G/xwjbdfffwW1w9br4O3psz1nkV0kIN9oOD7/bHfjg0DJ3VnwfaiwuvBqF1DZekUhVil/CCDXk
cdIjGdPcTCQJFle94FA/1jmwer7iK1ldapkSuNkTqixSDWQzUAHSeMLyzmDuoLTJRyDQzqyyBLVd
gP1hE6x37rvTWpHhGK2HzK4FRfSKmFhLte/v8lbypziLrINlt3qNW0PVrxfLwzyG27uoIRuUq8Ue
o/2Au1pen+hTKW+gj+citoUeNddgxRABVOxTyMU/xNGFUtMqn7Q5UKnNC7PtfJx8wJoTbL2Akov2
TGN33XEqYnTHw7kXVyos5rb1IfOPMf9BLMD0Adlo/eb/VqCMsSQxeyyzdDmDkz5FcT9tOBED2XG5
J9Ec7pWxKROjqhcPjbfS0IZl2cVV3EiKeXjt2rurNgHdhVoBGwgM5LZ47e3yzSWNP1g2o2hvDtFH
fO8d8vDSIGF+rd0cw1d031ov9OgSIt3ruOIqSnk7arfOFup+tC0NQ30XY49Cn/pSOglvaNe7ZqtX
nqm+FdJZ0GufbMVvTNFUVkoK1MYQcDsaltnFCiggUxwpczH4IP7+i2Xyi/nB8E6ZuyD5TY/BWFMi
tf7fPTTb0PynGFgBHeXLhSjCFnRbO0a81S8RzZ9YJnRlqk4Ia/cLd8zgNqZztYUCkcFHC9I97dIN
FQpdcCdX3fg7q7u+e8T4Y50bPG69f5B3d8kR25ys5satFXxdeYvS52zpw25TbiYP5Dv6Kmk6fvOv
DujBj+P7RkWydHfewo8nbVbD6/pKGCpZX2/AY0rhBTRESJVvGzB9UIULQqd4MvuNPE0sikKPzpNP
td5Qe2HlP81GeAMTSFxNFIXOsbgUvjpP46iujzwI594MW0UZWI/+ImUhNr32dMIea1PyFcWSHMXg
pG4F+DcguAuj5Z74vJJaq0Fqf7a/ED5/QFXix5YbX0WrsoucRWTe6BmOFeP+Y3FGnmnB49quBTrS
Ef1XHMRh2+frf4iTc726nfdaILm0GP8zIkXzIz5965wPey4+0Sjl3L1HD/S0L8ByTa3Oqt3CIDGl
Mq9gLsbGjKyZeNObfPJoINUPs5hoRaWAOC3NgSZFdEEm+VGNvr06M/R527v6WYICopLlGtRfkhEi
29alSYW227GduqQX5eiDK/CL6UHgRDQm+kA88+6xaIclGf8YZ4I0uwPgdw/UOhAIrzUjIixT9BEr
VFHfguj5qqWn15Qxd+xDhdZfwQf1yJHZpigafaDs9KB995Tc+9OtQCUbdj33tDwvoyNEJ+fxrvmW
MpIgfRPsssUe9OyaDb83QD+fY/esLeH9pCp+PZZIt4rpJvDhZeJfrdTO9Dr35IWpNzhWJDsH3rz5
YLTRzhrGAMW3hII7yZ6bHvL2HpaJCKilFeIAsSIZeJfGPuN2/iTz3Z1+TF7oA2gzKZB1+daSFDS2
iAGfkav1IqeDUa1FqlM0FaLNf1EEVqgyGOXJ1GkCh79S3PXqE61Qf27h8p4rrPlw4Rj9Eiuqk+Gi
rvA3yCDvVODOMdYJkx6AKWXTM5Qo6HG8eFGlT3o+iSzvWnpCjJKo8tyZqzEm3r5hXD6PxYSEw4xE
v+X/HsV8dB6JV1qYrRBMepQf568rF/JvbGMoRV1Id8CPSrVgyRS/aTnDTAsfHyTRsCzkVjyhrRXx
KcWOgQLURb2oeaYE8IlfeeZGEFJuxFFRGf3DIOg6vnIMVf0GMech8vdT6P3cDrPp9uJqfyWdn53L
QZ0SRDgHMBZJAkYzMJfPTZrFElqiL+jnEOZ6LKwOzT1Du2OiZuuHjmRZlRggEGWuLQNBkm6MSYy8
Xb6TqT3nDsUaEUTwz+RWFfuod+ERUmxORJnwGMPkXh7PKsRyZmhnNNXV64URDpeWeIBd6LcEVe/x
klFm9spw0gDotaCG83fxtRXXRbxEGDkOCLNf9oDAktDX43PhuOWuE0UL0CwOZArZk5aXu063RYRU
gl93ACgMMP/asi9gf1TY48exBuW0jU1Ltn4dI3retqtqlMaW36Ic312cb40GKnDEkb6xv6oHhh+r
/Ok+MpZlcFBYf7KDZOjwjlBeAWDl3kbVjW+pdm0ri/DBtC5Q+61iElRxpa1f+lQ/sOrOp6Vzw5zP
AMlEba59gz7AU7GsEuS4wO9IeVbrVBLsaaw5zJoGG18nSTQnQOgu9CfqIZGFl8xXuzTO0iXjhSat
RHiWlyucZWuZmFPn2dKiIlD+jy/yfDYUsroBUx+3Tb05oF5fWr6kSDfgWj8AkPvwMUSKqvqGLuDZ
dtbqXzIWJwDd8MYwmnWI55KMyDuRtAIclX4/C6Y7WS5AkVXQy7iCt7qDplXUn41OeMUtU9+hzeuJ
PRTdOWfihpn/GF+IYdDuTNifYbPpBv2XFkW48N25HI0lDDlH+7zfccSDMIND7lOdv3cVT2Q2SICC
FTFJOnWeAqfG0MXNhtOQzHeZMCCG9g5oXURR/YH+aO0YPvIhf6pcXrbZPB9bQcAMVfxZSBfwlpQe
S26P6sJPMlTxJm9id6M1gU3p3WpgiqBkvvfahnIcYlW6gre4x4L6vBvUueWm15XybeQxnz6m76DQ
+QzL4cZ1Vb8WIsHLOcRd6yExPlKpoca5Z0ZaP5VnTMuzUGFwYeqmDnCavp46ZvRjHHQklPg3vm3D
2QgDE8EJBt8onMGz5kkBZFfIpd3CUtnzNE8khvihVi2H4eR+GAd/f/4xV3aqRJNAdH9iuonp/vqC
TH1+wD6E8MHdHbkQQTtf6oitkbrWew37MXWXzTpg2fvuUdZZXT+c5m0HA/YcgkpV3BiV/cOWnmdw
tXeBSOV6VIOLZBbN2wO2c75i4WeGKyuS15AxL9yRV57M7AutrS82Qg+76yLBui8yGEj4qCiF/TvS
w6FVwRk3pOHhj9IIFp5OdcLW2r4BwlZSd2WLd40mgC95NEANcw4gkGL6IAs2U8MgPmE1ERLOmLLP
l5Cz8QK+0LK8XHd/8F8IR+1iR2umuiGCbogHXl4izDYo6/9qYLS+c90SDDgcH/vE35tk7C8ocP+R
bc2vQavn2zfFfSBV4qdKjzhYvyL3jKVCDYXssvS375FgCylEuplSnhVvE1ktl52TTdUAzNsMN8Fb
g2SivkUlxETsUSCD4l3W4auVgq7OUkoBOHv0eKv6rapVaB9T25WDdDUaHMXnz8No+PP7W28foFVZ
8OF5H440NPxoH4jo14KZua4mbcoO+TNb7rUzekB9Xgttfv/wQR38s5R3YcEN40XNMnbE3mf9sx2z
q9T6Ahf4Sdtw5w6DGXspWzxBGHExxdNLoPBRIbc9Ob8Nn56B0Zc+uveaSD229UyvNVjtH2akbJMB
bQBxVuOp+XVCoSWLhYyf48h0nzW8ARN3CZ3gMu+a1LyvyOMRK5QrAqOlG0V2elJg01GKkXb6RIjS
BA3hkZ4VeywWzd2mhIaJ3+mZ6JQZCAAoyKr7QVwBhGPt79Sf/3GUsrmBWZwffakxl+2fR1gD3IFM
6Pv42VajIaZPS4L0G8tqyEfJ3pHjBBC6TTNS0hEPWGXYV7iHr0Xcs8+6f3peG1XA7C6mLUL/e0yH
mKqZhKKrRQ3I5O/5h6wWmiVCsyk7jQM0SSUOOWVz9WBWdGJ48mgJhMXVbfJ8oY+hijtCoJSz54gz
RiZYhHgmOYDnZKm3p2+tmC+6RbpK5W6kTxvK/N+FhcN0d0nIKSzZ2L7WgB3J5VKWruBTY4vVeUsZ
xIEPAcXAfQ+InksRAVnSdx4vV9LoJFtzwCT+c0QqqUYfoeNpQs1NnMuV4pxrYSmECEJUSLBPeJ8J
0ABr4BkeyYmKJuk4TXm68eASf9ahulDByKUqMNoYTq8bWgYHXTmjYAGeSma390Qk8v7FDigWora3
Re/Zawb6TeG792bJvYCkQ8KrCuuNID5D3lJmnav0QMzVmClcpyLNJ2GtgT6Aie26XKYF2aYN5oBZ
SlNp6xCY7v8gF+7pev0SYv969u9VWmtfNCjfOiEdaKFYM+FJ/WhcNoimTi+h06aDtTuCYf+6Mxyp
g7Keu1G4EzGRvF7n+xi7HRcPh06djbbD4CPzGdDP/BduojewcnSVpUua+zqVGT19tDm9AW3MzEd8
nyhUOqirp+YkSCPpimUXszAaBfdxZKdkOxVx68ubPyuelMXX9ET5GhSeYIORco3V4ZUhfZvS0Eap
B5RW+xG7YPKndwutXc+tmiWYP0z3alnITF6uwcz4JK0cDnegELOM3FzrfuVDBoMpQCmn3Y/mLxUk
L8lCP3OjxIm7B6V8nFvbJ+e8PEiVW2xfn+Z7LHjriVYTTCmMBzufvTYHOFfxH1w8UyZpf78b8DT/
/l/xw/0DY/iyEG1UK8DB6LUe18Y/Pf95wFMHBDfVtEzL6DaYlMGPZEUvdcX1GFu6CJVzF8TbZzcc
K3XVdw2hv/N5auQRrHb8xGEd96fZNqVmoI4WrzH7LFkebZ9+g+T4xiss3HmogN0Uc2vYVCLQllGi
8Z2UeicF6zwsYx6ZbRDqbGMAboU5RqF31QgSqvN79PbMj+qBQulSgdHJYMJ2Dl4Uy8AatkwMtGEy
I9ARYsXyNuUsv/aKl06M0n60edU8CgZY936EssCYqMv7822L+05a6prfC1gOstl+rKbR8PbVnHPw
ysxwcm03PoXMrUSEOVA3CB6AdnsHWqogn8Ze/YA/AG78eqI31Yz4ppGWfFpSXKUXGRbyguj7dm0g
1s0YS00Ywjlxm7e+7/QtahL5IqCtvt78Jyjsi2Qjrh6wFKbylZKL+cVwSdlLVvWR7mSh3kw1RLEZ
lJiyx9qTNQoSvkbt2Gwk5BnJ4/LsHtqWlOjErAq7bD6Bpd1cjdjTBdttL0RGm9qiRFPiFDL7u6bz
9Z00HoCCQ4B2F7fTXkhDyNeyhBMGNunDwFblvJfBY2drzkFM3n0erehkQEILsJ57av3VWeuTsbwE
Pi1Dlx/Sb0TxHt9YdCvqDzEfFc2lRlRCO4hgUuS3FuJ1jxgKWs4qPg55suCAWl05673iY9kvV2Fa
aKcidBypkUjCvG5Ix0cNmVic4AgID/vaf4BszGs81xlAfCUJRLcOgicKhqsCxJAJB/s+Mcrz1dnx
WSmulfBTXUVKEsOfBCetW+vwDK0ClhMRdMn8bB0SBkyuLqjWPRQmUdavFCIFv2t6ZBIMK4+OFY+T
+3q1t9iuyWMU5bWq7PnIVgvMYcVO9fqpBQ5dSy6biS3XWhVgk9gmo/wRkSnjVaaHFAEDxGRuxmDu
P3V0no7uChQZkIOi0jPA5AlfDTmp/Z8OMbqxmjmjWMM2hc+364vLLwLtFP8CrueyUqmXd2SW/W4P
WR8CR7rr6Zdv+IEAl3QuPTHd5Anfxt9OO7B6KwGxJU5rakwfbbDn8llpWFgN8vbrvQ7iUpCDjUTg
FZgZaAwcUDx1sJalAD2QOzOgtr0o1bJ0cYpTrqCS4/diLgaNetJU8QEvmplWBF+ebsduvrHRNusS
4Aaaf6b8jcnfVqg/uC9+cu0kLhxkGaca3yYWGA1LY3j6Oxd0neEOL1JUC8BrSnBrQO/VCjvC7gle
9dMfT0WXZeZNWoEcElCxYvp4mabg2t692FKxGfTvGs1A7BAL5MywlvfXczkYkTt/Fn8qHsgr4brO
ZZSCCjS44z7GymRERzLeq2aW4N78e7T18VLzpc2P2yk01/2Ht3I907yvSjCbrdT/HopTmvmXKWkf
6TzTzW5qlhg9xUCRGfc/8DSiaZiSZxCRVph5flIS3yVCM5tPkjv9RANgPTBeksdjchKIu9rs6yiJ
EfqYmg+WYa6a22Ls5kmAeF3Zqkr7+/aO5mtraFxfGxfm8FyAsifcOYWv1vVvHzRzCAgooRXSuSAS
3RzbPe2eBd02rP06Mv31C/vAK6QIkrWYRCtKKBU9MWFot9X3oF8YU2kLpuqQFbIboyDdt6236ry+
xw2D8OVJSzR928Pj2BB/raCu5wf0O9RTCgojo/Yv+lMakqr6qXuyfHy5pQQxk4qjrZa7RPBU/2RT
qctUusfle+zzr8uIz8k62OMNQW9xaI4eEgCRinM8cmtMq5vmGaBNQ/eidsApHfVmIPJ8o92a/rgV
L81iUEql/N5tdIk0ZtYrrw5e+bwjR+RVc+H5BgiOenuHxgxlQKpHmLZ/HCOlHxFlhtRX7fBpkanc
o7BH4Rb0p9j3XCac+kx/wVEUKCOhZC+fJvoc8XdoeP2fxMFl95jRU9V3lX3iwu7PyneD1ZVIgDLM
qqsDfxlbMOPvQQLFV8/j/2LvJMSZKF8BBQ6HTxt+3rZrgInzNdH5XehvrbCHxrUROsqpmT5aMmTd
QYFgM/+9qKQPzA9O2EMGrmoLnzFhuadPH+jxkVgohJtm2RPNKS+ZL7+9VgfA5Z5HNyh0oqIqU5/e
2uRIvGphBN94J1v8pYyDpnV6+lkH+Mcuzopz4P8XEpRjGvzQ9syIkc4TlVpb9GqST7Wk+Zc/FCSA
zDWKVQhQ1PxBna/arWw1ggNTcKNBBu3Ko4OqMbo8UAGq4LCba2NgHTFQn0yRWEPVGPxwoeDC3wOs
L8Uh0FXTRKQcgk49ZjJ6mMp5X/RVxOSTGpvJ9FnCxq0B/Pz4GN9FirJXT9ZYl4MnCjao4aAlUPfG
KoZVEI1x/xUtlXT10Wdo9n4bDMvNCTiHX4wHIIPiPkhlOx7jgDdbNRvzoTKuu1jHlWCAmdrH36uU
4CDfb1F5erA2plGhs2keS6Ld6gw7SENBbPr7NEfUOak3X8pr8q4ibfjTwFyfMGKIa3zbbxNaHafb
JSQ3MfLmgVdxTjayLMiun0N/EsfAi5b6rN1cx7YdZbsp3wUQP9zLxZXsV9q+T/pgQn5qqYqV7Q7a
1gTQy0ehsvUz2Q74erxM4YpHM/OScln/T8acyzutlHy7x5fWbrdXwZqlQd9HrN/pyJEaEXUC6c1a
qtE3op/p0X2GGy35V6gPcv6XgReqEqrhiIfJgZjsHfKTAfWxCRBU8IG3PdIQYwwCovPQU1eY1ysw
oScVz8cw/d+g9Gg0o5xKDsdXbdyoO1xGaJn+sVEr6eFcNDENP6Soytanp2ncLyWkFLR4u/Rpr62o
EoyCCPNZYs6AcskxGKDKWorz+r83b5cFr8SBublSFA5/45Y/iHYUbwlINl1V3LiI4PXM1RgnoDyl
FfaHb4o/r5Ne+o4C6yddHtmtnEhTEcGBwfbkrI+GRkKawzmLYhZXNMSc8cjdcqaKhfEFbPe1jS3K
u7A6U7P/gez7eNz1dWADS3zXd+/bvTaE0xYaTZFkDXsSzAcRbSxwK1BPuHqLHUrOSNdeHrXWQ/NO
PwmW/pLl03IumYITtirdaqy4VnLiY1xSGC3PPJFEP2YdoGuR6KXSv80ss7sdL/PlY3zluV9TtcaI
ddqR/El9cjquUC7aelHgVQ1s5YLYorDzrRRxhLhXh5sFFYnDjsUqAzaB8a4BYMioqD2aP/uljkJn
+8ELWrqzs1awKf16UX0bDSQeQ//fWYz7I8SnhxMvsRMSlCIbqUKEXKzNH7uCY6D5lsTCxMQNH/Ls
a7H94gcG4c3+PaQ5EAhccfngh/ZbQSyrOf+KyZxcbTnxAUxK9OkQRzKsAqEddFop2lJKH3rw84u9
KWAY7U3XD8jbhcjGp2SjwrJTAFDA/X8eLLA2RnOyHV9pwXGrUFNXMf8GeC1qmIOXyOQWpyUq22N5
2Fr28rd9UCRyj/MDlnyjm17jikAxUwa4SoLUUeVaclYdDpZcG1E8aU7LhfwUpHKKY1OoDZKcqhQU
WzWrbRH/a2bmmcQ6XNn/pMhwOUQk9SzSh9p6gYImBBQ/8hRzLW+QZhdkWvu8SPSSpNv/wyqa0DZ9
NV6S/I35LPOIwhA4in7kBMs8nh6K9K9fuhzC2y7Ap5EC45T2Z2QXnxkLOWR7AHD8PbHtIq3UuUGH
zbPEyFWlC8iX1OSJTpu0tHJZDZOHJwLd/PfJpCGRJjMfiKGMKyrZvIkP+nJ2hpx9xxJIisHQzKmt
Y8gjHmH6Vh5sgCqxu1azv3zr0+O98vrOeDVdf3aPJJsevT8u3v7RCXp8iKRliR7pQqIZ5P33LOJG
a5av+vMDKbhYJg9gME0SiQAIW5cRxMgZn0jAy5+bvFnTajJ5XHmm8Vjp1Wnk063IEIifGtCU6cOF
8dpgHWLhzHbJ4wQv4eGtWxneJTivvzBPxi1I6XNOG3wb+pCEYL4+QFo7ePlmHnUZiwSAZQ6+XYM1
gOfqtu9PnOA+RwBkWPvl2RGKwRInib04QbJNEb/pk8DxOePqjMz9Rp/LDJexcdngEKGzrGCHF40G
PTcNo8fGDx4/+sNaj63HfVDlEbMI/A1mCUtuej7euEbplZCRUBWzgS+x5yphVM3I3KExGNxBVtkj
8RT/O769myyqc8PPyZNhdXXhha1YmYnjCU9h0FEfQ/POleE9QKAIoNopK3sxEbCMnNNjv6JRKEx0
hiueiXQWhYzAvQ6joLqpIFK+M6qNqUODyGMt/row3MrYNoXta7nDfEyRU0mpRRPkpI/xiXMkBDKt
LEkhbrKKKEyF+29yc2nEYye495LHzVqW/A3TOvrOMqQYK+2pW7jLzFwRX+ckxydrGwPsZduz77on
/mTuNdX984VwQb9+42mClCFa512goI39P5oI22j3XEoyto7pXjzsMw2nOZNRi2jAeEoVurL/Slc0
k1SQpRbe78fVglFr6md4SQ+vG1KlzP9vMDISLS/L54UzH90DK1UaiQyixeIxubKNgkEaiQP93xm5
Hsafdjj9u1NWo1rEN3phdkWfQiggZziCFOmJBUeXMM4MusMHjQIpTYYkdDeM43EpXue10lLivO57
R35oYbhqlUPBwQs7qfOj9QZWjvDbc3izQZdtIvEM7uI+8L5ra3/PWc89XWBdP+MdNt4dRYlfaLnY
CvQF8Y3kpwqCylwNgCb2nKLY3yOu9zIj4ZYRA2vcA8pIJ9WGgJCTwCFYA7Rkkjt+FUUVQ/kQTtIO
0/FMOFZuCNGv3oeAir0cqpIpQoXCo0MaLjAfYq1Y1kSbazqKWQPoix3SGbhsQH2Mgip6hn06Rqgb
SLRklvfcAnKA+boOU6u7jMKqGoXhi9NhOlChkCw+vQuxxWoEm9NAHHHe+3QsrpW7nUdjjSctkxxz
mPuRkZ2+rokiZJCv9Yw6BSRbzJV3YMs/apzNj5jtjSI1E9mx7N9oasHzmdoqrgnt1yT3yUbhp7Ch
5q7/Xub8j1lOYcDqs2uLBuiFZrAKORJg9Wx4KgIhj1SwFBDG5ZQzD6XjFrF75FRXwypS5tA1MywF
01ZwndkdwttZ0Hdv4Vk5rpOgUJ4ZxhfCUidFYdrXWsSz/ULC5n9A3TjzCJlZvkDPrv0MNXNah0AS
8Yv/mAtBI1Yvsu6iOpjcbLfpNvz0CKlgqUBbg9lcVa5H1iVIMHUfq2ESe7Dvaxdt1YPsyAr+SipK
1iPRLUgXkam1gm748Vs6ubVmxc4x3ZrF/tQ2kYD/UKmL00Fr0gR18CCqnEQMq/uvrBEQX5Wj5hRJ
lhWyMJmHmY5WpR3w0QSztwtT/h/6d3Px0Yo32PEI2TN092UmcgPhy5W+hpeR1FWni6oiWUPXk4Vo
5P0BjY/k0QdTiJpQmwPd+JlYBOzEbMC35KR2Jn7UMcV8yG7xftITr4uCRQTLFd8fVXQ0QVWG286B
pKM9Z86Rm462Hbwpx4MSnapRrto4alXGIm/PhyrP273RfGUncvJrUgrAoOURHY8fnRIernIIs1ss
Lq+AYeqlH3YriS7JcrbaiE9nI/tUNGSu8yL/MgEaO/gK4g7BRlsNXJ6yKPixUUIIDIUWbTmzivkl
bOQNACuiVe8HRyRtGs43FJ1wn+grOdAcFmVCBk28UwtxBontZ3Au4oY+sABvE96/742Mo0z42FqG
qdl0FCaREV9q2EBehk7n2ANUohacn92IBhVuoXBKorRXQEyUNz22DLzV/YpJ37aF6cgRLyPxOzp2
dRFUII/tRs7ditTatQ6L2vOok2DNDEsusm3X4DY3VvbzRd/Ip4CLpcW9Ks/aJo2xWpNxHfsYJIdm
L3rXIivN7KOszw8rXB98HCrhAIYk4QWxOjRWem2Djshy2ny3GPeIruzy4OM//5woUmkEQFUV9NtW
CO7CEd8UAT7m+T55MV2XAzAbPRD31JzChUkTh2y1/5RduBNSOmbz+UV61QD7baPNlPPh+TM4FGPy
/Ff5PT8p5KtVMBeD0BQxEDxqck9xk1Tr/mbDU1M1/JOM+HSmALMrOtoh+WUNUHvELyaa3Xb9Yy0B
7bk0wI31RVejW9mlbSzkt9PM2Sbq4zITB1yrjJzFfCRGMLDRhjOXkwZiNis+74HQgBcMbt9v/+VW
VHk5UpvrxxsIwxumiCWi4wBCDoJJTJrFR37w8FrekmMGtyNVz1wFMzHbbf5oJy4U7XfQ4V4lePLJ
Xy1lO6ufJGMo/eyw3Bhiu5humIB54TKe7ikiElgHIXNW3622N3SN563sFrHivE4BtL4tNnb8H7DS
m0G+f9GPPDD6SUVY+9qlbmjYOKRaX537POJDrLBwaWsqE/K9BmBNSGNnnh16H7x3jYHZ+qJ6GmTV
HU4hqihNsGvA7AYTbIqk+Cfwiwq519PY8vIaJI9JMajPn6GrxukV6RMCXpMsNj0sjjKdhPV02N/g
yZ14eP6k2lCPEtSip26I8Ya+jKX+Wezk7ZuO3WNi9uQ2zX0nZ87qJH+6SCXxjFMgRr2iVB1vEloi
iHF4wYb5mrjXKtcwvikk307VuKAhgl8fCuUko36DSBte/z3pv15MFPyMLMcJfD0aV697U61OyTLr
G3bqFp3bpGLqyq2dDiq7A+34LdSMaNCr5mAco8lcRUOkFCKyMVx9fPp7ByMcd/7S5qJFiuQvOnCj
B2UWTWPtFDZ8plDDWYurvz9NbzYGWex72qzgaNMrAyzApy8zxMnI638BYZRxANBZt3KfLOcVwSfi
tvC5n3DTGlUHw5k5Uz8kUTZ1YLcmUrp5QEdtwM4N0G1Vj5QbMt0QQqdQMZHdzSXybEOOF1KR1tfU
VK73oF/Z6RwGSNM9x42H0kklNRQ8Nf4Ewtt2Lm3GctnyNpVm/1a55iqq0zVYs4Bqm8e9wCGUDEHs
looRc18adT9Envsqp6FNeOJWnZE8nW8UKvR+rFl3zn8GvFPuAA4NjJFA1ABW/TI2E/3q42C+L6qt
r/dyMdIQRd57WATzFJXVBf9yTw8TukqFEMUDxqzweB2cw4cgaZk0QTA6qvK9u9U8QqxM685KhQZQ
P2VyQPhx83cSELZU8gT5ID8+i3Pj8HLxWCJxqyUbrQHXUxqKDQqhGoKCsfEMw8NW8wAi6GupqHP0
rLFucvOOWtS8nmhpvc5wsQTNVRdTpP3ElTrsDjeV19ej/iHNhqmmjEGLPHcujLwCBGrh0mV4izoi
22Rmw5LkKfhdKPVc1bOcGFY2DaY2d31ao+7xB4W2zZ7IXP5acdH3HIcwB0AWabygdMb4zRfIQ8uq
QEYslaoRrUBaQDu6JTNHiwQJvFFQzgzGDVADFIjUkXZ4p/9EWeCoCGGm0zC3p7bSbBdVhFI/XY/c
CPAEMqd66WN+cEWQjwwVISF7bDSYaVGqaKbt5wycgaXN9ObVZvRGR/MkhzjsbNtHZCbuLKpShVRn
onYsUeQQxhREZYkaCbtcUO5UNRhf0nS7pgAB5bxC1itWlGlaeFjvjQ7QLYtfzUPHn7k5UVonLX+c
Re1WaUnn6gWyRYajc9qnWqQWl+rUmt+VSVc2Fb9rf1vQCkxLS+F4vU8mhK2F6BhNXQObQW1+VEJP
6fghW4m2vgVYN1s6BFDh5okw0QEzzEI8bx6CpX9x6iWFwS5b8hn36ZUtaSpEPBHHvPxo+Q9RkjPg
ffCxta+Fvmgc23xg38xElYXAS/fI/kWpzsy47Hha/JNSIkKJk2w9al4AtBrx9ratkf7RQpGWlFGe
8iOzs+lnEzkDPI8m35qEFjUCg7AMGujAAZgiZXO1AygAW8eaendcTREb0qVorLGwxb26Gb0+TGJg
tYeHzgFY+/G1nlmeoalG7M8rtYx4tHo5EF9Gptb9HOd11hR508iNd8lXT8b1VoD/ekNmgW4xPhos
fbMUqAZRgNlI3bdxtqAHjtr8ftYVz0PVn+Gn/Kayy1iTtPbdzsR/XRONB0N6a7afm5u+s5lH1K5z
slje/+3d/3Tul4cnJe/+pCbVngLfDosoJJ4rbTdcro7JucFX51/+TGxrp4nVMRIroQQl6Mq4XFm0
RGAjeILw9bktLHdVU8yVTi5q3ajCxqGOGF2xHub3VPQq9Yr+URqJ+7Olx6ubupghlIj4PaknA30s
aGNCrAqzFk8kYa8zKoRgFn5GCxhALG8M4MfrYGt/cc+yYdi/Uisr3topjIHhtF952xVePDP8bj3o
5ottorutyIdVqII/xKVPYBKMv5koT7ef9FVw6nLwrSOYVy4l8PnwoNUo9SuI2+yKyHNjNRufUcFx
9sNlxbY82NMMgIq0qvjqcNry3zPVMw9+DSRyqBNJgmU5w6DzN2oOnFEqHNi5ac6s9545KVzzbr8i
vL2F6FjdLkgqrHHMKy4D6HeOh8u50fSaPXxG87pgSUO6ZryULQBLS8/M27m/1KDumr79vBu6f56s
WD66GPfvhAppDyLrgCX9xSzxCJA3trwzbu/JSk6WBBSO2ihtlt2KVyN0AHWzMXrfrgRDZHG0tiP4
4ME62UUs/noJiV0rlmnnj1LxE0nV4seg0t5c0+4Bu0l58IpoG5SFCm/Q4YoW1EoyNz3WA0AO4o/v
hZ57tJyxQdEMrmqq5bot+18QhmzXwEQCgxH+4s9D/pfUPjfhXzarh35+iL/jDXXIygJF90jkPIzc
SMT4vBbEAd6P74LKbkFdFKqFmjnEhcRmW6dV1/LZIsfaYJH1d7NQPOA8Lg8ma5P3t9L6cDMHeo+x
VOyjFYcJwHzEBaZHDgb5vJb2tR2aQKR5VxR+PZc2TM6jIxjmsRpyiJC/FAQjS7gAPxgo9JC93T2g
Tr3K86j4dL8k6vofoUiSRqjGX/k7741s96ktNeX+HLA9egHKoSWKF7qBvpNjEwULe6T8Rflz+6Au
afVRwUIJZG7ZEqWkR+4TzzcgSfvy7nkjje6KPT8oU5CcJ+1dL3ufIxMZqUCv4czRYnkVxnpu29zo
Js2ntBFgf9KCE6AfhqKdpMTrogvGCxiFyR3AzHZL1bTcKRXtHPQydi2sTW0ZKGxnPgdVfXSsVPcp
I7HRLVAM7XnnNEVpB/wEw6UmJfDVUrozugMjgl87sKmqLl4KNjsneSFmmur6d4WmVIlo3pt7DNxn
UN3PaAKQ9l96aj1oxFyPXoB3lNUMXP50QhtiEeDvIEVmpkxiMTIOzVAtKKTZgeyymelbGuvzYejG
hoVvV4cum5Mx9cmrqZJ0QjnOwSwN67r2mbGWVDxeP0uFUpk5owR+Dx7mmvfGZGE7NJigUloPu7ZQ
hYXMDwCiSl7kYgJ6TMbgZiOCUF+7BpEUWLnvNchF9SUMFB50IEP1HzFqZNIxqkNGmudBG8APAL0a
ldzyDgIEetrLlWcCeXmk3NhS9IyCR5ZWf7ztBKlBM0gp/DeHVNj4kWxCeRJ0IJdiPH1nhbbu+R4X
k3UFJVZXOCypJh7+nUPLOA7vKISswJVcFXa4FEEXWvJhzRC8E8nGgH0HVRqkjv5KCfkvusmathr0
lJtEdKEbNOHbmsat2YrhvxecDvTBsSmh/mf6HGAStAYTAKMG+yl1LnJSzrT+qj4sV70xlGqaAXd5
yRjjs1TSMs6j7LcWBGXPHNpHUpCQfljo1f0dwBJ2FdSbIa9Q7RcunRGnMr/4oLdlB+4or6dbfM1F
M+Fvylc7AICEF2141rODZ0NlT2eu+X6z/zYPofntymwLo5UjDY4QHmi4nw+FYYVR9P46Zc90OVs2
v8zfRVwPBdRemEYFk5Jo1zijyYGIZ0wBuh+F8y0FXo87xLB59AhMGvzo7g6nti1EG25rpsABmdKZ
GZc1r58az+uynIoNPc8ewNKivkLyfdgwTfvSX95L/8pR+6kTr2Yl5T/4blIJNpuS9Z7w2+cxg0j3
bqVJwBBgnh9ys79YXuUMIqZSf5JE3Nx/8Rih3Z+234Ldg3VUqYurv+naebsvDgTkUmHTeAie1DOM
CXvZ5w+Y/v8XHFiVH5MhqLyEjCOMb0xPXldySyWW7gr6mc8YCiQIw6ZGqn9aH7w1dsDylGupJcew
FP7rqxRyjpo4AWm/uvWrDIXFqQKi7U3bWcVgWylZRrWBCjX2HZ/F+Q+Xqc9Pt97C+rDhdRfi+3q5
w1aNFP148VMyLqEgAPAe8wNFqH1pb9+kUTXcqv6AP6K888FG81PSuhDqWwZe5rlvW05xYNtDuO64
Af0scahR+eyTvsw4ilQx3oaZ5DnoVMKtCoYRf5Jg2dSrEz63tbxQvx2KeXYgpq8sshihOK8NRL9I
f8d03z8qwUlN6I0ARM9bjqfGQCRi6nvB9NaJZgxkvtSs2o00+gXCf22Vw//GQLIVfkH+0R1mfmPg
XnQxjyynATn9jqEKGcGwy3i/pIW2kn/uRV08zGnIlW+Hzp7kE9kL1ZYE0bYvFimhj9XJSl65+CdR
WN0PZS+PAGKEPy376X95HS4/1T1omWgbIfFMbxMt4tXDClxc0snjKR6u5Mp8BMqJ0CzcvhjPv/Bw
KqJID43m7ZsHwTU5Yws+WYtrWfWpabs6Idslu0B6n+1E3dLZOqcgjVwzsLGjx6yS/KyhlDd7Bm3S
waU7dr5tnVavM7dzenxP92u56E1MXWBA6a7ajdKu5bntX98zkjIAX07D9lDUIFSYa5Nj558lWjjU
GtX6cy6hoiZOCpIw0GBucPmJaWvCCzXyx7jXJFS1jkExqTfSMX7JmT6gD/9DeUjOy+3nse8ZR+0f
VNPU6BAQ7iCKx5pZN3PJ0UL1kVCS1nepTZ0bsJzZZ0QyooemjypmdNyDmCf3YF2T6R9HDBte2vgu
US2UzbY1Yb1G2nQf81PjjGOmCu2vhf+MIs3CnhLluJaJElb79Kb2wPsdO3+qAaQNPjMOKA+M6M05
1nE/hf5oUpQJuh2lhYpldwTzSNsYO8rcBhnGwI4aNeWUN1XFpw2xjYDpJCiycipIg4RvzXoQj5dl
eKF5PJopmgXs31efaH0evmnC3Y7KDIp/RSMyTtRp1xNw8zwOKNq7AXfRPNnXq1snYmSHk2ocqpEw
tdVdz+1Qe28fsqUMipCVChIXqBc1fF6BvC5u9r79bvWosuMfoOBt/fRG2RhYZuWvTrc99JntxICW
AZHl4suqsJU+YHvzU96bSCFppp/+dr1i+6z+XkNHMJgKwyzcORCK0fSbC3IvZNKmh49AO47dm4SE
oW87IKSYTR34N6GugOLuIY2nz7llk2sszCcp+yBeOn0J4ugxGVq8x2SZgQ8b921eLctibUJl2EPt
RIkaSZsRxYRbTjKBe/dJkAZolaEfisQ7R+re+RHckwJxylB0MLAxs2/tz/SPrxeVpS6JnfFrrXHq
7USZHKjjnNqbUMsyTwPcpD2zVesJbKhJkUsJJX0ay/2xlJQy4obTgaukpoaayft1yp9ci4F7X3qU
Ye9P+n12Rb6eiHEEABkScQC1ftvQ3jGlEvZkpwU7983kNUY+G4apYzXYUU+O6CrjjoT9Ji7JI5bL
0HonbxdTVDyJefHVV6uJjuIRuYru9I/sWIU59OW03wsq9FDWlueFRC1f1bXN303VKNZsyuKnwZNT
kEWpMe/IY2/cz/VwtDj0Q2q5JqzFMdDWrvGo8x3YClYcIghkZhdlCzTKH+l8ZMvxmvLvPC9ejslG
8ak0ailKbwKqBqBdbtR6nIevLJyr/5t8btJ5GI0ooLO86bv8gF8kUftKn73OzT5SskWxMjN1WvfM
C6Ir3kM5Nmj+F/6Fg050089Eoe9EMNJL+XpUpCXzFpp1Ak0UcxkdeIcnt/A8UYKzQwgJ41GLZGW2
zrssjWq7oBcNKgc3dRLCOPTlfuqK/fZedchYGJjMCvZc12clQG1X78HIH0+wo1KocelE3Seg1sca
sB9U9a59f7MKxoR3rpIVpmwbrji3cE94VpsethlFXJhY8dHlZ79xj8SakZ9/dYiih5p1J4Mv6OZ5
LjsbyDxb9yP+xxzOMCa3zS+hc4q5WbPRETMgMBjqEywZUGRvKjj7477WHqB6U+lVIC+7j/zijdr3
JFKw+O/jgTvs3qsb+Wjw9JmOYlqIjgJhcJvwDMi2sRZXTOn6G/Crb/cbHV1PBJvRb+XbL4xkDdgL
ATbvWc4tG7H5/1RQZQK08RuoGLlhQtDiHTJFq7ScebxUhTaYKpRRgemdOcFHss+JXXeiH+knEHIf
YcawWV5R83x139G8BcGqs9Kxo0w3AqQJa3qOb14fdM5Gu51pZw1GlNI7ulvhZzUPkX9GBPEPJPTP
+VUeW59+9wPQp8mNSGqMkWsefKHWUD8GNoR+E9Um3Dr1XYDNUsGWPlNOb999VJQ4MnaEB4P878Lq
taJYDVhCBaQxFYkdmcLYMtajKvGctMiMbofL6OO520q6mEpvrWV84XRd/htrQHGsrbHN05udirhg
0bCGo1Uc3D5iRPUUhTiIcyDti8E4sVTBnHQ0D8CwwLb/a+pDynWS7t/s0ZaOSXHltrv1R2ZhYW8F
sCHMCp9ojNKpGqD8FKgG6YzD73sFmNqMEQ+BOV2bDBDE2kkqEOzoaOLwHGtu8wJb6Z6Qfc9KDkF0
mrz2UM9Bmd6sqXBpEX3anU8Lwvyme1g/HLwKA3xsfz1iQMKbYZQrtPxoe28jz7FJvC5FKTNOX8jg
ZdQ9AVgdMSWI76LaEm8v1loJBzejdAXNy1NXergHy91vqQ/He/NpO5HcwPkl6SKSuay4Be5f1mo3
mcJGCBLXC/9hMKMcuoNRK8q9lQwDnxMtlONxwNS2hROn5dYPzNLcC6qoOBE3mMirMNPAN4KkKQH7
rZt2cCqtRd8+oBIhb+5276gHHveb/N1bGo20lfFoM10EUTEX9VHaANOEaL9UA0oI/E8NoqIQ4cP8
1rsUb4CtPvQhj2vhZKfo7JYl4Ck0dxJvBqm4p8FRd9PIZS+znQkq9cvYjWrvaXroyTmPT7skweUm
6St9fHRvMVKjKTfsG6F4/TGKFOFFv5HLYs2LWpUJMb2Cy1ha/oJKEnckVkp/gQT4Fl4SRIRCrPd9
eBsdhGxI6zOacjeYlQ64QfA1DNqtFAiO8BR9nH+nU1T3ZSWBakXBwXj1vCKEFJqXpW615euXEhTx
aXPxWVEqF7iFCdTv0LRagZEmiNpls0SFGSbbPn3wq1IBLMJQMAJABWgdHM1bGM2XFYwRPrtBoFZq
9LO/jMGOjWQ61p4fUqzHndCugrr5R8TWiiFjiVUDu+RZpAuT3pUttrPRfdh3fVpP7K0qv/oFuw07
eZ86vPiwWwFmdWF222/AB4z+9oc9/kgYy4ZI4jFP5j59y0Nv18UcuSTZYLjkLGPiZqHvt6Y8iw9k
yBrB3uUfTCoGqKEPTQSK1yT4vB7iH7UtABMgo6xEqGWlAejIO+JMwnuRr3vX2XO9dm67iprpzYj5
HpKRqUM93onpnEyICUgY5o5LR7dRaTiVbV/mvJLWaPy5bSDYoR2MxeLOXZQqBm0bH8RnWTaefJK5
/JrKTNcIOBbcxDI/552mN/dHCIO9SPnS2rI/gA+THcRzcXWNjFEL0FYD0HDCkaJwj/M7rMaiLcOT
w6jO49JIRQydAbcFmwQCrEPJTl7oxT7hVo9KT58awBNdWyTiCo4+O+0R8tHSb2R7iKtjcOyoz97W
mYmSLUns+kLz607dnePsC6RstkyEU/icZSEpAhVTYU7BbwthdhtIEDD1qc1JVoV2N4DbwDot4nv8
W2pRxC9qDt35nmt0Cn0uMaG66hucgdOUPUYfMsNrXkA5dcZt1YLG9G8WxbosP+sk8QB/NBDJm53z
cASOgi3pcTrWT46ytwuzxBsiaVEc01hwoXgV+HwnbBqSNiF9CVQ7+8Cp+DCrxxXhyWQzIeb7TN/7
A6OMnx/kSvphYZPbEz1yWYefS6GOgMpiAmHJdgaeQexnIpWO6qCUUdyr+VYnaBS5PdsGyoP15UiT
54SaXBmC3BEWdMopj+7n+a/M4mtv4Cdtyxyv7QYQvcva8lGcmi6zK06I+O+pCxLwb9PdITVzOMt8
mzLAVZfK1XcMYuWn+GHtnCaMokQnLSsd4WmeQxSCfFzN9Ujklrwnb/e4Nx9w3jr19LvuK+s5/byO
TVtao1IDUKNOer4/OibF8m2Z0/pe/dyCQeCAWGdmOn6XUkLR8Gxduo50nnHJMCxE1IoXZI3X/Zro
3f1wZ7eVhAJMVssgbcORtQebW/h7wfbPQGzA3R3JdmovmhY0DkLiEAD4nr211lhVUxZoY8drkbKk
/jmCbfDj+YbT++Tq/FG/YbNMVgaOByOc8Nar8rh6y23WvAivrsY6WPmZPjQgosdOl6ychohc80aU
/GCDl9GcHT87qW/QG5oRLTmx+2/ihP0bhtdli5C/t83/HA0sBe0lxvqVjdMkWQpQyWr0/cKc/8LB
Qmk9uawGsfrybfmk9PNzFGruw/A9e7X5dKRwBKkjd1uV7jdubmONUEnPPjJQvkLrcMlaurkI9uKR
7BiimYXE6/EjCZmFqym8nQO70AVlagoQMJWTCgMg0o55SnAxB/586j1D+IEsYOuymA3Z8I99ZExM
rAh13+oROrzKD4+pg3H5Smg2qKLaB3XnDXfQ0M3oiHlYuBzrdMyRMva6OpqymH8bKEP9UNvM94Ft
UOB5fCXBbHfQvgnIaWwyx2ccHU8eFErYNnwWGMCpiCxrPrleZYIChJsrk6cZMeNTALh9wuW4XwIO
mOdPyehRnjf4U1MghM+17NPNhUx+HDJ/G4KO2X8GUUVFVyMDtnnnDrUjYyhPwjQKKGowE7aiiloR
OeYb7bnN/uLPO4pnlzIQfID1tisd3H6fnHaqKfmSdNfBPtgwJ8bUUa6MXWaQBPrOBpIL+QN4fftR
UpjkI2gLrTgRm0x4ziwZTr0szvBwpFlNYE12VbG+hPfyUjL6QEXylSMVrtA8puLVF74v9vHbeSNR
jycEZlajBnS6tEqX6vA8L2q9BWC8CQVpLzBnA3wmojbPu2nEEudRfYjp9xYB6bspDMsli4ac4wU6
tRWYlO8tgQeoLUvPFwpxsw4FGkwdxNPZp9KZsgpZyiqEEzsTnvWJd2g9KH9MhZuwwDZf0Rp60SZs
WbDE8L+DvRpGMLv5rrCq/6igh7jiuKEUUat+hFF0iOvzr/5WOYOGl67rKwrHboRbE4Ri0am5foeE
NBk7ML8PpcjKBcFcuMbUw7apyWT2ExWvCcMnoYx3Tql1Kmx86peJEieGjhjaxpX2PjyVGQs1m0dJ
9zJGRrB9xt+/EiUFufQVBdinZP5n7yx2Mi4d086yKyNdI6n4n0jcOgOn2PGmKJKxtu26hxc+TqmA
DPwO2FGHK8qz0GChkVoqlDJ6AAhltwh6Juvlxrw4sv3FwJTNa4ZRMHUNSB76Ol4TQ8tw8GP+uPri
2PaNPFeTsfvq+zIokF9nbvvJK1v8ijWI7QQq+brC45PsL9H3E3bnQ95c/QDCpLZRWTBDIPV8wyzk
RjdNTfmzcUNG7Ug8zATKU6SfwOt8ti7GDYVgTN06ihwjhrNtV/wreVHSgQsDAl5rQvZVx0fXvfb8
9i2S2/DJnKexjpkUJkYV7aDxJ0Jxfu2igG8h5LgOqfN2t6iq3SSHiI37bZDXdV+bfPKyhIB2HK9f
lE+WEh+CW1oL3ZQ/cKPkZSbE0zsG7ml0lfeIvPsG5dvTamdtAt93nuRpJnL4pPfMWZgbpyGz0nMI
ivtbdVA2AfId+9kp3EzISxNkQpdMdkpWr0xod/vzo4g1GR3c2oiJfCDFKMYVmLatKXCBeO7+B4K7
/1wR51Zd3inzhvh8jf2+ebJi0YmSl1njc0GsA84udtqvOZz624nugXwCTv1Wgvfn6ldqlq8dGopY
ljtu2izh4eUJRZ03Tuu0Cl5SWFpsWR1uDFuYpCzWSVlBETbdtZ8+MaV1JRyWpkSydzPbgZQkDcd8
ebh+owcoD0x9tPS4+DhJ6fH3/uFVXjwtItTtYg6dpyEH+dMyLnjocsrO0iRWwbyhLgInfY5MM5sw
2k9qK516/DqTAF71VHSqnrMsL75T0LgK4/xEDqYDsuR92V+Zsemk6XbaySBimNI18Wobg7lDW/6a
GMqKSJBJsxFgTW6RJ5afJtTooZXmZr8r8aX0TnhaeI9Ucv7Ka+PGhFZ0m8lgz22GgeMT5np+3fra
k5hJQjAyltwu96LYjn5ZI+8HwtbVHW0K64ZAjw8GC2XMv983e+PwWnQunvCcjG+rpPcCvNfh4Frn
jB9iQBI/pYSQtlF9lAhxiMqWiFnbNMtJN2DZGx8otSZZu3/Vf6TzxoNxu6zXa94WvHZ/WVcXv+MS
2YA6XjCTIelNqhO8+sGyOpEC0cy9WQcJ4CMJ8fDO1DxOmPHjWqZrBJE/dNGNR/v0NSXmi/OxpdNh
nC6IVbKpDU4mJ3WGk0cf0hMmxRwgmfq+A3uj5FheiG3ySzln/pM8VL396sZfd1eCV2W6ALFGBHsl
Hvh2Mhl9Bj4ouwpx3mL5okm6ND8IjvdkYh0LAt14rpKJ4Gvgc7M2FfA4KThc/K0O/tI8eaiwJRMW
KE1hv4cWzkb3p/A32sSK7ihf8fcfuDCAQyNgPA+DpF8lY9vDYDzmZn2W60GhLHOA8o/yMCVhtCQr
gcrkcrNbycslS5eSnYVsswDBNiPMCm3Lh2AK9c5kenUclWOiHUFe9FiXDYQVPvnBw520xk8Nv8Y4
ZqaUgQ19nIkuBR6oI7KLl5DxdM6tydG7Mr0xF+aT4Bqkmcuxn1FLYjNkmjXC/oWAU202AJjSlLxP
W9SsuAm/+hmBHZJaCDBZs9AWTWFlBGzxhZBMqIa1qOhUchqH0ypy6ylZwnrE2IKjn5sIrxiqDtFp
h85YGOvfcRI47XlTx+Xyw0vuSqc1E51wFDmp4ocIyBaSuNzOiP+vE+TbuEAcxGfdtHhz8tdcQFA4
uI77y95V0md8rOxoo3UCZB89fO55bU3n1GoWjKKy77f8URuM+s6GID5mlq8h9vEnLZ8CAWizuWQz
9isIYoXjgxqMXNV17eS0WKUld9G4dmytns1X8Z+YI/rMpTusRmt+1TZeGXY0bUWSz7KlCZ6JiPLj
jXe99WsXC5RGRuXpXTU40IaS5envz04SNSknvQSPxUfTSrTW9mfJ9TIqrQcCk+c/ufHq6LmU4S2/
NOhjwXnxLCLkt6xSlC4ndVZJUEdIpRZJrZCF0emIGQVKWqYgsrazpyyoqYI2Z7JZ44L1qP0Da1pN
Dtp7lKpvSp5N2DnOIcewxttrnv5B7f3T97k7bacBv5d+kf2b85TK/zLy+Wc5JioD7Ckq6Re6TARl
2b+PHW4El+Eb574vOdONhVNUqtCrrQCE80TiM7RWw+4ShPaa6Pq6O2ZAMG7pGe8vVmSmsetfhxtL
z31JYQNUH6d+7Zz8E4mxIuyM/kag1E7/hSdTrX/xjf2GDspsgdpeWQVZPoWAeNZupEmkXluPt8YW
+468+fR9TnN/LkmoHC2GzDKOjKiZjF2Wx4QmOX7nH5wVwwOELxXYnoOeRpuxpty8oy1zFrHPwTku
jeNt2tJPiy2yvDyrd+0C9HglPIBWSOm1Tlo+fj9R9DPmWrTIRnraYEr/v+R29hgZXq60xwJfEzuA
8dIPX4fXH3LVyYvd24sbqXJMSnHH/sGr3TdT/D4+UUjWsgNbYItiEBYugnIrBpCo1cacRQbTc6OS
IGspd8tXcBcXFIrjc9uhvrUyZYMrtfcg1TGpMedQZATupQ42JHb9k9xgRSOUjgmb/bG/Qtu5c0jU
82ykNw/m7a3gYRzDiLtP5MZemcRYmbVPrOlf1z8DyfK+94CSkXdt4xpsIUqMvMCph7RgPP0s/8uA
cJYJKSmOUzB+jD3dH2klScW3ntfPrtUBcq1H8sxP9um3sR6XAf0D1etWD61jzyAuRBcLhesoHsAC
99jWTt0E/Fb0uzYC5LaJUha1vgFM5NRskUsXA6MrC+MZCnnEL/rlpHK4nEUPrO1j1oK0desvWN2B
mdPwNPjeYZmTCPrEB5uAV2S46H7DUsI6Wqkh1FI4fCAAfDJCCqLPFZjPIEXK2ZbgeRzW9XE3w8+s
RxeLlRmVM1UD3kUN3m6oizHAvwg/phcvsASjQYq7autIHBVSBSfZdBnuWFflyu2vZB/TYZkA+NmF
l6QZ7OQQxl+cdpHDTPff0smTfZ19cuxt1mZuhVusexUnUrCsrQt6ODFgvlH1hCctTQLqLw9CqBQP
+sFMneYbE4yYcfSzpKgRCAnOGtJzlhMFY5u/QyKO/NgzNDuZFsdwihjEB7zMWiqmxR/Q4HwgVZ+g
jxFwDkZSY8tPztv79mhbFawipWYkkhLehRBRTAxj2iMwEtxi9KmNxnq9kAGw6NujQegWwhKrviO0
DkQNuWheqhTNlr6v999mvg6l3/RFO3AvG9iNBnWqraaF8TRYgXpcvI5DICCCOoR6an5euSVFHMrF
s7m6zihfGv2O5YRLFCUjmgyqnZ8sMeXBVIhuUVGceweOzho2f2n4tU/EaGZEYPnC4N9Rdxko5qKy
zBNiMlQmfKdqhjfawQXh0BTqFpuR7f/rVAoHblJjLOrDSJ+hl02ycJIhzRkAvQQ+71a230lCqkQ4
2zET4xb/2b8nDsvjUvjc9ArNWds7pXzbNWSmThUVqeqMxbovw7SnYLl2VubrKRVAVft5bXxoAGga
kpukCA1FvAwDz5VUaJlhaamZulM2LTQ7H6Z2GiZFvB90G0ozcwK8q6Uhyz8u5j1ZS9DWeGSl+8T7
AdYUZudLItZE8e7PPoXHaalCybqluEjEMPJqX2IcZtpSWQSuKPLo8fxyUfTA9NmeEyZ8sJLz/kZY
53COjBrXYoEFdTOWprd/INUeWt4P9n4WRk2Xl2b6ocb/L3u+TsQIoB3SF9Dgc/HxRVuh/mPZzSw7
FrjOhSBdjJ9oy+PbmkbY1iaDktMFqHrY8IHd49Rbf5261itTY2qk5pxTi5Oit8QL6DT/gHnIKYAZ
VX/+ESpUNwzRE5Z5tOolFfYrzG6MQDZ5C3zBNXc61nLFoNtAjD+OuTPqJvUoFFgKPqdI+vtNi6ZV
4MPX2aqMA/qPomA1m0+Y6C/KJ794DThKkbkNRauiL0zF1XohttDJtJf83Xr386d5yKcf03MyklU4
odmO3CzRslJAqFlEvNIT30KeAVSltN0EekYPsta95YCR8EvReTcNRHcCmk6jNcUBGMl8QLyRmEJy
ZQ3husTWHY5iANs4Z/J9EzaPzXIbrYmYiG0KxB/TBv+tYgBiKSDQcU1A5ALhGHYWuuuxGK/OvoAp
AXanhqUpjE5lSuB8yzZ/A2gMJj5DnyP2faWqLDl0uz63+FxEbki82dpLPn7hZiVEVyuUdbQYHmwK
qpXUghEni0z3L6FjHc031zrVpyagCkIB1a0mc+HtIFFqsVNHX6umRQrT8b96AiFREvYjRCYoFLEi
rIeVSsc3qOtV4hAcmpiKn3EcQG9OHkhj9fbEml9lG62ErbxiJ5Et5YVf3QJtqy48LFHYbE/LNa0D
02Lky0+lfW1lKxBjRD7woSBjfNbDWQeCm4bS6q5bdyUHWtqs3qX9u9mHIPjlC0+8IxltK/KPqCUj
SseDwOadLkOSKJ37tA1hJAry+Y6WVdF0SU6ulBBp84rUkJe5dawJLu1ghEkg7bBTcnLj/hmUeCyC
roqfoUafpqV7A/yIHKX4eaz0isiOz01fYBgKx4ZcADW5zkAEiNcxYZUPC7qft8nJX1DGxURFyT56
WhjRd3Ca9YQPZcgtfH9gav5geQRjOtqufsOVdpEooofYipT84WWErCNJ1bkytIyv4Ap0X+DdWSQL
OtLvHiT6Ph2X/VGmrS+dd9Yu2gGkn1L0kHjVNqAIBy5flfXzHxyWVEcfwz9hdk43Yv64Nqna45qs
nRHKi7efwxnxnlwT0mDU+Q4amwCpD4cDq/c/mid9eKwlPIQil89LrpLpO51PXE3xztD74jdyu8th
U19KylF5hF+JO/kODC/yAUzPpquApxRolQOCUSTCbXdECOEPr42X3gAlCjQ70p1/HSAKJMqT5n/Y
+gBpWEhnYEiAD36dniilstgBVL5wup5L9QhVS0g8UN6ilo6aKca03/Ts4BKADDEMOTIJmDTPRLA0
WVPtEre8GCql6tmXW630+V7YTDo235Uzxcd6deOKULKFsGaoEL/eY8KfWK1mQEPBcIKpTC5rbmn3
MSS8kxJLrfAtBq62kPDs0JXFxnYrLxuWJP/squn09zIgGHopnwy5G5vb/Y3cRxsEtJRxdBzG3YkH
3kqSE4jfCmyvKdicuaqyVz8p9p/6mReCQ5jlgR8czuGxT/1H04Sc6NqtJAyL4gGzZp47Zj2xUYtU
++i0WkCQEoG1Ba64GPBkqbYWQSI68J3mZFzEFt32UzREW3KgOM7zwN5eAmXJBbA94VMs12R16ubc
XYt/5x2vTaIsgcyIHdsEBFGGNGwNuD2KlViVcfoQnuAir6taBOph2GvHcdB9YQYXSQsDzT3JFtd6
LEBQdvWCguSKmF08REsvg6uQ1eSik6vQZqMaSHyfdRW1Fet7Rv2U3THQZ+5VEhBbXlG/YsmR+sNK
dGYcpJ7XE7ef8EOO3bknnjhYnNOxcXzb/87eB3DKW2Jjt2tjElrvdeHV+maLiP7LoIV9Vdi3fAq/
7l6df3CDPfiAl3FNkGDr89F2Rg/ianWCDHm3xk11DDJueiKpdXLfbuB9IahC6NZMJFrGRJU3+pLq
6CpfwR8Q8uBW5zFSoSkbqR932GR3n+SuMg2bl124Dgm9qtFFLQFxGWZpn+hHUw9amnH8smQKswt7
HrySDPXgbPXZzHQj1xeSXj1OnEpFuIj6XvHSGCdyTXSmAeKAx1OlanOaOnsFVnBES7gpKDp5XzdA
GysKIXBr1acRgDJLFzgoomupog+HKJ+MafKIUJ+QBDpTe83jhMjObDpJTx8j3+CfJYXZ8J+dk89A
DXrLxcr4Gi04BmvAQ7rlCBolbg/AoIbgD2dKi+oBfnhKXQYbNojKlzZr6JPvlhdvY0FmalyY1tyE
dATfV7GaTznlx47BVYytxb1WvRe7Q35ZcPJbgXckylsCDWgSWHHQ8DVWUZM2iKAyipP6OYZiXIki
dTtu/ZC2B99F3K2gE/6seN3zzwbsNkMh/EPoWkyBPmWWuDlwY8SOuHdoCgbAOKpDzndEGvwE7WZJ
Ze4bnZvwChlbZ4gefPfwpqGun4EMmAHOgiAoUcJYj4lFKEFwXdxQ0MxXsZL4CznfBP0nwWONuI9s
CjEuqz3eUhXyyYfyrRJ/WLTc5SPqHYWx+SlwJXZf40Hb+I3lPDvaJHCFBX3Bgv0n5AXA+JLnHlMB
S2pFMGG+Ra5utN68p2PaabxMhJjJDGQ5ZKE1TpvOMaQOPzw/CFCjneWReA4N4hXR4aSDXP//jZo9
RumtG8DK5/KJMCpuFhGjLdxh+OTJ94yBJaUwC/CGwQKPBajIzm8HragWm9nxSOzdqFTcHNHYbUc4
AraWIx1u2Ne05hweEFq7bdo8flDbbkot9nIQyOCZY5UHwWc4pcxRmOwid1MLza3k5AaC43IdHJJG
dKHuQfby12iChFfL2j2YIN/uSv6f5Bfp9jflXrUk9zfWFu89gwaKz9KoROh+Bn2l5qvqmT+iePTi
W1oYFm/Sc/TCIb15giucHGUqt/fCsuzb0rj2dCBLDZtI3Zee1A1/hDN2pfyoYx+gG5VXA+x8nYnJ
8TBqsqUUxYPUU5KXWBKFvfwbQ4XWwEe7MPLL7ZuTThcPZpRqduODLXWvvcLDlctQVHA3E5gFeGGw
HPTKt88EpClTbOwMBN8N+anJH56Pi/5wPQap2g/muXLiBONVqtipdc79rXu4qwdxNYT9sDNaGRXD
1yzQWoyPXhWw6uILxa3Px5XOT1D+vkrasb88oA+EJuoHUgJMU6Tgt7j7nQaFsKvoJQiKUU4IL4pZ
t6Ml9QXoyjXTYtXPhmZuMSdiWN4vcbFbDeCOCglSt8e46YRdnaWeT0Fe/fB+fCr1BH3KyDoILrSq
FDMkvEnAc5MpA9EKfrTHkTsDz1wsyG6TvGXohTAivuHe5X70O2WQI3/xFH2JLDMUEIZ6unwnhnba
1wy4QIxE57N+9j4vVfH2xDz5RhLh2LUsCptS7nez4kwB0QjkhUbEDE5L2vxRUT9bFmjGtabE70CA
3Gm6DYa7y1g05Yz8xK9ZfT0nPYeGFNFGFreNSA3l47itei9IGstM+040MBghe6+JGYTxeeMDxtKs
yWqyKKDXFqGkMGz5VeWeRs9xyCwn8BKZTigmAeagL4fTHpIHyYKSDBF66m+p9Jmlxhiv17mtoFsY
iiWx5f3p/ag1yK436uYTuft6US8r8P2z0t3PTNs+2qJ7xa+78aD5I4OWD7YGvgWDSiY3cf1krsSc
cM3sE/Ii6huaI+C+a8OOvGityY2Xgpty4ji8YU6CmEoCiDvZ6wagRFNRdj4Tb46M+1ztYZOccg0r
fAtRsVFOtBq5tx79xR4a3EMH7EhhyNxcXN9DXroLXndIAsBhPrfJJFt+ztS5jpeiCOXeWK1KixUU
cfmeSlvfF5LIsCcMZFbTvkzYsE/mIM1bWKrHqTT14g66QBLrHrkWLLKYQigpqSafaaqy+cjU3HGt
QKpSWBBqEY+RRyOsGLV2y9ve9vdUDHajRIHcQa9r/ObZeuEwiEj/h4RKIutPbfDgaUEmHhibc0Dp
MSK/pvQihou4cUi4roLfsDqyBYJVn3uJsJe7l5s7uRMQ09z5o9VEUsZkPAPVtiseitMFo86fEtYK
Zpj6Jaq59/MvySUh4OeqTcLfC1acVIwVr5KWEZnbsyyYvia47d33yDKt8stMthcfJMROhnb/tZr2
JG5ckeZ/15JY3vLhE7EDtbHZrwRaWpWBNhVNnW5i9DEbeuCuXfreZ9puynOt0X7NBYNFci3m/IQt
UmumbNkwtqQr4TlkJJ/mCXRgXWscgjYHYh1h1LcCA5WYX23t0PEkUPRF0MbO+oCMoHgncd8I1oMg
vU/50S5fUvNsV83zcAntq3wWUrWCxObSocFpwUEiQspNAHA05zcetTYaJ0rwwG2uhYkgsUb86nbH
mWZyMBLQMR1gBSSzuGPCqEtGfV1ksDJfZszjrmg1S541w7DuUN6UNoHvrbvqe66LwAYSh10LnBlm
KceDHjM89w2Dv5yIkgIZT5wdKrKHe0LVvJznABi4ZkCsmue3tFrpU7IBOtbaidzfXILrpLA1oQ68
MMNxGmxEucv/G6Pb8RtcYhLAvXi0o7j8MFwCWJFLrXc2l1ZX8kwLdvME8JvkcXqInEurfdyBVo5D
5Ha4K8DK+Drm26JV509AGlblje6FRhThznV4KfikSxx38mDnh5e0VFK56aacH31m+rTTOhtZ76Iq
mj6a3Y7i3JDZJvtu4csr/o1VczkNaj9if/LDCsn5XyGKeB65pTyt5TsR0NObQwn9uqIUljzjPQ/v
8GSu2iMNq1sPm98tBjbJGldcmWa9kDRvo4pMCb9vbSITzWzr2wX3Zn1mB83KqKekoDnC9q3OBTw5
b99pvFMiyRlmPDDr1IZJIcx6y+AEh8OKno1Lb55ErfID+dSIwAxk9Dq1s+ePnyt2OoqymRm4PMNW
Il15GhDXh1NfOU80E8GRtaWLnp2nUass5TiFZmIfVy96PdRKhNAw2jjscXsH2vJlszOI2TFw68mz
qvzxmS6uF4OJZIYuecPp8sgBcTJ7pSxn6JSJlpLPOvjxS7icG+wl7bXvKYohadrE4o6ZtjRuZimT
q/0fMBMwVs3aPU8KCR3hK13nTVMKocyIzGRJlXbOujr+RF1swtxgsXc8mMlMdhTUZFhi/RLUa2lX
IX6paFsCa7AejN+7SGgR7B/s620Z5mGcdOASHHK8wzyMPkHqc5XiIjYfD7Zuj7vp3YA3fwkc8oeQ
//JcnByMnjGgKnPajRS9wzDkb69+i4OngT0JrvmGjr19m1lSjae/oYLB1OuT5+eKLcmgG3y+ie3N
FylmXLgYpuCjg4DwhbS3Bx6Wr12QAAh4LPAcmDk6bWV7Rsg0TAWlc1ehd2SPyhHZRh7junoGC25K
lqjKXzaFy2P49YLJgBMt1g9xcpwS92ZMtR6yphV/MW3fy5q/CQmM4T0OQJ3juwJptt0vqN/JVDD0
WMHqBvQ1Jw9z7Uuny9y1oiNSoQdCx5tc4+vTDlwLAnt7n5nu1l1flFyZ7Der4XMDiUDkfcm4XlBR
PPsUNKEkdOI3vkKUsp4RAY8a20DSD2/o/N+DK6mT7Zrd8HtKQzJdcGPE+s6u6NQo1F4ecgJNLZXf
bkTGIWya40X8gDCfkYhDAHgl1hzj1AExzhHEz1UL1KnMs8c6374sYl56Yx2l8m8kfGzZKdwOplN8
u/Zh9oo7O2NVpNymOQp60f039QLRgTj9KMHDP1djB+nkAajSbZ42tYXpcrzHyK6wPrfcP6y7r9jV
/oThOwgXY3qywOCQxQUaJQtJTDa2CPsomGmjc/mZwBPLHxYvVqtTxMDh6dM/1eloNFOcC50Fx71Z
z1rvdXee1ipP+SFP8XuXLaZaNPx3InJHLcgPPtQb8uGB2BPxW2xvgln+VXvzOZp1T1E7Fy02kyrs
ttvozF91vlcELYS8M7oGHwZ3X8a9gFW5lv7jL1EfuT4aEPHCR7C6Th6NtRGYkDSf22YbS41ndzRK
CA+SIas/nwJlNEJsfWL5lDg19wfXZFCZ4Z6DzDDJ5L27aKgCTaVamtgfOoN4vr96eq0+STriBem6
qtpfc+VF8s+066a4IP4H1b8FUFuuMZrafGlYXxjtKTkS1AOmLWWV6TY61xua+AC5aQ/MHUjE+4Wf
DsQL1bLcUigwILz0rEEfV6qTEuGjmbnzZdTd2l6huFjSc2PJ+LEWF3Aur7RS7E7gLP6EeDZlsX9w
Lk4abhbC/xJw1iGaTSz9Ylwsvl9UzI/yDylLx1NQFdsRPbg2pNx3irYgUSU65CDlLdtMkz8SHG7H
KBK8OIKqHcoRvGADrg69ShIAr3tuUrIYTF4hsJSQyk85NBbrNCH3R9TQeO8+E6c+OW/KyUbXSBnU
xqIBb9803lqOXLsvUzB4c3SnFmiEvYq2CTJZGJkdLI7YiRVqqQUvS30o3lB4AVef+00T2fxMTEC9
9P8xXRitqFZdyAKZi19nIiUZz7YDnawyjWDRwE4IoDIAT1rVcTQbF5aCpYnvp3T2YQbuT1KRChMk
zikYDrywKG1lpsAbiFRotW9IJQ+edb/WcwapUzrAUIduDdurl7UHGy8aZEPKjMLeGn14SQY7ds76
foZGDTU/gj3aH02Esk4pKloCteTwWMO7Vse4+zm2IYhxdV/Nfszo41CMYwt3k/JZZPNCsiCJ+gk6
OEAoccog4q4Vp7QBRjrguFPJdo1/gEZExnliGNkbiBUOb9lOzdPE7hr/+YLwn0OBJvhhC1atqfBC
Rzx7WTSrLnaRHxbYwxdTweNW8dYQ/j1egsS3rd36apvrwktKsOLJbf79WXr+OKM8evLpXvEsELG9
3wT1I0e+7tfup54P1TPlNaesOAykQl5X7NpBSxVBjr7k7Dp5xGKGcyz4bfJjrvhaP45mu7XMxatt
/jgqJRDZpfx+uZmOXtkejzkZskDmz+Vb36ooECi7UDY3Bk8sDVeRV0VSUhGWo8R5nrnB+hOTUmGT
w/i/KCUaAUs2XpomVLxdRnUFWQJRqzBBugOVKieu5ktC/nT8t+vg0JHfffJn2r1cwK8F3dxnjdbO
60dqnE8tpNIPBmW98hkz0al5po0Q23hanS7Cll0VDJfof0ozS9SSCdqnFG+xHu19uFbgZ0WI5y7m
LyWp1RLhELurHBQkQisiwoUKlJSMiC3fl40bhA7ad+hAr/G7La6AMGu123GXEr76Q06/UbSqDhwk
TSLzXH5W892SG52OvSpI7dpHgsVlSroUe0w1WnjQhM+CZtZHEKkUlvq5f2ZIzmrRrYJCHudDJn/l
m/k/cE23xjS/UGwItaLnI4tJRlMMMfGRC4uk35yZqzDoQaiesd+KUZhug2w6o+adIFLYC+M/gcVg
cgs57E7LhepQ7SOccj+eum9A2xQi94SvTsUONPpZBujw1bENL2aZN9owgak6lXsi1Wx/CmlcNI9m
hwzLf65CtRJtGnlmV+q0fqBqGOCZYTtQy6QrKjNBuO+NsHSi1BiwOLFO5J8ByNuz26FqxK4qdEaL
KzJhi2kkqtQF1Rlpz4bLmlOQ9ii/zq6dTVieDTzCCYwUtwjW/7saQhpBunIW/Dvkts6AaeMb/XZ4
q484cm6ppmi4XqdCVHw7YDDrb1FflX/Ha7+r15bZ1Km+cpOJ5/t6ahtqq/b1YOp0/oKgfwd7w6TO
Rw5BbjWrkeqONGPmF60WxmyHSHFxDaPADqA71F4+Jl0MWn/adadZdVjHuhHBoMZiXhuYfM3+5pSH
byd+nAV8juUkUqVZ6lS6D5Fqw0ecTNdQ5UjvDmn4B1qAh1XW7UDMkZcHH3yoJm6xpkNJFPzXuT0c
bJWBO6nVFSGeSB382swDpHwf9EtUF4bQ5P3kW0I8Nas8g0lMqF9J8xkdwb17/wML2Kl6C8Gyt3Q1
0JZwmnR/pB+nXoBzwUJXS8Leqt3E6E/mkZ9X4JcJn09G3mO5oV13wfMixvZZyTtvH9Efnwroaqc8
aXS621gFvlFYEVGHJs0/U0lDNh4xB/Bo2TXqkWCd1SCaVSX6atOwrdDhaqhUditZPGDFIUqUUeKw
vfHwWjuiCTyuGqHb7IHGV6dMJ+IhJvM81RDCl2oOeVtpaSxcW/OMyV152pW9tQw3Uyo5S5nuRhe2
FPBvBshpRdjYltXxg/frPOrxaBz+2XYHmhx9tiGzFCQZMJOR4QjdSw1/xolQx01GbUDViitSLYRZ
GcD0q3plr680zT27o+3slenWYg1/HhWorBnTeXFn1smbhN/IGdZvMCb0a418lzfL01r8RrWW9sQC
wrrlMbKK7ibS8gM9LTrfAGBgcpBAj5HI51zsnDIFit0yfzxcwdhzFs8a0sEJSGnU3QSrGeyp6QnQ
XneXvM7P9ccBW0JYYVGF7AFh4uNBv7HtXslgCcim2oYpfqWv/9XzlRz61P6dQR8XweAA7XegqChf
p0+0RmQKv18VLDoyfCp9fEkMh5qLDK8vJiQJhA2gVbp8+EgoWLvnaKKN9l/2ow7cHG/oQWKxA4Ek
86UYqAe5duAqklLM6anNnMVhqE58Et7auVt5DO9QFAHaCxYwyQXhodSF+tTpUIN620kAvDJwxdr8
RwRoimUMNtoFFsvQKgJEpQZ315Wdt6FIa01jokZKL7VW5Hnht0tIatcO2RHkNIfY3jGJ9kh0bMpO
YfQOa6xH56WvrFJ/gxjDLq1u1dnGmBZre+FaLegyaenFSYLQktOWMLeQ+benklTtjasZYjt+78Ka
arOOSh0CKRsVuyGM6VnoHafwggLLPYUxVQfjqy2CNbdZMyymHlYzFmq9hEc3KPKt+haIWEHrzztf
/SLYrUebTyo/a9xfPp54e/z9HObJ8VshFuV4H4Zx3kyiHmvQVkTwHvTIbyIJPEU1OSXVAqBJ4oa9
8eJ/bmSscvFrdsNTYp7jxoj1CJFX/zg7dFYnUxEIBzT0AChrcRVCaMpuGPvBU5ku9EsGy7TCtn27
T0A2D95dN41Al6B2pcMzBVSArzfGyuOLP/owk/H0LIRSGwr/YBWXuMiPQsNIBEFwp3tbTGw0FmMf
0aU4I/LRmgQ0wps7kXUyczdqcAHvy9PjGHBEZZKpk5FlP/zTQNNLni/ooqvLqCssECc0gRpux5gb
PAp9xSV9e25ubSIlZRRMOQL4t622Qov86OtHnnhXGFQZroSgHtalTMMzuwZsnisNX9qnqckJtgiw
wCgWVRDBoGcoPdnpswZGAPLmbYfZDYsdh/c2HOw7bXuQQvTaNhAIBK2lBj9NqDn7hVVL0qTWsMs5
XK1qItIUhhaWQEyt61kwPvQ0A/KF9YfIJ8W/wrqY0OAm/ksKZHhHJwKehD2fJIyY5luGLPPCA+XC
xPOHYUFGHl4MhgCb3iFI8WV3nIhXl1oqM+h18pyZOO8nBCNA3lzWEo+t6qTWUMhlioV06x2oLwJp
Vut15+/VE/1DheSLHeEER4ErX/m5M0I8R3TqZ09VbdpGj2aOV9zdl1ozE/WIFPN7IKDZtnSpI+FZ
9sUTlH0xQTFnQBBunCgZm7W+hqePq8Cl2ZRqV1gXiRmGs/JnQC9A7lXBClXCNHIHXPUkyCGjgAnM
wgvBwdCd90MPfSyy8YVM2PTh1k1YIlAz7Jgb8QTxJ30Cq8CV3DlwDer/BvFmEVZDJePJRLq3N/pw
PBJHytSaXHJAOwuQzYcyb2TURjHY/YvcpRDf3PMRIg4eIpRn3jU2bH/iRbbp1LP3I9sxG6MpWmxS
OEFGb822G2NsenYbteOqtNk6IGfT8uCm1iqczxp99AeUzv0iVx4xo+WhslJSzDr6mesKB7wZOmFQ
0dzmKIBslDZcA5VTdGUpuCzsFscyc51gjGXVyTV3RTr8+8pLVbKg0gt8PE6tSeMSOrIOA+3zS69K
J0MSjr1Rdx978qHETxLQfAI33kd65PwDYInEg6i2ch7V0zwpSsTQdoIB7DgDg1YWYvNBXLrEfOjh
6V9yMwphn4IHJ7n1ADXOGtd6nYAgLyxbB4ICmjhiCe5Zn3208fwytoBczrijho9i1b915qo8ZGbk
4xZ5MktDv+iaLNQMGifs/yJOc9a3OC/AwFruZbFnTQrDK1dTMSWJgbHc1bbmlhL0HBY0rPTTw3vD
HPVBKJMmf2Uk/vFMDhFem2iFLd+tgShXu7jKjiauqw4SOkY72nFXx7y+fFELU5FSe164bKM/eSTp
hGsy+q/jifhBTz1oF7g+YB5epxoDfoilcYJvT/wYqTmAbFIBPVk6pGjhlj0AGbY7pVQCnGJ+figo
XWnZyIWkwfETRNcD8Vrn4q4y4nP64p7nhWgsy/Z8YG8YHHNnN5fYFyha/dMf5RANfwuypgiiBRJo
xgH2O6ubg1yRnLj1i50Bl0jh4veGmt20jLRk0xtdyqcEHngVJOhlUEY/rWCHXhOl6koWQ+nvpFje
ZgIa3QTsKsRqhsV9zKSBWnFqdVPv7WUpRQ3Zt/cMh4VMil1N1jU9weWbwrLmfXXtTmzwS9ECmiyf
uqPxdQ8tJnFJl4lgW9rl3NhHw61E/QyIQmbVXX+LHB5kJUYCQXEO1Jhcg00bYXGW1OdlQ/B9S5+h
ewF4yyv/U+TTBMe8WxV0a858WVrDIjZvuZeUIiaAa2ctfj0/0Vux23V5mIGaEFq+i8uUQXLHQqCM
2Z3EZqz0uhuip+31Z5EKBreu7nz1IE/T1w8ZKPmOYELShNf+fZDEeLLB2o/Bd5UeZ/Bi0o1VIzJH
okfBjfqvJ9td2ePxhjgxb9YbfxuOBcciEyc8nuo5j9OfrimKgwa5TSIJMo2yjFRvxRRhue7fEoXw
+MLNXivETh3Aefc8qIiCMQxZcApxORaDZ8/c9KdffQuIu+a+pDJZ/R4yOd7MTFYiQM88TgtpQ/eV
Xd3788VXxtkrzoWvKRJsFcvbJM1irhZnbz1RnpSdTJCdx2Q4ZCIvPWn/xYsYhApkEoR7JeNSwfxh
00wmkJ9hMeRwP9jvojqSDX3pnV2xHx9w8M3BQ4JGJzBXJCVfskJfK18OnIiQ4NzpTfoWjCtaTRMH
5ZE4Q9R1GrDOlBDPH1jA5uP+AQhneMoEOfFnlavxDYbjcer999pE+HHsZh7tnCVcisPxrLY0UGT7
2O0dPjm/p1O2ijp80q+oYsSTiM2fAN2se/Go51hvAjfbaYb3L+VtQuQ4NiHGME0gxqJtgC4WVCbD
/wewpvlidrTnk3LlhFa6mrOYPaKSCE+upYlGTWb494nCmfGjQGhep/svpmlS3AQTPKYkRAU8oAXm
1pW7SwkinH1KZ/GVOYEcUfnxxi+KZDlj0Cn56OkoO9kGiGBukUkAnMnxJxIiOLSaScNE0Z+YPezY
CmkGihgFz9rAIGjE9ZO86d9VSv9mtqQM9en3MULzJ6AaBMOzuqLUbSd9Twj4ZI7cnOs3aXrYrs5v
I2z05jJjd85jMOP7EW6BOdYJdlZW57q4WULFYOyB7VQd3wsYdBS2yrnQ88qekQsiLnZ9Au8rkP/E
BZ4U7nLAUEaJDvPLAdWw8X7ZMALIu7e29D7C/WoJiFdffDAI6BXXcDUIWmftsEh6QlwSYd0c9rch
xEL7ZqBDGOwkWHuYnPst59TWYuoTN2+vlit6akBP/F8yosi8IENXpOUvGkxMRfM0uphBoOnvfMGg
GolEaSM1MC2hJZrdLwoq8ic/Copx4eQGrJkeYaATsLTmR8oC87knptRB4sUdICF7RlAmDg6lYDwK
k4KJMmsJMe9P7YjcmbVAPQjNp6lSHgtSIGgZpkJXewRft1iKe6jXruvnCKrbvUb6uPT0IXPAAsOG
kzayOFrOxVO5MupeWgfx3idI9ZQnstulbU5Oqkb3I6OpCaaHkM7mdPGg8Ln/MKu/nYnQxXAn94XI
JvmwW8FsXsU1CjY9Ge/qvRbdAOXpje940lM5f/WIgqTdr7djVWSuJMz3FhQzAK826GfVlWzZ4a5N
4/z4/TUJZIXW6D4c3dfUoKwxnWsa0U0WSIX99vSsEt/M8Fc1p3yPxYYu17CSnYI3sC0xiBWCfDi8
JuIYOgjx4ZuxqJNkIzkYs83neHuS4TvsBrACEmQbu/vlgO8KsBbJWCCY44fOT40oPLg8PnwCylf0
nPhTrcq0oVyP9uqNfvtEQQ39Lxf5UFUYzFrcXZqLKvFSj9ECdP+RplMIIbPaUTuQ6YtWLrdOXTrI
Y7JJiqdx4M5KCRdwEGlYVT2hw4q4CPpCO3l0qLgUobI9O6FNn5XR4/LOdq9/Gn06+soyK9HoQwAu
TKioSPBVZthzGi9SyY9Yd3fCjOZgkNxUaVg9rfqgi6RGkrx2zN8bSLMmsL6T6iWWafDLoTvDgqWW
JQRhRfUsKrUqyGPxD3TNKy6jCCoZlXm0+tk8maQJIXjjg/vVT7CRaXLfziGOFJeWtUqjBZoudLEX
w+TCzhz8hum/apASns+ObSGgXZWTUbWoQLnT6Wz4xbFS9WlKOCCvPOMrMovANDk2+dlu9rG8lzQp
+lhyQBfz4qKpltVHUy4djqAlQXz0me9isXcPaYK/GWpDyvpxBLBpQKiuW4V3JRkFXiG+qbynr7p2
JZKbWMcaL6/kba06kr0zPpnkGyoKgqJczxjv2V3aRIVXZa2Ta8wq+efMy1hZ0k/oGW7dzMUgPkhq
CYX6gAvq6qvnCuZdrqm4hQ2BzmU32MRYb9rX7e3QGL5THr4qK53drthVuJkuKUFLgSUOeCyCTYjL
0Nxfebgs2kt8olbeiVhUSkljOdNeEKYrAc8fiAB6B3ttZwrD4yIOLzD8CrGqtu2RQplMCWVRbl5J
CL2mOS5rzZDMgAtka7LeRw/nmF/jBCdKD4KsZ4WGcsIAdmJ4rUvtdHpTF+Oy/hx+zpxxfwH+HksB
EmcsNpJXt31ip1IRCxTslwr044cKfjhvaUuMc3VmYRe9HhZedbtet/hJEVCRDc96j1uoaoVEIDtI
BEBnxWpxQFCMsOKEF28b+t+lvZzxxDF81mC65mqtH0NEB+6bJrE5K4QE1WrW1dnjaU3uJQvaE7tU
G1PmeAfwfZGvzl2SLWYctMPQqBoFAbTCqTP919bDXiNxEi9u6hp+5lY4CVZK56BfK3dhtmnH/Fb+
XPxQ/9vi0jV3KwXbOrUw3VyFJrTmgBBWUAw2Mjdzc/oz76pFSTlRt70uHkZeRsnE0GD/HeuSLwSw
3+JBRq2jSBYmVdVwZcSCP1FQxurdrlOOVxxyl86r2R8ufZ6079qmhUNGJNW+3gzF7VOfjNrBjA4c
KtgW8FvQGsoP+5pbDp7WN5cOIejTs6QMedNGfnul7/3MLdo1/q0KPsll1uWtdsGRFbto26dyvz6H
f05SfC7+xpHc1jhLyDnpZNTtTC+d2Omp7dtPV2mRqaTrDvzsGNKZyzApSy6/JjmJBvPz5F9A67f2
St5W7KqUp7BtdCriq6c3xkq7I3NVOaSafrZ8s+bAQr1j/AhZSbnm+QUy1K9QjyiPiYXgiUjutdg/
nrjFxtiUMp4xbfSMQC1bPkYWoSw4t1GQyQXV0Pr2SDuTvBiQ++CY0y+WQKmVsOjBeFNJMNXWsu1J
54QCE5eUXCm/ERwXJyxhtZTjHzAHfk9QhIgbLAg7Wl4pk3SkPFmFgKkmu1nI1OIVshI2zixPB2oU
I/DLhcPOHC2mSnvOCYGoJxKOKNaYGbSwGlRi0xq8sMdCYyWTIqpKBr1hUNV48/WGJkKL6+919N4B
8bIZz8PzdccAdIPyL7QWeuLWOsRbUcWedrGvYYYGzK8lRroyA5NorVFLfLMOr7jb+EQFGDaNC8dH
hnYR1DqkEIhWivLGfiMDXM3gylNUe7ARG7fSNRQot5buGD6RdQDIf5AbfS3KR4hwQmDLXvGWCqEr
ktJw+reshiPtwshBXb+mfDwTgjtBUcB0FJmGG/cN/ul+zfnbyKSpw5o55dqhlxySJUckh49oT0Tu
CujWjazfEe+0Z9LRHBnCQHuo8DmF9LBs0WP4wPW1VhK7mZ6MzkZRXpq3Q4jnQyhncBKwMgGmVJte
lVlXqIyUvFisy9lHnGFY8v4ymH0RzYXGYpiM7A6M51vbm6bFs+biLZOzf2Bp5uVbvPNeCe3dlo/n
Lh7SFZQ1ldD7bbD94TgIXRm0iaK3ppoo1wrms/Dmn6Er8fKlYqLZ9mxTgBzx+4azYS1Jbn15Z+5m
AhZofNjjGAf2J6cgJ6FaPPrbvm3f7k4BBVnMjBI6TxA8XxRREsA4Q0pwPnaPMzlxCs4eCny81ybX
eTx5evjXBnOfJoyT9lj5sIR0UamcUJr/tCreMM6XmVEU6U8t9NGFUK9BwO+6BwzCxN9CunfeT3U0
v9lb0fqjphUROeZdHJ5mEGo6kntjj9QvI18W9cmD3kCiHIHQFc3Kcexp8p29lqb6Yem5h9dF//n2
sgxf8QZGrlpJMtS/MixQGV6+OD8qWCWlffris0PRevkRs4p/UHYd3fLGzxM+2nGu5oJvhTCLMtzj
EKn6m3Ih4IfDJZnXtmts9xA/w+1xCEMRoc5DQ85MSWcVmwMRzn4J0P6+0lt7RgbAAz2sRC4niS56
PKWfBmMH3rrVVKdsQBRZZkDkjDBq9nExUAiTbW7HfrinY+iAzF3gWqr5sfurTukkatUQKrtlgaHO
slg7l/pTich6XAVVgXJChYw8kaNhyJ1SkY9BlBvTelVtkuhNN8TXeL4GAVjDQn/mbKAS7tI0P9Nl
knIQ5k54w39nRw8dz30VuYp0WZKwOKDVIVdo1TrPRJyCpz4APuSdbxtfHeUWLQz1F+APzzSRrzus
CWzTHcy57depVwjPOeaR7++H0+uTxe1lF3Xw2TTibez/6hUVCcifyyCDG6kmb2J4e1dDLILxm0Kb
ajGZJfu7sB7fmu0lN+RnGbF/w31WzYRB74pClTssQg7aUby35yD2FPQkNA9vNtd69YSjjeiBHnYb
jyJQjNOJ3+nUFUzTUMQ4YB99XbBMiHJzh9zhUAOvNlWbwcHBpFThasHen4pUrVjFr+j3Qzkmqwk2
9kT4YyUtAX+fpYwPpAl8INjfxngwyzjNazAZOj2aiJbjGlVX3omgiJ4ONzjcC06z/czwOAHEzVTP
K1o/TN1kHsCH8VGFnDHqsloiFM7JCLKN5Ojc3aVc1VTpN3P9zDB/e6PrG+BMK7MQlRUhsyBRL9VV
0aa07j/dsEnbtOwSpR84jlyBvaBasNual3qax3Po3IqHqzna+xu5QqXcw3iqTVx02ZHRffJ3whiB
Mpkfu95pLymJsiXK25pNys2o1xES1TNFfAPVlv4AyjzLF8FmMfM5k5jzsMN676KLPuwR5WSByhnh
YBm5+XuLts81of0nZ9puBzBHp7mfuwJJEyysGlcTsUgnjtRr7qDix2oWKjYMBRd3y3JNctOhEEuL
ZYaMsMBt6JViOoBPTD+oM5JjMwW3hHo+lyDwyB3FyDdmUALlY/qgZntiJsVef6f3iYsX1huSkG0c
7LmDYpkhB+9UFb9jzzxl7QZeroD7GV4b+rEBQTzP263WvQ6mxgpQGdT/TWCQiB1K2kbQLKiP86be
s52elJ23VWyCyWJgEdybp0LpAglkQ8fiX/BXQ5ciNAuvq4R9YYfvN6bG6oKP+FekL5c8zOGQeEA1
12cSMALVi+OXlMtsA7RAN6qtbdvABY2efo/SeFcyUPSaO01lXITw9q77sCDgcf1p8E5YDMscbSCu
u0SV3CfPZGRNA5QiToSqeWxT+mV+G86tIXYF6tyItXFHuezaBORJK6m6JvmglRmekuxk47eA4vy6
8atNauhZ+hQH6CcVcR0gejJVHQTxFwgmc/EnTL0EypIB8PYjHVn90PcXTiyZjvMcnCZ0dvWucNel
ZpTIGUt/8QI9anXeFEIrHbOWE1GlhurjfxkCE38iLHgdpMlZ5VWYzn/g45MMJDf8bUlbeZNjZzG8
zcY2bxnpwzg2tgraXvXi5e2C1fVttUMUg87lBbofPxC9mdhbExZA/XBC30sUhKik39BfoHpfoOND
i/DTKzxkdqC0HwZJm67yeTdwkNVCi0HpXm/SL+NEOb5DrC7Q0TmK3WyTXmTmAxhPhPsAgku46XnJ
Ba8LlLJY2SRgg5Z+sId3Jyj/u9Jxpq72bM87bT41LxbETT3Q4wqHoWmD53N6ySc3McPLK+sq85D7
qDFQub6AJmoI/bvv2WAW7izbReZMLj+kc6Tz7gTAit7eVPAowFFCL2jEvkVCuFOHz9DQEq1COwD4
nRmfPLvw3ByaW3lRUAPZ21GE/xVrWRJoupwOGodTreHMa70pPWkA5MCgoEe9Jk2+nCa8AfRIZqOR
bcezYEHbza3V6832GF5ziHGqUQY4B+lhEVKuzxWRGZTliZgF1PhR1hoXwDY3pqYpJbCynKX3etVo
miVc+kNc3IkRIcWhRXVH1z/CsTXdN8wDX5zeV4DBJJO4H0vNHiXwt21kovX6PrzSJum6x6Jc85GZ
T/Tz34/IU45dZ2lH2+k74WZKroyLC1swAh+uwhwcTZmhBRxvzLi0GUO4/ftvbB1k8IZPvSy5fdyi
MscIhX7MklpCg3LbUc5I220ySLkeLP4jJ9IB1XKyUunXN4+0f1LTv1AqyEl03nJVk6ZgvfgIOTJr
iNn0YnzFc786mfiBoKf4bVT1PbKnlK9Zn860QLw0GpdwluzxtX3WFWVO9ZQ9BgffoNRjYiicVoex
Lb/wH9ik7ZYQEZ+cY5WG6nnqyZnuzc+74j0TSRdVaZYOoW0Yiwq1Wfuqanzc6SiAkWxpbk0AXFyR
Oa14q5A5Y0JvPbW+2xT3n2fPw9p81s0CEoahUYIno9i33Bn+d7dy6CCZM4NDJnBpsvUMtaZ4hz9F
dHTzGCR3Xof0Us3kQKqZs9Xd2PsKP2lSj54g46wZSl9phrvHt2UsNwOER/Q0atW53eYvoN8X77NX
pTPKfd5FwLgmEBu++OGLwuawqU5ipG8qagE1BK4wyG88Ug84okvoYu1zfz4v19W8q6/Ok/p4BVul
kAu83gwz9Okz83qkeRHgAhwQPKPqED8uc+0AF1RS4gPYyrn8GGfXi4/ZFnUsScwT6LP7DsxedfEg
urrEi0BQ6M4d8dgCYjK5MvsqeEPRRPsYOCeUf4BOz0lnDiS57vSclyPsbZvc+soU3Y0U4iXbAirk
wI1zkU1ZAiRfPKv9mBSoYpPwgj9tpoX4r2IALK10njCQefNDOQY/E+q/dXiRhPE58TEN+figf3xo
On9veXiqFbTVtHQ5fUmKms+dOusD/d+JjriH9TCCkMAAsNREOEpKI48PJGeQZNn06j3A3L9S+MZq
TVEajUpHLee8KjeVivuyafLFYuVFpHjRUtA1V4qR/MkJ1uV8Vat1p9qlWggsjBRpLWpVKL6tovn2
yx0mHrNKyMAIFyBJuJi98woevSMwGE4HmplS3h2aDbtMZEy/MUkewKJBywh4A5zJX25LsQpuAuXW
AMQ0DdNY3qc6p3eq7VK0vyFof1KYXdEKOQfVRZNAx2YoEk48qnDbr4qfLzxQg5tHZnQG0SqIAVrv
UiTgylYFcqabilH6xhAF1qqZ/PdRBfldfJeudnfoCHqT/eIq5jEsnzOsg78WkdXio+CTYmhpfBuw
BzZJNo9KhwVABhX1/jI6o9Bg0D7s596ksZxa1x02TxFLaYp0yEzjo31IV+Uz4YkUNnmhDJYZIxKp
WNZLysqECWKNubMqHkycC1A621cPRWJJlHuzGnqUlKQgwQF0MeqXfgiVN2f/iIaRhj18ihPZe2HD
3Bcl+Pz7j1oOOKAa+MP5g3MvCV/tZwEXOOCZzqKNzlG1U7o6UXq+q/k15A9roaz9y0jxce/vp7a9
aPybV82DULCwR2cf7RnMi4zZdhFdBKxcSR0HwFJ/xcjgpdIJ9I4lI8jDTwUm7NOvWGDuAYQsbGFb
Ru5DbuW56AxLtJ+AE5fvgTdAjjteIyFpNrqTRP/ELGU83AvY5FYs28p2mGnrCHD9dg5N6UU57Puq
F65ZeoNOAcxuEjTpsHdPElC3btR+eKzVZXvYsCnHY1v9k4z/dwswdyfQhMn0IYhriMOF/OaCfO1L
RkwfpScqy9bd86pBwJxemfEIBElLX1Liq7CVYmi6xVGoJtxQshvRedJ23NwpdNEjURHwBx4i0bgv
pRbN4rl5muCFCjIZd0M6IyBT9IjSzVDpW/+Gkd79gP+MNSYaqfkySTBowOm0yjR3n9mg+o6GVCK+
TxamRy5xPaXYka+OOthHa/bklufh0NK/Oa3v0YoAD7kKizvclKZREW1t+njtU7zf4/11kvM+aJTB
aHmk3KrRFF3x7TGy3nQrGHHXL5DLIcXVvPfToa5o7VFDqiv6Vm64mLefUXmbPw+Acji4PJICLEQs
k6bDu30wjHtJ2l00veAgW8zW72Vjoa8tUEE3XEYP3bLiXVG8SVCbR5BUYMEFu9ko0sXap6G1sEAO
xciZIujn2+asP+Q+ot2gCuXMmz3x115IXF32zyz1bMIzJmPmHSExa+bUsiN36cg4906yXiB//3lU
nQ00ciYR0qVmB92hOfom9n0qoN5GqWrPNFLnDDnuepr5JfYchr6+SDuvI/M6iWSWVWPMSc4F0ZhC
pnW/8utcBZRWL/FYtQ59C0oeSI9gdM1e/9QUgJ1yjebOiyiNsBCjJVxBiyPfhX0Lr5wH8eun/bY4
Xy7RuKK1vmpGOpNq05IvnvAl1wWS7QK4kroG26cSPwtRH4aEmV7TFmL/1qWt0OxJxkM8AfACEXF5
+bScRqjon5ssBGyYj1tGp4TQUVVJRBQhF7niZkSyt16mDGal/IdSh/Gm3YTKDSvny1oNlmbTgnOl
arW6Kb0GYvDxJJuSAqpocdOkjC6duyB5LOO8OuBrFBdxUYVASZ4s1BM/zJgt8wvB0GyHbCWsbmk+
t1kIrV/KhWeGpvl5CFD+guOaWX8W9OUU5hCgtKtNm/cSOo2xQ3VQ4N2ymIqw5H2wxu0Anvmt+zMV
d6D7wGXQJm/dNI7jZt3SxgEzPBAa71Rph9CmIWC7WciE5JEgC76G6FWOklmxugIfzzjU93Ax6fst
msMJ/0sAjZ1NI/4d98voGxxnmHZ7hcudC10sdip2BrBYSjCbtsGDpk077odyB2b25o68FgZrNrPf
lTtgx5r1MwFynZqs2YaYvpOg2mWbveVYbCsl0nUgWNcKuqzI6kWGiIF0Cg68gu7Tzmzk6VxFj8/s
v5WLoOPndOqxyq52RHFBnq8kKf+0D56PQc77FhlJLg9RjqnAcekJC3nPCtwmJCfayLmdRlsOIsK1
PR8JCD3uYc6evJh/5gLOzkGy5d44D4IGU0NkwjFMl2/1REaB3xlyWZqAb0AK0M45HlEZ7doofG4v
ERfOL7gFaqskzQ3TMKpwPlreRVIgCimt3oLUAeGOwyRdjWLevaDq5lCepsB6MAwqozBakesHSmcT
nwgQhQ8+S89vhIGcbbbbe4eWBEfo6GR/rCU3hldBBJMx5LEFeHPkM2ZiV+vf/fELPO9LWcGqNXw/
f9qu09JqRyG+1EVQafBKR+0DnmQP2l3GJJV2D3nBnevrqWMnjZl/MWBNbijBnnc0r4jrKnyolZDa
Ngt9BF5bLCAzFWEOqhZTlYFbtp8ZVVxK0SQRYvo++QeQI7/hhPRwJCwCj/fjMBEyZRjqPaT5Bnkv
A796OtnYHsGgrB5qwST1Lw6ehAWE6QSgOdvlmNotNYYYUZMGsiEGutJXhxZ8s3WuoqD0dcqmJz9b
0YIiBT8GlTEU3vR/dBOkhW/abzegdYAbrf1DrPLjnQnNeYc3eLKC6EGdr9lLoSkDLw1MLdHI4OP3
ny246rT2N06h4TzdV0aeSjcxL+WGqNZESbVMfJuV/5UEL06Qep6yE6erIPD0uO72anfqlgAETP9H
ucxjY4f7GyrUOjqT/dXPJwnpuMWGN4TurVsAsSFxotb4rMXbNDJ/sOnW/uIEGo7Fi6LBRAZKRFQo
E7dvAGmCOKZN9aFds5OP1qv5ELA32si76cV/oDgiWvvNbdJkxtPwPaeU4Iyccv/H/2qX1jiNLyM+
NouheZOmaH/bD/e095unCiyCJiNtv7ZqglYUvvCjn87HkABOVKI4TTZKIJ9WxUI6uNL+TK9MrgIQ
eKTl4RF944nsa0ahzb/FJzzABrbf9uzVvVR9ouXH0+plpt3vleZcW5c39NbXkETj0Tz0HB9BBuUQ
AOZFDsvvPa9S4pjqBBIgFy+stkGkxmEAieBKRKjVKt/CjWHcHTeFtjaytbuWkGHdOxLAZlT0PFZH
BPKDBvz8ObJOeZaQDKBYcDMYxDH8BDcA+oKnlrQvglC0mzAfGEL//eX+LP8In3PwpD4Gi5Wd8IPA
qVYM+0vszvWJp1kb8cTGC3B4L4pRtV03G6VQG34RDnwmZbJE/EQ2UaDcpmSC9zxILOVzutvfOQAM
L3zwwRdDb+HYZtnOoN7rDzHcSczZgxYVymXTrO4yGJHGGGCRFd9bgflViP8KhwdYuDQrxHBckyQd
UE5zJiHJuyLAQm0nelEydEo68dsXx3O1Vaa6eGDVfpNbHkWRiuvtuBcWuiKk3sOPtJyGrADAIJV1
dJL1g1+KtPEFOIAj+sz7AlqYGjcmUvfGuop/CERpjBm/yfB8FJnjNfaEQ2OY0aSC3NHN6HzWjXVZ
nlP9OmtE6XReSKCpheiPn/0LhcuXtef+HWozOPdaIoEg05dADXiRwtTLl+tt4MmFdUyFjqdhgi1S
cQedQOSnMYKSCrPeQ+BOvJZhcv53FLp0M8z6pxDI1Cc2HabpaeVOaFAVzwSYbEtZhV+YHDnisQ+S
k5+pBVS9ch4Uwwok9IHuKHDQ41P9I8drihQ8pcm4m2ZvTfG+ATty0PYe12EUHB1vd6+nd5bkO6rD
B/4hdEpYFwOw8IevJHT0SgVbixnlR3W9/h6nUc2DvxBOGEmq4PakCpR0LMZ6xDdPv0mfrzpa6e5i
HezvKOv9kFZgQzPiXuJt/+ECuNF/wIo+kj+iroG9pH8AB9xPvdLmhF0HOXi6EOxyLXWtWfKM64ry
9zQrViVsW33IXp6PtA07g9Bj7BzXN3Jbz1ojOMiBsRAU5fqKZ/B5+GKyr76HAmFEvWkZkqCeaG5p
Gtkg9O5ofLCeUk5IMfcnSw02Lq2sonG8T4UQh9RCP5eUQs4jCPAcoZ7r9rnXYfZsymaa1s5rh+V+
+7mVCvLwmvFljiwY1JIPWPXVUuyi9Ce6WCFM04IymyrgzFxvhUu/KmPv9fcM1r1iWUW664L26uLi
urnga8/sWXNDsCQr9KjfOdFMpVJHvys7nH2OVm20OXG2UPAmlcbT+EvHoMs/DMX56levNKMKtIXq
J2AavGjUynrYzVSvdl0wOb1Pwhgmm1+dnLOt45z0frHIYzW/2hePsmnuOOl0S4GZOgnDSDntBxvx
TPCTQj1JpnnbgXvM1wmtWtcJl4bIl++AzIOpFemiG1DzQowqNHcyKTEHgAYNEG3c9aWfRG3HBe4L
5BS18odw98latQpnTr0B6jr0bJYRz8mNjnmd94DrReGQ0tiT8XYngqkxLixklQZg8Pbm3I5EFNpR
phKI2LzuD3ExoLa1GmQz7j76YE4OADcGKeq/xsiA5BMGSdLcR1SQCCeNzEjmaSyD4MnteT6H/vgE
2G8ykhKWmnRP9Mc2bA8zJZjsVDowJSKgpo8Fve67bR+fxO1Ch+mwDFLF2/kGbp4WLdyE3ChbOOsn
B/SB8SYnUG6xEXIyVOG3hKxe5FWm3ukKrV4l5L07dosDxAuX+p/uU4OVwphSpdXCkj3WDiiuUT0y
vGjPqADhQErqhUNvTxXFY5Zax5P1D6nBP8VsaeIhP+6ldTyEDnAiB74jWl0koaz6DdXZwvVvRQ7v
2ZelzmpvuFoPUmW0D4z+sl1X8YnZPx0j3gDA+FrWa0sKzgmQYrqwNs7yAlaJfocWfyEeW978lR/+
6dY8H2f6DvJpYSn9xX+QxNYaiBGx6scEVR4pSqFBSlMKpfU5uQLhcRz6RwDwfD+EtAqirBT/XHi1
xGMZqJkruTuZslHCtU422V53eprJDRktRJmt9OxlQn89xN1yLav4JOopOC42PBfaeyDBQZaqq0al
5zUwlqSi5H8LbyDBu0fmna8zcnS9NV0wDgiYXZSAywgr7YYjST49mgAcCQydnn++P68fL0XjS41o
tcluOSaqq8AUvPiqqR34o64bG+NmblLhAZynhFNEysjtP8e+lOVj50c4+eSUs63S/uclhOotzwx3
ZrZsL21sOWTnjiY62GvLZEsEQo7cL8KMA3uThJET0gr7mBCNlws6BpQD3nnM9JHx5pec2RwEU8R/
svpXAOfhuiTB9BBjqSVWG7ECLBPzc+fTmx27fflw2dr/61b7FOPAc4I+MxoM5MxStubSNGClZ6Xs
TuTwb9t1RYyggYl7gn55J/hsjyCpKelTUM+RFobZWZaQvXAlNvY27RXfzUSx6deSJFnRA+Alc4qR
6DimKDFDP8Oe+trHQep+U20S8ZxpyDpbf+UtcKgpR3QZ9B8Po4kWEhDGRjqp1jDwS9mFWrtXndxF
Qfw2SOnVMpgPr8UHEsQogo0VkpFZ5WmOIiPBsop0P2n/CEWZKPih/kR/ssTbuBWJwA/dGndZynoa
M4YA12IGI1gNKOafPc/+TPKFWq3XggXOW6u3CRRn4OdYKLs08cqaoZoSiojr9aPrtDZ9EVeakm2M
NxFSeD6okdJ2oUT5/q93pD+Ec3ewSBQ7VwFQY56MUHODANNSMS2c80yYsd3mS1DCSJH6HlwxlTKq
pUEA6yx/p60rbyq/ZuH1O+OylvfCuM1r/kzPFGzgYqa4ybS+nwkEHSOiBo/vZ9lvI0WlGprIj0aU
l2o0pKAtMMb99AHgoy2F7JIRUCvVRgEmRw3IK0uNRzI3EbR/FAt3Ufy9LQkB+O1EkhpYl6KgoGM+
FyaGPCsYNQ7iOdJmfE/0AnGVs78dZ9P7/v434Sw6NoZsKKsA/4WE9fmkn04kGC9MZVT/n5JgRyFC
RDxgeftgv7svWmcGM6qoukqujFUlxLgfxWe5WZ9yn49ED+xEdY8Dqbp2yrJr8blAhC/hrL8Xs1k8
YlXpMSGuXCOnxhUGwlTGSbMfm3C6VnpvsFjSx4tfhHrJqTcnHwE8Ah0ZthzysWypAKb77mgyOxgC
2PABSb17YXCxsBJ68MrN9DqxxIWnAgqranvS2A3GWalzMABnLROJPLdyaXSu69rtZFUlwrAwEA83
Bt5alq8lMLuPKulDDzk6piB1emwF5MweLmWuPwWcsS6n7px6OnVPWlNLYb9Tx7U/sT2dH6E/gBLA
aptpiKvu2Axm+UmnwnXkT5zNOXHEz5qAw1M/b2/AQFzmdnoBe4QNJ9gXfam81VUHvk1qjIAjIZNh
BeC9uQ6ZEDH37bPsatecOQ3xtE9EE6WWvkbCJJ0JasuP08N3I+F2Jvot9yn8PYBdwdMzUjpuYvzF
hnMmD4bS1UBoRd/lrHmVjJWrpgcKJRXtT3WIsumWIdUO6S9XjJ8tBTKEaBXG4bC20nu11fUe3X/S
wSpSNQCYwXNNEZTSEibOYz1RWX+wiJV/gwpMnDhzyas/+m5WN5f+41nY4e3UeIVx+25zXQl9qytl
IIIA9i+bM+Obv8fRdkfVDzIrA+NdtOJqpLL6+fU4gtkHyi55z/IT7gqSRVlCvRxS4pvG5dobEWLB
Y+70XaBmdxyY8Ee6/d6Hv19Wu1zcEOLQoCc79V9iE13d1mulyI5xg8p6JTEprrs58eh45WNuGN9J
qQPGpcLu2TEq+MreMXv+0JovhwtppJN+wT8skACueiJIep9y6b5B3XwNrQb+Vm9BXlWEOnbFgjzF
XrHVnpLO+KN9RLx3xBK/eCP6V7gbi+L4S0qfkJGTbqGqK59UB1tZZniHJh492tNnFiAkOyF4a4T5
ozBeZ0Sm0ej05V2eCF8c3DWKYAaUwiIek0JTZPnkPZfXvrniGSsS7hcsGxv9A28EC12sI39d/d0T
lVWzrHMYsB9A5Cj7vztfMfK/QGagu+LsqBsCPq0K0Eerxi2wAE6587FjiKwiyc+QVT9FoXA0oMfl
85OmEofCnvG4O8BY9zhxEn1zpNrMgxneUDykJVlZT07mquuyDSqlVDu8TBRWDIPXL4fsmFOcKlBq
Eu/Zy0yScslUYnzoqnfml7xafjAIGH+Zoj8E11FYDTpN+n74s4YFrprhVcap58okwR5LzEi/cDnx
lh/J7x/PBGzTEo7Xp2oLBltjDwHSAUnVmPa4YcMR3Y+KJnSxa0QZ6p6FrOc1kfkOIx1LiEfsk1b9
QjjEYK3Vr/VaQaW1YNC3SZBBVn+jDUrrAlRXtMLoxECMlv6w3oGUkX71J/RudWH9rVrTAp+zP8On
eoFW5m8ETYS0McWsVOZJ1LXhA+6Rl8cARlavR7q9nUv7Vm/AlP8WJ6FQmPTt/hMrt17/k8VCIz1l
DRMUisiqvoL7cisMrTR+Un4vQf/K4k6MtJGa6Tx7yf0At1qgiVsM5ntUpk0Md9aatpxC7ALabYBr
kOIDPIXJ6/RKE+1pHRMxOMJ2k9c7RlxNJMH+/qeD1BuvWHxSxhLd0IjZVOtMORDtMLf7a8dcJYIz
7t/FqDT0kWIUf+JX9iRVrPylt6hOuVgpZU+ak+4cKeZR8NmLTwTh6foKicA17OqjcK9r+VVTEiOn
4aNwPSpquIIK4SNHMQEGypjYPXzElTYPd0LqFU3DkFXRmMS3LxGhEWiGC/mSkfa68FoDYTyNhiBf
PFBau3fR3YCai9bFMVM12HSt6UavSbxGDPCQ20aGsqrvgJtK5PkZzzgLS6AcprWCn7wOnQIAlKv9
5KUEk91OTIb7Gc83yfXb00JJSc4UeAysXJNHu17mM0VO8DI8BK7mJPgzjD0RWtpz6OS6BDHSvm/r
fxeMHxzgA9Ryu9fOF5ROQGywkQgAsc+Y2mQbduSGXnNgzjB9iajKe945O5Tm+VVtV/8U3nYjFhDi
+R4sRxILp6q5Cp2EJLFh2v+VTzbo5g5OnogXkxawaTADyu6rcwPqR/fWtOlZiUUZ+x0ME+2+MyZ8
iGvTTHyxtxS4NHvhMk0FDDdoGtFqJ5m48tWHd7RWP35rjE44WZKN4+C50RiyAAJGOcWkXE3A9PrJ
DBYHGb6E8EhDXTpP7bAoqoNRT3qWBuABi4WfAeZ4AhkQangkhUa9EEDOt0HMdbQbxYQdc7KGLMBd
zL8WqYum5XCgCkNZehuBNuMxZ8eNMLVmVS+/jiqg+Ir7u6uwT8c30A+4RXeMUSx+bAZtlyMZn9BD
8qXNWsGIpAJuWhLhLRPAEOr8RGj+Q87e+cE31QNU/+L47QGCCMoeHaL7RtKSHDcoE51h5lZHSaBj
15SSydQEfu54zOIvlPbKl0qbYEWc/ro9fMZRIJpMHBVqX3+hJtE3i9z8i6XY8PUSja+D0ApdXmjF
eybqhHVyK0gsTO1kh+2pWfkOwPiXRNc5xUpXRBHk0g5GV8FNz9djZkid0xId0tj0qkw44jn22gdO
YOoemMY4HcAS/+lGiRLKijsseb7Xa7Eq0/oz+PbOaI1OJEBPDTfH+IcaospaUtpY+6jeGWeN+t6F
JGmOeGsjfVLuYOuheZyKh27CPBY5YOq57nqUkAbGc94gaPgRzJHA8HqQ0oQIXjUW6bOSI15d99hy
STvRgLZClaHDSe6iSUHotMEoDSSXHuh7hOWHUSpY2NaPu9ljKb7r6tgianPZ8aBCqBP+AdGhq2ha
hmZnLyq5Ic0CaIUSstFxoXEyytXjkp1cpnHrl6m8tQ2bjttBmp45SGaKwDnQjuPcHu0qScdYMOen
FzsfYpn1pWFmUi1aK6AMVyB5eqLZrDbFhbjvtF9A1/3KjGCLlHB0TfUA3xZ1I02s8TWnKeMk1dCH
Q75iT4Du+yBGPiW9wgiiY6ekL7Twuum5Br7mfAYtE3J9vDks8bRlWBsxhaAiN1zLLTVFtV90Hm5+
2fsZ7UN0A69C/uwo7PbJTOM3OKSd6d2RY3tgfuX2cY0CIefx1QCQ1+WpJlKq6QERde0J5OJm29TD
l+ZySor2i3RMOoPJjx2RdCVoG/Jay6cut0rbpdku3N+dzHwflKA0/DJyo/ydqKkySEIzWqfwZzHB
AZRw7gCkSX9Y3vhZnS4B+Z5FtBxylxgQM7zrRYpTKO4V5rN2kGpFiGiiGNDoy/shGhi7pNrXOL5u
Q8ZT60ybyDWpnKtYLWiPGdEf5p2K0Vy9CgYx/gxQmbntrw8F4CzEmGloL1buQsNNdCHlTIDh/EZH
zBbPBPcFjx9NhJ9bNaVSfVifaJJSD5g0gKNK/DxEubxEBZui8dgEU4W+bt6rpRq6VPx/ZkZpgbJ7
U5EIc8VwOxS1QVwrtTSd1+Q0hxkiWcvzFV88XFU38nR/JP2gmlAf550fdTsu1E7hABtwhi1qFqui
iNByl5KB1K4VOnsMu+zyw2K9b7YMibCof7bDjB7A/NZRw5lkcZryF47p8qUp28M8DanNewk1XT65
rB+JU4dt4zlBgk1DucAVbyaQFKpyBDWOVOEwB6oChVxWnIaHKlA8cL8AccW1odST6UhUkRC4tx6S
PN8MpRICUXxkirFRcQX9twdGzrQ4y1c2zRY/vHkJwGuZFB3wVXFWKf7litk5g0KXggtQzmtaas4D
Qqcy7fvQ/JSRmT5aKfpIjCvehq3NBDzJT+tBZa4/r8GisufC71fGLqLV7lNX/L4hifqvN+gyIFUD
I/uHwtusjztEOpmhSybcOQZWLjQ462C8QQ+zaTZVMC9x9TXyAmfS3bpnI4ptfdA7KA12pcY7F4w1
LoyAxKsosGgKRl9+4QE8zpowP7TW8+a5snhU1ttsnE5qcOqPBUTVifDoqS4FbwTeYY95b+fZ05/A
UD37EhCDNnMiXeFIKx/yYDmZd6VcoosBNgmCmpsXFW8KWQ7j/gq+Sdxl7m9aMm4qzRdYOP8eHqi4
mt3fOCnS86gmeT14oHdEEMYQ1eEP1VoR6J0N/o4E2PsMUJWPiE1+yktTkM3u0e5FMUdrvvwA49mV
YycGJbA89oVrElx00kRgVxEuaxT7U6hWStWVdVnToWwnutKwi1B+AGB7MEMPOzHI/z2aAhrkzp/r
zkVvSKaM0sqrUhd4mb1em6edBAN61vdOFiaVoyS8oYOUK9/buId9xRO5NXvVG39Zfrs2yZZjiYPe
cw2aY3chyVzO1vUcNh9AY1a73AXmdwbO2AYEImbJwoD1mbEhQgCBJuyW9HSyZar8MSHDJto+UQoD
DZPoSumoKbh/9fpH9j2PywVFShEpBjGr3jhgINeX/msHLBYLEhR8JjT8qkyN3hSpMndi0k33VJtP
J2JPtzWlVSiDhGjydwRTXye8T39y5O3LYsJiTPmB07dFQo7pfIo6GzGLblPCwVTeK6l81g7Ppspj
BBRQMTllXDCbZ70FyE3pdEt6PiCJMdPiC/H2Eirxdkvh/rtLxYHd02i4akBPnp/GdRGQkLZtVlGH
DQNU5luJ87OMlguv+O6IxeJdEIBZD70MaZyCdpD6EpW1u1cCFB38uSoKjFIcLF8Z6AW0hGDKiaek
gPL+a4U8Q4GM7t7ThsdARFe6wzjDXbPPymMYZI7msd30yK9EJf829XPsgvLnswMlwlecZ3RSP/iu
dtS+eCTJk6BqWN2B7hFtvyemCmreL8tIRh4+oKPkqUe0Ra7vQnF3RG5hlK0uVamff8MRVKm+fFQK
kVxff/Z8KSNo5QuElAlH/ZRo9GgPVFVQ+yoxrAds8z09fgYATJIa91I0Gd7Z4sP5fzySakNloqF+
PLaS4/XAkNRx3ngt0tPfpZBJVP6sdCRQ4MqsMGPbEXlekUPnlSmt2OTbtSx8ynXAgjtMcXA9zVic
Bd/XvWz1ypjIOZBizY/1+x1jNjpFqmo4WQMGmn0+uWZjymvP7MHxHZzxNLF/stC3WC2EsJXZ/ACP
KsyDqy+TIYyQFM0bKnVxqjoZGusMvT9WLqRVgQh0dvDop5XOJJSAahp0TZzVXFVN9OYP/DqtRQKy
96hM2/dJrwCfQQfgqSOWUYb0L1AEXeN0TRJNGnwt99SVYvr5oZWtyn9iFS4wG0YmTtTdzQ/TAuy+
HkuPgWt1z0meAfjOePoOv+dL7/fRl01dDGAcOjWBwAsBSY0fBjazBTJFothXaLwV94BbXbQgOAPp
y1fzndtEKApoD/PZ2fmbSQrMY75q2aq4IsSAuqTXbb5RrO9i5wcTIbSih1a97Te6JygReQ6o2P5b
1AAPld0ITKQymmGNYuGqMBPEo63HTXpjk36jSx/KbLIm81YkBQqrmVEJ2UjGJecp9y+BWI3XrC8u
qbaFYLKTzotD4ke51WWCd1BRdWTTMSVTzuhlfVm+vk8vKwq8WOJbobrjnux70lLNyJypwR8pRsP9
jouec7VDAV+s6GrzM0YhLojzUbp1DghNnz0nEdx0D39S8KdrFWD6m8WSOd9/9zlegt9ZYM4EUhf3
Rq1blHDddqOFPqDTjjtFzV2Bjq+8AK2k+RSOVxpg93BsGI7ltWMlwzv2vCI/259/xyDxfTiD6yTa
rFgfn9lNNrvPstbzW3iXIexEbYC6ZlZXuDAhPWcelGkiGUf+c8aHmzQLHCeowR5el0capY/WKkJS
Z/DR9npsejXPfNfC2mkf+0D/eZ8lqwf89WLfADcFbxccnaA+SnMwmvHeqR00Mo/YLnUmdCPTK4Rl
JL1cCJh+v54GHTG1sCwQ5QFO7MKsXMLUE0jTK9pbjoCisXoLxLcSMC4KzgqCJcndS+HZIXdSO9SP
mYZ3IQpoiWhqF0jGTEJZcs8SaP6s6XHVMP/GSj1pJR1H5hxL+upIS9Pvmiclbhkbnx+RilidWX9s
W2WBwODMivafmHEHmp2ot1a7ywvlR6H8r9MoiHXvD733/b67wTYT2Zq6kevgquT+MuN18UJRkwh3
o7tSlfJ9qFdZkDoyURmV9lPxzmQBvzV7TgHEVP020gWkECNXnC4Ysr5BGRuvN6468yHDC0UJo/O+
PHRwnrQSebQgn4HhDlP/M+O0yVS5dgJGWGV4p019ahnovpsBVDTH//mqLk8b719zvkR3S4KjnLQ7
hvvCoVwECdTF7XbwHedokaKRVVyOxYu476eCSFLIZR5mHI/JLINHit9ROym6Tb88k+buIivzGHQR
IU05A4dxYMBveLxUGL50X6LKkZItcMlL28kqskN0hu9to/80SB+W/UW4Mdp6jSdwaotvnqllnTZ2
FjoXCJwUpSITVcsM+ol25yEfgAE0qu32UPgpGX7eZxtUPH3y+oaiJVLLbJKUOD0bN5TAiSInw2Y4
sZpDzz8hGxu8Q2DH0blNKI2hOkW4tZDrU8+2/VJq1MGQsYq+Hgj4lDxBfiU7At+J0MxZ31jjZzG0
8ZXYAJnP0cCNFYiBA3OHJ15lqB5dIag1JfFJUsAIop4MyUpfFCiBhNOe/d7xTqXS7+Si/ESdWqfy
mZQQcwuAQO1IxnzVyBA7vTytfXFbd+ZLoZZUNutMN/xNfsD6O9O1EBCfAgcvnLOVK02rypUPrkXk
821wxRKcag4cyV4cT5HLblrZPaiZi9nlBB7iPJNnnYH8dsKMqHHzMA4OxIEKw9uQ59BJhrCBWuSB
tMkaY4CLMTBJmEuAaGMtw7Vedc+aSodJIkTtjPS8qYUacJa3Oz8ki3t1EuokyWC30N3HJFEG6zbY
+UTk2A9MM53/pgPzOPAfNVNUATT9qGS5ziULqBcgbU/0PK5UtL/Nvld5vnIJYVqn+/C6341/813l
7OFMeIM2hUHpWGsg9CPOgekaQgQuFmbEO3OcjwK5PKPorBAPQRy/dZTVnPwMFpdwGZSAvZaP6AQF
9bQyxWrWENye1MZmA/BwS+fr5sP4z/WpBExL4dAP+G+P3Xn5c/Fc0PD8DB1zpYLcgKL2FQBrovAr
b/99RrqH4DugYNA2u5FSSMyWXgfNzhMblrudWJwaxWWCl85bZPtiZWD5TevVtVF5N7vGxYKrKDay
ZoCyDdEtwauPLtsckFDt/GflXc5xsiPD6CBXuhrbmcUpjJX7lwcpIZH3WJ4MsWoB93BszgCDNTGZ
dHzsNtiXkyApN2H+LWoBaIvJB6QNzf6JKCM5UFN3ZI+dqpYKOzd0drCLi5jTGZvIP+zlFrSowTS8
XoGWrQ/FlcJBIBbniqHpvE/fvzmzosoHpwtVLfiTKNxJcoCTZtp/Y8+JkspUoWNOq/XsOGfHQnv4
8JFs/01qDXzSlP7wLCV8oVjnFo+5kAQPwX3KAqGkQFVWaDi61naq/QwPy4RCLheLS+L1WsLg4zHz
Fd0PUxzbt5JLyMmRyWdxmzWRW4cNc9J+cOuaLMwsv6cjGQmSugCxDROCnDEpVpR2Kt8tA/saJIPl
xaPxZnA3PcvK4nLpjnDfacGI6/Rtn935fxSa/vspKJwcR8RaoMBuYFnlQCQ7Bs91rrHJw5+RSnTX
+NBlS287/rBwq6EZBygHgnQVp/om2igwhqEHbhDOYvqk1Zpst++Ku5IEoKLnoMOJUlQi94Fw0xh0
7/6p5i4jWVWwWwjJKffTy7H2JFGTrOrwBiEpw2d4j2/zwkGuJPfR5JDvXgUsVP/iWf5LYmFNTze3
Fr6wdU5wb1iBGaOf2/G2PJz/XNdAId4pEOb/iVzgKyTgB5VeVioShW0Tzpie6ExT+uNSWp8ra3+e
konLtLvCmygfhj8QFo1qkPpfJLsiNRVEeZ9AUgmYbTOToyJIAwJ9E+rLffseXuymgWtS5fgSwe+g
y8QGMoSCr+pm9BkZdbEWNOMC5jDeAK4c4vYexPRafbbiEInyt9UEAaj98UBFYgcovmJLCbtQpDXW
KN7lORedLxabvMokJ5i7Vny1uJHCw2KPKtxrF/J8VixQQbv0y5zmGEvIBjnCsEGYeQOuXqDFF22u
ijNMT56jkzJOWstUUkEebe2odRae8Wt+LilOqbhTzlf9xR3J6fke4qNFAQmJgLQQetnbwF1ova77
5UeIiAHUtJb6Xj7BGtFqi8WoLfuv/1zJu0iaBeL3IQW4TzJ0LhFciOzNlrFSeFbNySoz7hM5wRv1
ifSzMGpDPd6LSsMtvl5wGo+k4xFQkRofgkYnt4eNaogK3cXxbItEYNxqzHXB9ZnsQemnMiKGq2H0
ddOIFSRjcMUf8VqjzNyJveRRr5Fx2BUNWvM6eJqswvk/3OCSRbxb8N2ECp5KvGt8nXIw4xtSynex
1/VumWJ0/XkqHNXFVDEfpFVUU5WPT3a43YM7LJYDUvJX7s0Wne28lrzq8ScQOPwAwSbrQlS2ngsF
aXx2bC1Cra/ML3OqrRnnGHJxeifeuT5P7T+hjp5yh27snDsCbRkLHnM9Ctd4oX36B2KZAutz7+IQ
DVmobSumXfNGy9rhZDbqQZmjLeoR0NCXHTsecrzKFDkP1ZLXOlvxGyQrn1yuDKwSQYEzBkZh332u
s6uwC56UXBEsLXKJcalr0WQNYsdiYUH7OSb349u8dRqJd6JdoL/GgKbrYJqqlUDyiwmuHl2ede+p
XD+m8KuW4dBdC3EqA3Akj2KlvLycfsckg7xnVBfblxcDgtsHXZobVflWs6rG3yvBtSqV6kX9Kmue
wQuRS1megfMv6KERFF/hx9lCY88CVQ7sgiDYCFOB/4+5n3zwjJP9kZsQTcObl94R0OR/eBrvSodB
MbY+j7Rq72augFj5XOCpKl/8M3lwdN8iTw3bdjMD4WJEy4Fy3uTt7acgYWI/oymRXDAN6I6lBp0k
KHRviWem3bcK0Us/caJSLq0Pj4Es5+2BzzmCnPvnLvl2h+Jx8eEblH/WT3Q0ut7asTGEuTb7wzSi
5NxydMPaaXOC030X2WtP/Rh0MHWsOMJra/xokRTEWKM14HVjwjP2qqPgr4GR9nQwV9GP5xoxq4g3
OgorVlVU/mrUgYGNBKPoAOysghulZHYWSzLPZGrbyUOtSu2bOSaop8D77iH2NorzkxbCwQTZH54w
v06qznK/O3fP87cBcdI9C1IvReIm20ffR1AEHrZMO1NazJrOOIh5DdlUkKjC8hBaX2g05rBlJTK2
ETR2X6ikg3bdzTH6L5Uh6sbl36VkKfm4tbUKm9pDYqoCY2HrXIvvAWYQbm1gsSkztiiGOfL4gIhH
iwz6h+Kik6gS1pnxxQn1A4WQ5x9YZsDcDOxV42SRS3XRoUtnBVSuMnKOuMKouhVQ/b2TBLxhX2jF
GstdAcRGQ3GfUVsZKzRxzb5Xm12Ow9TfTET6zrn4kADND2jT/v11vwrimoA+YJn9138LQ+h2aoXf
PSk3gpxqiVgmGz2pXpb9OZB6VhjK5ova8fylsz/1twFpfFHCW3UOamLWajCOT7sT/JJZtfbGh5Bn
1TRRp7YReeyXdTOScw5M6lRN0GA1/Qu3qRVEJozvoiSGa/+NEhc7AdUZyATNqzlj0Y4GlZi5bOEe
J0pqpVRMqkgrZuPHpBtDXo2Sb8IZd7TCGKhFdngRXibb+hJYghwq3wyXk1sgqrLQr8ARvWl6JpEn
mGkDeWeXHyTjbGbv24pZBbFcFNWlg23iSTryoenvHHusDRXLL4v8qjjPHsbs23PXHMGkwO6j/FU7
6o7MuV2+yC2ARjcFMhgrfxDsP3/fdAGbGG7XQ2dCHLGOUgdpmo4or+V5rsIvMAg0lcFhQV5i2YzN
VbEvDE9ZmqgmDyWRrgPEa9KuLRzIiU0UJ0di8ir0jTcwddXqPl/UrW/C4m14pjTy+SgYpQF1LRex
h61vNa/bESNGjUB3fPW6K8/n5BDPvSSQJnABxrwmpX17aOigyyQrnMZMeS8AGBRBgxNsggn9k8SF
nFkzEUO1BWgT2S/SieE1z37++VjsDtTbX0hQctukwQUG65UP2rffFp2yNHxMwon6xq6r7cHzhiaZ
VCqfhes7GJB+sL30LxliTjGqPCSDPq2Vhh4PPwirVgz6MBjgo6UWl2QJMpHqtCmi7JI061rGgG+M
RlMSXYo09Updo2AXRdAa5v2ID8y67jMVY2Fz/gsqltIFmBoh4XFVXyZ3iPCPyeS7gPK5V1XdNiPT
s+nWooe4CHzjz6MtQoHc6LqCGZbJzOwSflyHAL6UKLj41Maf2sHsaLDgMMu7mbo6Zy+zTHtL90d/
DLIZdl7JMDrmXyzQF+9mVwdcgedXy67Hq+HmqDy7rG+zg1PZBTn80KuBtGzcWGlp5Bs+h56k81xN
zL3LSGQcI4A46k7vtGVtBZynBaEMMdRcYYdjp+Swk2+uW+WycGASUFJbEelGwfRZg5kDG06ktRkU
jj2y2Y/yU1+/u7e1Z5qWmSAIa4NiZS2vcO5MuZM2iXmICSf2ojPVTVJB+TLRVL88xiCemY/yRgOt
OPHOXfJ+gJSjq8bGXRoEo8AHFRuYLiQFaNX36CcZSqUx92jf7ThTfoSaReJ7U+cJ92pDAWTAfgTD
YtsF4cLJfICzn4vDopUo+aqkcJHAqis0Q8t9zvakuUgwlA8fi2QubY3RJYYQy1fkx87VpoCwXZap
Tb142213W7PJ8OOwAhjnGDNnuGfO8eWJo7+P4hWwpcBMqTW48pBKVO5nAoYNl28kCKJVfm0eLgUk
qZ3P8tPAdh3Bqpnp/gorWPv0ywiQ9i2tlbiOdUftrRYlZ+LzL787UMJathJ03/oiW66YXVVeRYy4
KILmymd1YLP6V5ZmIA5erjlngwIiM38bwDiwpItDu1lMIQvmljQAoTV+5+rCAjZ/ihgolrKRys19
McjRGSpuMz3SuSj/nTqYbNtgXw5cQ9cX8VRhX0/e7LITUS3XS5K8L++LAOLH/rL4ALqr/PFWedh5
dj9Igvy5g3T8pLmSLMcfT6/m7VB906iqfSIeKT1KiFXuMhqqjQ/JbRSJzHYs32T3w2mKLdLjPrae
SiravSc4tW2pXN6unosScTreciGzoTBtV19t/6WTixqVEwBTzifEXN7cC2zDdDQPyqvwxg274+FH
HGGjNcxs70B5mz/Gi0UC8MwYJPiTOvW68Ofrq191wxGo/9EZhwAoSuEO+cK50ZrFEpsHjzQOVgWD
3VScKYW6HfsQdvORggqUtxK0qdKBN9mdnxOwm31x5Dn42naVsrOUjpO7FoaSoKMACwM3Z3AzMRZl
5uEQND74ckmY3ylwASxmIAN7FSI90fRmazin0o5JHdji1i/2Tuc6VOJ1bkqTHJz2k/MG/MgWuzom
2EAspsbDQnLjDKvQZLpqseR/JeTAqukamJcxKbsoT4JKfJ5+S/vl6ekIWa4euHaF0oRMUMmvb/ay
2Fxi9Qz/ZhyVuLjInPBuIEcCEBQPgzQjXdq8lRwFPcxoA9FgDJvdCKtsJwXz9eQydy15oH30w9wQ
9iUdqx3ZfB563tRzVRTFq8hFGE1MbI8ucslI5O3bJ1IOC41paE9A52kmDlQCvfHizMG99qZVolmP
OYQfpOWt7yknML3OP9K29NM1I/cNAgQcf3BHFt4QR9EK7iaV2nuBekpFxc+EOEhsBJV8TUFB1YYC
t9x+h2+NKEnnvl4XYnX/jW87YF4bZFdzwtKa4fWHWGnhAKvA2LWo89gergnKvpg5+exgJbDfaDwU
kiGRsZjex6kv/0+fFSZRqyxs0+jQ+AEW8ASpK2rmJhv8FCOuguZ+pmZJvLs2PS5xlf0p2VyIk2lY
lKTUdKnpd9cuGkBglAluyEConJaqJPBasOLJVFhMz4l2A+AA3HKtkSypsdteJhr4l9/c0blwdT6I
owVEjqn/KE3W2PbbvKXBGcOC7tMTj75Sq85OzcBo4TX3PcYpTubnpN416shJKc3sKzR8BtdI0gIf
num8lmT6FtGVSccaeGzZHVaX5fgvSMSelAQnLyskLJpMwqg5yqEFfMwNsVbTzEe3hVcM+tYnUIaM
YH4jDZt1lPQ788anWoyOoSSmLuErw7ifCdsQmwFup1hrIMAsjyaeov6zocV6nekAElJWrUWx97Nm
oEBS9H97zv2EvAPphtrI/n/wUs5yp0xAcbCOqDAtLkBz/ThJrKGyPPXdvCGPwdar+3AYc8glp0S8
io0QdlA8xef4zbU2Vk3CBGRDcT0Fie7FWOnVlGDINpojAEeyoiXIqFMz029J3Ic4InERNOgjYQRC
QYmOFJcOFymmUp+6jjORSCyuG7wItPzofTZkbsjg5lTo1zTL7WeerZD1Oogagn6ex/iAV9o9nFf9
LiNX8o7bJvj4CPTQFKnvMu9Va8+UnA/4S1cyVZZ4+BaIZTkSzUlqnA4EDRHNAW3BZPUjEDDXfzMd
tSJs7U0Q2AkF0sXhNzl2lqeeV+oKSdsGYm1KeQdnJ2xwEwCxlZ0GXpsaiaUsjxDGYlysFKj9sVfs
C5nNgR6obUMEBim1KUMWyG4XCJaxD4e13krqN76PVp1esCl57wYn3n3ykC9D4KAZrG7f2DgMqcWE
x9ZVbTaOgjEJhAl34cNdGCc10QqJ0tZUUu/a6IOguXksGNbSlTM+xT7V4jQ3BiYEjRIPCutKv+ea
MOUdIucNqU+P3qPpVWHDywGnkjQD0ApcLI94Bt02XIITRVQargTqykOk4TVuJJgFota5gWHfVD7i
sqJqKWuCnwPDX9PQhHtNpIZU2cZp3hG0HmLGQlXGQZPrIod+stz0PfOkkFdcaArdwHdTpuLyNTLW
BmivnKTbt9mBquaZvWCcQaL/PSD+Yp3XsjbfLLokBks1CMbtPWurnLw9KveQgT5UFc0JXIqzSb4O
+XmsJVqgXPKuX4XPcJjypZnMujI8IAJLbzExKM/ZMVXBaq33GtQ3LzU4kjZ+TveucmkG3UsD6Z3M
iDNA0zMUcfstkWHAV5rGsNRFxX0RF49ZZaxInWHFQJnbcOXUY1Zd/E1pPZuz/Mqz2GAJku5krpvN
rjVaM2uzMCls8IPTQfk2pW/Qsnbj1cuOceJDYTmvN6PesREdiD+Jcy0kIARUmooP8LPMmhBRU0LD
3ch03GE4PPPYh8o5HxniQ+EQ13XeskITWVPza+P2rhEIuhnQZoPeUqDsu7RZpbcbsm5h98Tmusle
VlxPBlZ4ropYcXirdNNqn5fkZUtywE3XBFFjssfPopN5HjnXn05zLzCcgB5SS7G/hVV6MP7xLqZ2
RQRHkofK91sOj/mqfqBp6QyB5tjCzXM2+DG0LuIs4xTGX4M+rA66b0P20yZKUyjSPKW6H1rSDDuN
Fhmjz4yjjFU0Rp3NiyX9ywxEMx37V34dwq5JHTB0t6pFKEdFoYNSA6+3cKb9jjLsAHZtuNqHk1Ng
2KrEXsYBQdgYA2HWLmX31hvZH/1NTpNButTAllURTYQxU4E1kBl37aYRlt0DLHe2+UHwYgg1mDCk
t+Y7KvkppMEY6HS2LKszPM3zZsgKissSUTaUboLr4gupOU7RGUQOpkxnCxFKMYLM6U0FYqnMJaTL
civjva0oCWxauYktyak6LVsgh2qdSF4xN2PbMMgFeaoa/TUgdaaovRhgOyjsiuhKNGSW4eNFvk34
J+pmo5uKzAb6vhH32TydaZHLSytIgbRf1wV1yxGpTEFvnCcMCyqnOkP0Wb1xxK82FV/9FUNvH0FN
fB9nTomOWaD/4FBgWkuJgaX9DXsomiVIA0afuOd51hnYKHnGWeRMTK5JPlQvMNrvHAqD/A2C0CeE
6mCFtyuvOIX8LO71xkcSry3yEaXR5Nb1F1sr1/gRfAJL4xk8n2oU+YTdk164p71ljbdgjJzIAjZK
8vuIWfO+84/qcxE++aB8sJyR4SQ9peRHHfz02tFx0BoAgK4oMYCeDvAYDd5DkpKEE9XaIASNqiVv
xP8qjoYLHNHhqZcVwfUwaWhd2g1C1J/whT5h0GbBvTM86M5w5sR+n0kfY7Bu4sBtEuC2uD/IwE3Y
xhKYyy8DoTPbRRf5ZoDyarhYQ2o/fcypBDkHMkk6wJO7tq3vbnjXTwsbXLFSxSRXD0wFjl1pRNW9
G1kEX5o6upcDmJ2nr4K5rGr1Iz+MUMJV8t2aj1WGOesFBQin0vM83NFRvsl/1mftUJ5YBYRG48Vh
R+UcjwgvlVaItbL+6E+NgSJiCa0lMJBcga/KT3FV68qQt1lD85awThkXmL0xjfvMx8tH7AIObQUx
m3hZHMmP/ezA70Bl5Aw4FHISiXnhpSL0gRTZZqrXMZeM0rOs7vEBuadW/3x/JVp8vWzmIXKgXgrN
EM3GSAPv6v2YH9gxEStNWJCWCfOQDm19QvVl3U6HrijTLAXnht/bn5GuwLMPcjJrPMPcjUQ8hMvk
u2n+hPVqUvO4KkX1vcqGLBgHF/2clrHm+gmbkuLISRViRP/c+EXOf6SmXClio3SGgilztsuUoXVR
85mP+zNnIMHtzAJyLZ1aFOklFXdYMMV2TXkMQ2qGeHn9IhbP1oAJxQCbKUz+IIgnkS9xqJ+vDoIT
Bi5iwePAaiHtJJS6tRcjSxlHIdc4a1E1ZXomXWaK8qx7kM6qCcytSushqGHzJHkFJpSWUsWUVAet
d+cO4v4wvLA5YWLfQKoQpzQQJws0rBk0B+9DzpH2PwoxS0AogLR2f87ob+TkM6FvnFsV/bFKXEE4
qBgUxlDnXqBCZwyfeZYl6Mr7whq9Fz800WvW8rWVGjb2KcsEUfZhFEwnpM6t5Xa3EM0bpc+x4N0j
bk2HO8nWBYZSIzGCn4xvKJIJB3C6c6evNmdhHRMYZXdhAV73+FIkb5YJ2tkSzYf4WjDNA/cTEzo8
BGIlkJ0dK5Q7DPtXvQsDvgc5CDCDal7PaaBTyAdex9M+SyMHKrn5kWKOslMKDMIly4kinh2s0yqY
OrR2x+WFdsSR53Zi5VQZ5/zGiRThjYOdRLXOKMHjQ5zhTRX4BbXuqhDSAgFx+6NaIhexwbo6+HPw
MNV9VoIyAztzoYRqXNhdCiWdqjjkelRK36Vu/UqXd5jyLIEPZwyjsQIJ5qUDZq8QzI9YwLhABb1L
LZoHbvs6P6NJm82jQZ169fEUsc/kRmEhRgWhBM5JHyjAToC0t+ufeVgXZVB/qva28YZ7Yyoh3hSR
FvpNoNEKjd+8TYD7yKfouOmD0uoL9Byl8+NkB0c5reI3zs0pQQwseW7bYxXZyV7U36rpuBwKRAw+
Nx3+3Q2v4Eie4zMqe7eL4FtdMj8wZ1jp2WgptMMdR+BzcNEDGc3hGdEWNWeOiLbEGbulSdXbmxKz
Otd0/EPq4Ldfl2LNl+WWZUNeo7g9bPvTYNSVgLZnvy8TxPop71w5ONq0c5qkQ+/T2HzILr4paS48
WwrfUjAYwFowZ0akftRu2N8nrTW7+94ASvJEDFbwdqqb9Qt3MIn9Y35p1NVbjl6ql1pS318HJcat
84pI4Z6YakpOdB2KgyFX5BWHGXCnB/Uwz0Q11nvqv6iRFS835HRZwmZEJGEMOSp8fUQG5aOVMFwW
KtQjsuXcN+kA1RXAahuSC/DJlvGGilQiHLOk1Zj750bDXiIoKQvM35X8vjKQnNpQNqnVg/MPh4Uh
lcQxFY4iC0oZo2kezGy5Atu9lRPTNcPkIoZc2KDojBFKcnqaSleL2MJeawGOSZVkkWDMIZU29UGv
ko9FfvRPvJqbYWZtvXO6wSqMwnkJYH7561o+0o0ah7JBIaK3hyuc9GEvlQpE09ykBvXko6OzYhKj
jItgjXZpEsUIHnFmmTN5BVfudpmorSSgcNV/BAFjMWlVHjW4yw75fcaqeOED5lkMAfhGMYN1HGSi
uEiqY+a7GcSZ+qn/WFKigmRpiNniU+nnnt1aTV9l4wHGUox/QpFPIfQ2FSspu9ymYH/quQA4QeZ7
YSjzpC323PH5mxeaEMYDMSmOE0kEg5uo5LTRWyKTN/Ot9YcEOuBUKd0aN35URh2Dx38TdRwhs/cY
lTE+4YUEOh81zacdLU/ZDoMhTeNHkrK+5SxGC1b8LGnCV/fGhPM03aXndBzNO4ytYF5FRkPRP5JR
57kk6C1Xc6VsZrvUY81OJS281SbMw8XYDA83v6YEBxT0Bq7siW/Z4N+zSDmH3cEVlVWM8IzSZGlk
RtkHyjvEUM4YDNVBGA6JqCagjXuTi7GH+ViPL/JCobWssbI3frInm7QL/zq9jMppk+eJI4arzASB
OrECJA8Ac3iK+m4Uf8ixGyupVOoDd0n4Nv9UHks82U0bJHGCLjh8b/GOn6AQNgtkne2kA4p5rJCX
NPnwR05MzcqLCyVlWpx7Lmx7AkvUt9xueXAivX3IECEQXkZEczZT4VlGhsNTaaZpQzS1NFBvQA16
fPu5uCKXZn+x6esGNLJUDJ9+1EI73LLFic317yNnUomWKHwcrTD8ZA23MO+40gprWLQyjdfES++E
bf5Or3ONklAIsbJiV2Wl/c7o6B94KvxMWzRg8KS5iPIo++uYBrmGZy6ZntNgrRuNqfJOL8/9Bca+
Y//8j40Iz/jRY+u5rqLtX/D+HaCnpxXPg1PGx7MxZGYk3Rcllhd/TL+L/rp8WmIyDysYU60D1pV5
J03XMyAhVdTyy41gbf27cJc1mtOOVeFKgacUPmWzN+RktTd7WN6BXYLPWP+ap+7Fgt8Z1zIzmg9p
g/WTmy7NledUU7Hu9ujzr0WV1BVs+1R6eE5QXogEMuxVAdrno9RDUDgLNeA/Qy7AUTUEMpy6NnLG
kVEyZYO4bT0KbxnfR8f3H0wShPuengo+6HLpb+6njaUWPHOBMq/wlkuO3909oOOafSljViDgDDOU
URncUhaw5/ZCnk6XshFi6F+UV/ASSfqWSOZ6Zsa94/DBvzwm3P5SfrEybDOTt43SHfRRWDQokxIN
eMdRtH/3tU6w2XOZlxirl4/V19mPcmc2KzyuuaCAi090FgGkrLCll7QLfTVCc0h44KdVxpt7Y9NE
iZrhJUTZFJ3L3aGlVOZ3mWEafP5ZzhZkbkkIbl12OgL+oGxZx3Fn6R/UZgZJu+wVe1J1vl6Hx9dR
klQjiXo/hDQiLkBoaVRdtFiInvI+DNV7lb23NOvnwJU0G78ZrFZabFYIgrMIKKlFV9CoIMGLopt4
8i6nQuajuYbnboQHV6f59hEorZo6jzz/O4qr9K7dR3aUgHlLOgiXLGsJUOy+ByxRJWfWElGoSQxt
NzQ2A7rXSfPXE7Nnoyg+VF1BWAy7zMqgoFCJYVzZJp3TpXvaG+vLFicetmgu0XRukbFtkASLLHNa
Fc/KDA/WqNK21ybdVZYYcZsq/gbJ3Bc31iYQkEhQEgmWqkH8mhiJYAQlWIV1F3VrEx7QVG6c70ZN
kN4UqrwDSTNjc2WpHNGmq8YMqOppv3phPnMf8PenSV70usJPmYlBZrLTW3U9dT81lUzlKt419D7H
U3zDlSWxAAESYcHZPRPw33VaWSn6x+ll8NS+/FBLVLBHk/FNqTDDqJ2cqsznWJw5AdJ3bTVmu7hd
sAav4Tyv0cKS625baEmG1JutrQPWc7hqq4gx4B7rgaPGU/LiQAqEtRUy4SIKa+U3Pu27MTDFEGQP
HBtkl9R9wUeAtOROveka6dkinmbcD/c3Vto+Wnjf3B6zGYxFwvXlPKFnsuDVHwdab/Top2pFaI9F
43IEPvhrhP4DAqmaZHxVlVMbGGPA3DcFU+mbI8EC2lwZ5dq/aA6VAKgDH/oYR0NoRFQmKARZJ4+z
L9qPlOw+sOszu/WQL5pqJgRnl6EscQbbnnxdIw0V38Vrf5kS/WpzLYbFjoNCkdF9ZrWkUR4lcmv4
p4P7Iqt3lHZXmwr6P2sRcHhWU8bWVEUH1TwmmIteJactsuOULKiP9Goeu/k5UHDkwd0ShgvYvXHh
jTdZsOEnZQ9cERC3KUVC+SclJZMYWWCTQzyValSJrHDN7Ruxzk1qbpLJUYZBiiM3Vibl+BtoCTuv
7fJkCYk0lKbBWvLnJaafhhnNpp8crv63RjRnkpnPCMhdehJ5/U2na4+25LSaqcBpwA/SPPLX/LbY
yN9X6tM+Zwu7MS59MiLrjlIxJq0WKEhh74zIzqxfA05t2DwwlVSH8c4z5MhTeHdp2j2Y2FKJlySR
Fg2LDH9lUDOZIZccb6EzHpg2BWvE2JCYTrOuUwHpmQhTnzv3kymUWtV8jiETkzgJMC1FWbSFojjg
pV98c9V5YfrLMknIUqG1yNcRkJxDWrfJ8xUXi6evFhvAnBO6zl0cySbiArrpFmbASZ7Meqo7uvU6
FpIAms0R3kYO+VXHtHINsE9uzfZaeh9RfYzF5EVHUQttNQ+g2+k0/fGor+Dr7hOv5PUZgdp63CvK
N8gUmuf2ypTiTRNuk9susf+dSHrlfbOw0vV43FS8lrCzqQw0TC20qARy7JmHnIlnUeGkeXpxdfrc
clOZGugT8pvC6ViCP9nggjb0hOGUT9W5cT+njevsCr2qHsXkpeGmBo18TzCNj1htmHt11HNnkE0s
FWzkUY9R2z/6v79sQOIYtlooOkHqdbHLpMxOXtH65EzyO3ewsikiLx1HHzYt2QvDZ3ZiWqalOD/q
zi0hUMeOZQcjF4X2mY3TFY5prjWb0wbNYlr504xK+o7+UXbwn0JP9pvER/rdWDZI6NGGqvW8fVow
dCIWwm0mVIQJgO+BnB6fgLa6nNcY+SZ4lJsY8n9MbyLYzz+SWKvJc9pogrfjSPacZMQU5zTvsqDZ
1L+Rg+SXCnr2KnuJU/R656x94esucxIxm6+qdIJzq01iS5CuMySxlMe1tROKPbHQOSeJxFAj30vs
2TEFBCI5N8fiPgSzRRsMObFpmCBqSuBHe62nm6kt7iyjrmenhyR9ySbNiOH65Vd4vKyog1pUnTU+
ZvQWAwK0BbiBQLfzgNRBqlEEh9N01SsiojtBnR+N5U2yy8VvOuORZVCqilzTQP6c/pvtLSU8bsGi
a+ebZLLXLiUcQjlSYKmUEU/yWeUFO5HbOzbIj4Pqwqv7rGQ6N1jPOf5G8EcyH64c5dHBoZIQfgfz
790y5bo2+ponVIDorVyXTN/QdxFzwoiYo2w2jDsseBv3yhuqKZe0fZfBdyEYiKu5eKwC1yWvVn9G
f9zDyLepS2lXWHIuEmTYn30XiZQRXiCVn5LP1VSHUB6iMHJsVGS4Yu11aAj3xH44n9mSSOClsIdc
VLAUS616L1lfvfT4E9mBHrpb4Z6hGKHlAOKMH4C/P2F+G7B7Z2gNPGw9HkpLHIFo957/JCvIL0Ew
yzez1O1xcBk3opbYh2/X3mTV2im04FlEv72AGbP1oHBum8Mg+JkyzS5bEXacTliCor+RnbOg5qe5
NfFWdbrp0yvSHIFj4WJBClWSw3DDWQvpw75C6gql4YZPfucGfKx4G9qzbSaCqA/wFcT6dpDcUxiz
Ivd0lHvvSzJYhdNTh8ufrS9bF9B1ljTJn59ezi5zoXZ3RM8IqA5KaCadO62Tgn/ZW3UPW2Jh2eVf
ilEIkLdFHEx8KIM+5e63/HMg/hA/AVBkZNSCEtvT5W5kpRUMWK5JMpTgnY5peISft8qx4tyCpteK
FVQWEMJypvaf9vxcRrmbl3qL+5Vki/AD+42wMyYibmHnqbx7cgw87rpjvnXx8/KVH7Z91IWqrsHA
I6nulpaB7SrGHcX45yJZdsNTEZ0IW+KdFJ7GgufwfSFbO1u2jF1hhPkwhBSyFtUyFQcCnHDnnh58
27k40z4AWUjOPzLYqyfLCPswSLHOQbU5gChzZh0rFMaEyrIgLQQZXfWVJd6LcO1Ldc0S3JNFPVfe
aGsjAV6pMQda4Qei9DJ+uWbPoe7zHitDmNpQXvd2fm/81ZAuxg+8GWnbmuNYLmWRL6RTXZc9Qkaf
p6Oi/BDoPfjdRj2wTo9ghXQOOQGv7fwOmBYZhue8BxADuPWe2MRvV2Hl3w6bxvOdiA5kpi9w586F
YUhaVjTACj4quD2k1wHAI53ctCyWWHAc3YnmmCjYJbxCbWYh+CfXVv9MdJUDXWbHlkOWBFURPRu7
RAIJfBxv5fns7/saLi+7UxAoY1R0X+TAAQoBJ//qQcXUtGQTJXC/pnlsMhATnIRkYZuYr7kIeGd9
lIUMzVU4vynZlEAcc0KS/Cm6XIW4jRPYSmATdrcvqC0MKthhHO9PrdHnPYuBvnkSgZiuD15RMpBe
zcXduYnJUTZjIWuT5NTn51yszWz4dv34C+JiZRL/3I0humOJAmLqIIKyqFaKVr6QxFwxsSwU2Y7J
l3z97ajHvJHiEANjatsxrfYDuX+vhMts9tLl1qbjCvNWCWzZyWs8UkJrRjlBV1pPzq8nvDpIcjiK
J8OOMV7C/ng1p4UKyUcyVGLF3s9Lnp5x/ZJB98DJCdm4xZt6SQdWXeCz7HydRwgbGKV/HCVfsihH
fXUJjflAwPvyrtZCSh/MNwY8iVcNkeOdADwwpeVP7v02fHgP9GKvHHdeXcKerGeVfR8hPQ/Brskd
sK60wDwaNbVrpIBXvqu6BSMJe2NGSdVtzCaIPhle+Ei3Mm81xJA9v/T/49C+hN3RjW1G201zFYxC
f7IW6Qni5rKIRrJUdqCDua7LWJHUtJSLSX2ValQwI2h9geMGSiDgLEizq4sNRAJ2L2wmygnpSfyw
s278QUzWV4SnyYaAZOcXwpNWflUXa66DNHMnVWcNQtrVqJeM/18Bb/ezSNfiRE7EJ2zJxybacMWG
3KgGGMkp5WOPRx/aPH5qcxuVC/xYj7c3UlYKyYP/wT/quxa9yZGwaTx2Qt//RBmH76wyLqZ0W1UJ
QGQaASg3zAuEpLM14n13qF/2p59nPc5MIZ9DEYx9DESvsqcxUynCbHk3Nanaw/x3ATeRPlp9G7wi
6Hs7YfpnXTFlD3Gf6wN6AIjIQSOb22SJb1zgrdzqz0JoNAU0x03RAUbjCjyAlrvuti/e6NMosTeo
VRL7C0JVGjb5YZc4LPhh29bUwiDQoFrE050SN436/dGFj8W6gPLbgmWCaOrD8qB4CbWBWiPL4phl
BN2WcGJ+So1C4AGqwX8G2XN4BYvcpMnE1+DJAUQgha2ZzaWAifKh8/qLVXMHO6caDAE7dYt/oVBR
BIEOQny3Hu5nXYtxBizPr9zSQmns8nYUqnPiyfF8Zv2X6g6jFaa0zJpoldIZMH2y42gJjcwE0c41
IzdiQETsbTAOLAkCUfPZ1ce1Bo/YKDInkXYbzDPidK82HfFlNGa5LyklPDTg1v0MjOZk8AkANi6R
t9w21WabKVlRpdjXb/ilr2/Cwf/JCqxZW5NP72csyHmY6Tq8fqkTd6uisHQk1z5JLZBavbIE4h5g
eydoUJA4I50DHup/FgTHdOsDmvA+zc+FDwi1jDIjyDuKecG8mULkwQKL0c4chl9BGjgBuusW/+nt
S5T/94tBzmb1GUjHKPXSqWq/8iZrrZitTr4PPkvs6J2wyeb8Sp/RFI8/gvJ4nhlzsQgdp2Y66T9u
McxpD7tpqQM2W/tUjswcqIAs80mau5SJmLYpXWWBW2wmLYX3Nj4O+TrysXmSeoxVkkte3w2I5OTe
T6awYtppGeWGHZRk6E3wTD0Va1jwavAF3AXE+1OYbr/1lIiwAqIcevJUslPNdkMuaMRa+KOiZwI7
OO08CT6cS6k6YRGPGwKiVaAgndar8pswHPuGQAMBbJaaGQa+hYAJVn4b6zyjWO8wrNJBETE8kUUA
8+1J4BR3KydhdMcKgVLL2Iiusn6mYd9FvwpzS9rVB75ppryWlRuVTxoX4raNBbyPSEdlmUXpkrW+
k2rst66zalyCV2Q1ucBiPnVOQDzCasZVD2UUSsXyk/+aYIBt8BYSBe4n8PVsnhil5lQYc6TMXO/D
jnXZcRblBe1pWw9eT684eHzIZYc/rjszeJzKpb5uG19H+K+XK20GJ/acw6LCnFcMJUPj8YZisPwG
FKFHbtRVSIM+2W4L4gOtL4A647GBZP2IfCQwEWUsV2jZaCAKt6i51jJzL/zd8TULaDWn6KDz00L2
rr+02LKQzqNEVI8hvdDbwKPDYbp8HrqFy4f6o+5SNJb3Hlj5AExLLIBjMAE2XaNLnxk21se5d+sQ
HmCBPGm8FtrX4niiaVbh4EWLwDZSCjdYBV7qjav6zLULIXYHgH2OlWEUxA66HouzpHXSHSyWiJqs
cFvoJ12iu4dd/wsJE+zTvt5/8clv6TP4rWGf0j3eIvjmLMoVaosOmhLY9oXM3h7NA/3Od+xlmQZz
8JGrLYHZ9kQ6wNPK7sLXeljGlxFl/qUZnUt3SRK0rUwuwdIaKAdkTfH4Mws2oRMAj5/tYnDh3+ot
4q5Zx3eJ3LRC6gKwaWe8/TGoUNlTV9SS7jAq+8PyinF/N1IY1ZE+a8gu9Okvp0zAXxDV1F4IObuH
sZQ30x24yoow6XA+T3gmsgXXnl++06yKU6SEDIIbCAVfDsFWFlCM6AWVT7Q1QqBfvpBVPRlLn9tD
7x1TlOxPlW9jaSOMqBZjRa6gI7zjhLl1BGIqAdFDKomPSvNzl+EalQoGuuybERF9Uk/ZUNRJfGL/
xw0MJiKhAeOUV26yN8EGkfvwuf3NSWM+T1JM2Jf4+q4kMZYRDs25goLnBCMnvzA4ZD6Ecp7t0iZ8
wzmfeSsMKUbgIreNuX76Oopcd790TyS8ckepV25kR5slx8OZvzxwfM00kwcnrb3+jeq/WfKE379T
Ipx38NTZJ27KGKaTmkm+5ErS6cbBKc5khKf8jhbEYg3yD8SGQ8fFUXhhB61eq/vN51lkpT6mrlKk
PXTxK4msmEJFW2q0LpgUdh6IySYXkA245wQRD64u5CGt79zUSRpmPrpgyJunExR4vydEphhWWdBu
aZKGU/5HGj7R6Y/f8opfwbhwdyll96NXuCDbHtVnggbOobglI++tn6KDRYnx07LmgcRr+CE03Ii+
e2gUyoHq+co+A4jKvyqvrB+ww1+QPSNeSBTDu1fXz7W4Etfq9WfLAUps7xtB0A2U1prTrNCqXccD
LPkDUX6BOgN1bBBO6uIjhbN9P6P8EH6EflBdaExArZDUVioQtBnfLoiEKxYIBOvWE2HphA0fO+nS
qNB1ayMkWZgm4Ncyt9XiYyZaM7gZoGjnMRH/sJ3nRWhaxNpiPwY0L9sK3SEun/5GIIXfYOz2LTKK
F3ekbny2035z7cHKeIM2RVObp5kdWguXzqWrDLdy1MsyiyHgb4PiexcnuiiNrrkIjUsFkNiPiUqM
0Yhm0Sfus3iVOinm1qGZYJVMCSeSosBzN+b8ifktXHHpeYG+nmgMi8/yAyJc6MGfm4XuaOPKAp0U
Ot3RDQ35l77bswaLgqXMby/E3s87Mr8Zz38MOhFHraYwxcK7ZeXhl3ZBNguip3T9QTGEreSciti8
PSbqPqOfsLS+sZ8pTaxg/7rRvBZIm/Es702QYoG9SPLvDuk9OVP9HcjHoNNNcY1CMidORhFTrP1n
iE6yl2F2vEnaYZxyk2teRWHCPd3YQ6PEEBoZoyYxNqiCokXnpvMsZ7JXOIDsPbt6JSwzAZiv2iqV
wKjPDRzN0un9tq9WJ3anV+oG7Ykv1orrRo+GPAMBpkE0hT/bmKoT5SItTaKINXyQNT2FyEqkJf1F
AGWt0/3uqYDtfKKYOMTq2zBYiLhfkKmgPdNiWvVw/+F6m61jT3bPdrJwnbuUHX5ierydNno/3lxD
Q+/2CXHrGnZ3o5ETx8Wpp9G+9k5rMsmHYzUDdtzGpR5BIQLwpOMHBMk+zkFsXcJacOiaziHD5J9s
+580pPN5znSA2SKByN+S1BlGaZlylayrfqjD4mBzZs/P3KtJTLBpcFCxOJb6avEd7bPD545ng6/F
5c+T7GoWA09WPnYsX83uDRmu0LuVbeHfl6SRcrw7DLGEZWGSVNW4RSEqAqbRx68yOKODJjN2iVb9
g+TIW/XIsveh0BFqjc+BSzlUTWHCxNn2/3S6aev4DUokbUW/Vq1cEY0KALXvdrtxBUC4BlPOYoFr
9wNw9hctW3sC1qyfeWpBJ4Oxkz/GYCwGWI/oYiKxK3gRhskGniuwYGF2ZMdQQ/KcrRuD9nxroLgY
vvVVVCKZWDAQkO2WS1u1xfAQwTe1n3fDbl4B3X7Jwb1jwwqmTUDAQQ8JUUbQT7o1GLfGW2j3TShH
0qTSHtrmce85jlsOge5sJTJbedTeWz6c57SWL4GP5t6yTHOFm9Bnb/fuAZw4k52Bcg7Wlb6++pFG
8uAs93/U3oGBDkq/z3PrzA28wbCYSz/0IFRczJzzRywya85YRf4NBKEnInBUon5dDe5rRqa1RYUe
k77uvlbJGpYLDbcQoUw1WO1lufA8oQ5uQaAK+JgDz+LV0ywKJUQc6dTN8GgSkIr4pkBip/g4Lo2N
8YbQ2vY98xWUseeUVUOjn2tSFe6ydk5WOmRuxvcZXO3wmDhg8OzwGGkRJPIASlAryzod9lGRAQ4E
2q+YXS+AGBWotIXeool/G1XnJWkqYNNjjzF1iy2bMlSAMisZ9m8c3Ol5+gnC08DiA7BPg9oGpOc1
C0pzerlhlxUgIrbQQlnJm30aUgttPfo+tXPTPcwMy/yaIheJCCQJ5FT/zJ+/epiviN2bt3t+q/Xy
UC4OjgoSIZsQNbknmsH2oa9r9Ucu4N9PiPjhKPSegnjf25LSzxMwzGJD3lbBkhr1Kq7+li+Hz4f9
TQxqRuPQ0a71Pdm1K+nZ0jU04dLpu6mPxypBlAQXZ/zznKSx6Vttwpat2Vmzb7VHUySvwzn9krrH
oHvTheaxOS757sqi9JVmr4TNtcekpUZ7iYVGq3pSpXfwYg5HFesKKwmWKsF5+bSgEyLVKv3zPxLn
UqkKQ36ubc2osIwI75q8sF6bYqfGx7eBbqhKhAABQ08xEAC1OlwiSMxLGHyxfD2iO1CegfW4ErAV
1iX6svZmPWgLoCzpVtaLWec29SPQe9ukJiljwri/9lVJVQ9tOS7ogXYh6x0b+JiHPRy6n0QjXpF6
G/9gW6udc40rnw8mVyz19ZHolmI+FXN/nl/xTPsZx2gdxjkJ/c3WaiqPLJHwF65A9ZYB8J7rQ5PH
W5NghZGjWVJNT+ctHk3Q32Qluabpt0nhFbd2XlAzAStG8N+Xu7jOUTLN5UDLvKhOmDAeEa4OQpPs
kBkt8rDmvPI+ygLx/X8LLkTyQ8KLo85FO2K8NiVs/wettFyW5Hrn1cERwDQHgFHccvRQHqtLLMaW
g1YgL2zSI68rwvWI7khP8oTR5LQWFyu/9rWSYpGKaAMiVO/Gl3uSzsus2WGgH2NHdlcaqUtE9UlV
S7yGHftErDj5wSbWjBcvzA2xZm9QpJmtzdw8/KRjJP+bogb1PFgLwaw3WabrKUMsgWpPkONOqwuR
X2NdXX+aqXSYSQviTu0Ne3qIwSc7WHCdk1VsiGYz9UduX0J0nDgt0ScCSWyxY9lROFWjd2Jan23x
PwFU/USs8vWUJu9rfPHilaLPezlbwaIO2V81Q4SkyDQPlt1j+/cnKHSO2ebrt6VSLUeCRo+mfzsp
1Tu9X78YF8dCrcQ6Wx1NADaalPuWeBOCKEaB8K38PBFBUO4MXS/sPwRQYNn69qGRllLLNqUbqQZX
L8EwYyinngwjYiOmzZQB/7DMn5CH3qobyB92bmNXFNlvfG4ppZ4L01etJFYJdFkH+EamlKNH2UKw
/M54bKbSKOHLrUlVF3JEPT6tBGvvyct3Rhc8kbjSJUj1dlxdjCgA38ps2Nv3kgVcpVeVFHIJXRfz
3xiof/cxi5HNyIAJ1jqkAWuKYcV66xTBoPnw19fH1NmdiGMZPCB7opmqtkESJdicRol096vlO1p8
UDKN6/R0EagLzxC9tPVDijDE7s1FQy9qQMQT7ZBZJuzILa3zL1WhllPPK4S4j7a5jlVh0DYaE9D/
SzqptPMERGaTrttbFow0yWGCD1TkNGvhKgrYO4AHt7kvH+fe8pcroxgwAHH6VygIenPEdcslHfM8
A1ATbaeTttOg1UVOppGzfFtGwqayqtMoW8Cce1CEp/Ol2kYkhgu06VshEzTD9tBNPivhiPXZSPUk
Dmv7SXmDGv0QzgTl994GUdeW8bUVYs8K+lLR1DmAT7i+FSDCzqlhIeOpp0EZn9DOjXqLzLcOV6t6
6Gfh9nzxuuOM89HapScftoVj8I4sPXpMu1ks6DSCM9MIYxLZIIBVWKD7E9Hdz+b7ZgNrAVONgJoD
65pXqfK/mFiY1QiMygOONTP+mVaEWz29jm0ObdTVS03odOV/UVZtzkDYoLufS+AwDkbH2nIny1ZX
AGT7qx7NMIqC0h+xyQ9oipok3EOconn4O5BGR6jtI7GtrVR4Ja7PghukzGzMdu3DWqSMyNvq+ab5
b3PN747JwL+jz6LhPuISWbRxVrNU5sBF1WdIaXxH2yvTTRMHELnoYd+A16fV2/f52g50+LGHuD8Z
TPrwICxaJJ3KEBaUqgit4tqD6/iYbpEyG5RlIWR3HEqPdhu3sRyHu5+nmSnSC/GGzza0hoV1SYwo
sW6rpuKrnVVQVezEUJjqyNv2qrciE2EwzKMrQVnG6JNycPl8lqSFDZW+rIDe3coWRkJTZl3O+MXx
61aS/mH3WxG6BBFhklMjG4ZvFQWnQXxV/jqGlAMuElQR5o4nCxgX+qVdKbOkEg+E8Tgd27xUQ/2O
5SkysO1aZzJJLRO1j5Cfhps2Y/mXQAHOG8kczXkETQU6A7239UhGa81U6mmcXfjTQlhab0p8MQ0a
SI/XXIySPDlgLwTSQizt7gk7ugDGGqQjEaMDkWeLr69pHNGMqrYHTjR26UtZGkGoaM9c+wUjpsHw
puSyYXWv6xqgh86zfVLhWDreAUNNclNzD9lD5+D9nSq/dzhdEY9Iz3ic/LWvE/9L5tA8rNb+mcZU
NVLvEs3I0zxNYxaWh5Iru8WNHSj/mK7uVWi2LHQAZZ9aKI17FlsWokAr+NRXZ8gQAAS6C061DeDC
ujZJcrUUi76iO9faURskRuMgtJMvOnvu2qursnEs11udX4eoNWajEUnDztb8sdkYqvWYnCDScmFD
lF5pt2OroJlgVuXSlV6eNuwxMV9HbkEothmZsax7VSXCkLUpHMPuouXE7it7pnAPvg318ckIGgF5
Oa5k9DbUjXj8379eLb67QZjheqlaVIP7H1j+ybYbzrKD8+crhqwTm8aB+Fej8ZVHPoZAHiHVDpB0
QVy3h4pQjrPx455j54uDNK7BO06e0cjwAQghltraCsxVF0E3ez9lVhIUoYadyc5fouI3LDsOAsqj
hIggVeDV8gwSwVFxc2P0eCR/GkKWAjTt5UZjUdUet5iYtd6y/J5S+d/Ds9n7U+Kp5P677Sz+HBfe
8MpKFFIZSuKGRX52edi/1hidoUO9fVAJ6IpHZ5Q2A3wu8gP2MtrjgicphiZQhaoI47K9Isa+m1Px
tVBJblSSJiFgXcqUfBtFgn2ZyFmnKpT9qwtxyKPRT6ZpSmkQToR0mkkGdexyvX6R3XEN9CeNW0+b
XvcJc1zpky8mUXwxSuGZ8+JKIwyf9Krgo6Z3xTSUxpJkwllh0Rnx0Bu4pnVynTDJrSy4eICj3ukM
LUv3FKmubm8SmTFLya/N7p9dA3EBWZMuq2BnpZxycXe1LRTFLvFakvvRKvW2d06vNXUl9h2stitW
sZS9/bRR4Nm88N9u08fnOOEn1XKraWbJPBQCj3IBWY1zxam6Xt1b5zncRZCad1PfBYZETHyae9Js
6iVqVeESgSscFFO6oXk5OUC0EBCxNclHY7Kl+eBrN+SUeWFNXcrenWJpR+Ri2HRyEjA/GTREGrYK
q9RRcq4uk8dnANEPrMAj0l0SZwj4LcgAgMKZrVRg1oh5X1r1Fwen574g7K+KxOguC1b6YdYxHpJB
u8YIIeROIZWTUijRmEV5RtBiLcW2DpdZ22SmP3skWy8T271FHHvbDXB6noxjy8n46xks0a1M8w8x
NIpUaHSeR6QT9caz8lTYwjFGX1FT94yHd6j4Te7mVeAtSNhsqnwbdTmbsccAF3TBF73X+pM+9Ix3
jUy2R5hkubdm6dP1W7ZLgyX9ywgNv8QBGcazMwqVyEwlNPWqERfLMXTqQQh8qGSbJ40RRr4MqoFA
qymVzrNOm9jv+A2FEDUTPaBi521QRz42PBxZ9YfwBB7p0rTQP9SCcwKnXAUHab9GV3b4IKPcLMp5
+GIQ7zCuWU6XZoiKnxGauGM+ylhsLIB5M2qvMs10/Ix+GE9v9GiPCAwXzUfp86aEaJoK8Xkl0Nu4
o47oHONIhGomRLKH5I9kIusdFw4eKu681srMrCneY8sCOYusdNIzEpEOMdEy0Pl/2uZgMveKt2fz
m646/b16+vqRcBJxYdH1GTv3eyc08NX6chePoJbQp4s/OH77XO6fOSqeY0mo1ESSqypEJ0tm/iSX
bq52GCLkiYN0W6xnjSKGw3n42FNJ5rQXTQ55kMxGx8FNHWEKlAVSxhJJv805hAxIQH5mvuNZNUJb
Rso+x1LZQXtXGZ0zii5gL3TbO654xO+pmQxKrJfQgPFmbJ3ZmilVFyt4GQfCdCLamIYQqB52YQQQ
54RLeh5HeYWTazwxqOo3YTYUNAbOdU4KO6SXIijKfStA2Zc6csngHxrWAbEYHhZ38xgy3vpkJd/Q
+rpgwDEjUwDKowlaZuVCUki9Exum1w74CorfIB6pDj1BCFYpRK65vnE8fy9Y35avqf82ktnzysY0
APjGkSC3WwvWP5kIuzXRRb4F660i7MBU/fNC8CdfTOKTjME+5cxkTCsOdDvv068ZdIXYF3J/YIAK
LZhxb0TpCoYPzoDSlea/eCdzGLIAxprHJtbV+xeKyuYfqriacRcLBpwuzJllulDHrigkEE5GOPrd
IuBUWZW2FgwIPXC7ls/SVAX4vF16TBGwEA0lN0M0Z4pNTCAjw8lCktLnuJtLgZ4bmO2Dv1YhomIg
KPXc+TC9HnButmBH4FCfCDeoKE07TdSBU6SZunxDZ9d/84nLICKqsO/MGS7LaJz6ODeLiY/RmjfX
YuACDle0wWyVRDAEYXEUSMfQJVh3miecBl6IldLwGSuOQGrGTgccuQMFuFGM/uTDmqTgySndW8XZ
QALMI9ioqv4UcBj8WVucb7L08M4tR8BSE2XxvXlwBt3v1+Vujped9xeg3pGCXYTMY6u3xofyPN7p
LUqYc+oVq+LYpv2hP/j3KQTiEWjLnmdFMvhI4FWG2WenyPn4eMz1JO64V3OCeSQa4mizsvijH0NU
cJtZZhzQPec9UFMaS+1ns4gYv1W4MLK7wORIM5xQHC3xCheZ7sH97pwEeXhM0fGVXKRQRkVaYucB
RiEt/2BQeJO7gWbweRhn8+BDimDIPzybp8mCFmu5/JVOT/dnK8y+PY5RQFTI7+2lpMJqkymkk+Ws
TzQ0io2eZ2wzRVls6eFm9AnexWKRNMX27dE9TKDg29FS1Z6Bbb+2kpx2Zim8QIYxcLGl8yLkp29n
tpISORNw3I6xf9IfGWSQsnQpa7bihQcnVNounFVPY2Sz8yD4RyzWDwc3geNTlCSng3lIe9u0cFES
qAcMKQ9Qazyh8DMB0jTU+q5qa4loTKFrmXCpFYbXu77uC4EHHCsipOR15oSldt9Fl7eZymmK72+6
1K/Lui5QSjRgZxlW5W8jQklHMYgaCYDHCRtsSy/75cuCx0wYG8CotwtjxoDchjFhPcgLAEYduT8l
zXVGnnm8XkUZIXklSSov1WP2MqbTgr7jdICZhL3IMdqVbSicZ5eaqf15ZP+X9qYdcl3uOG3SMIxz
s21Ab5TCCWWoGIPwNKowtNu5uBWCRwHodzFKzX//UjCVEvnNL6DbNfXruFd418WXOvPLn9bMX3jd
hGCiJ6rhAMOm7j3VrNjMAXLWTZxqeUGwYqKFxBF5mg61WqMXCbAcQ4CSLhdhbVDirQyMzA9w45nX
0T0EOxJ6JWQBsmpSGKIi0LlIVeah4wqGNtnU0t+Qgr1o0PUJkh7R/LsjpWYt0/GMYQV738F7W+5Z
uER0pBdo89rE4EfVrFTlYZeRliD1qsl953ZfZjCENFaGQzl1f/kgzoQuAbC4w9nIqKr2NqFYmj2/
UhYzNZmN19ibolI7tP7RmKn2gMiBkUNjHRtVgwdI6+ILNw/J+DCLraYNmPPIhtQL3+vLisV8a2EZ
QEwdXPLoay/srQfvFifEcSxPYYprt5WRx+AKUves+fBYWSDZUwTBh4jvGGAJItQ/khcXKhgu4T+v
hsMzOzQ1mmmSkxD0CBIjEebLvfcRJImXi5MHPybYKmMZJqcORLqkxJ5wnFNbAvIs3hsK7lHd5Icd
YPvX3fCcBIjdyz1pWE+F+kMvOrh/QY63ckr6l3YCxQMXyEJkKYvtOSi6hWZ0bduT3NwhAVQx4y85
rP9KH1wntZq3RER1Sc8nMmAQfOxhNfyaLeZi4YskXxv9Z27sH91YSAd3hkHjo9/4u+QZPAR52IHh
rpmLtXOEEZ8qdEzWhtr/BvLmBbvJNdjr9EdoQb4PfwZ9Eq/FGouN7nOWDY1iXlf2xnG9V61VtCIc
k35OEc3V7ZpKLwE/OMag3PwIV0L7DlOerWs5et7vqcYvsCb1EDZhHFc8rJ+Kb9TvsoXIRXJaHxB0
TbOrj0PEh7IYnRrVeUCJZsojadU/H4tYz7UdgEaeFRLDFMaZu4IXMAHqj3z8JI8j8gYnTo8EEbkm
xqbvVh4JcgwRiS5qCU6rvEeQyfmqxZVu1gR9nDjyFhdv4hGdsdsZdbQ+1xNFavoamaC52QsCOIia
MOiiAho0qSmjeUUFc3N1hWcDDohEQIh26JbyS0xdi+WDkNLvp8MEkDdMl66zvvtX0YVeOFefvQGW
E0/e0xCdEqVWlyVn2BGrFU6U9gCWEsGnhg/usH4Sf1tyD8s00Tx+NbHOh2KLBZ7M0cHwehHZQDru
l7+yP6DNBg0JaIQNpU9ZLKr96G1fVg0LNQeTIpWenXbzMkWrAzt5fvZ6xWFTQTu9eQ9r8tWGpdV1
sPfEMtGriByzKecBGHn2kqD3NFBgvY21HmTDTxCRUoctBqweNxMMcTFqTMHA0iKVFDRz+mnEVpQj
DMPyYgwDkIu3CRmBi4G8tvX5eMMlJsdthQWqKG7USpf58RdGzFEyDtkSD6Q3jJVfkK0C9qAi4ANd
7EdZKnnUUeoulvodzRVBCZ2IJFefpOU+S5+UtPqMa/C8j39UqTmGq1OwNyIlmWzUClfkKAQczjaJ
jd0wxjnVQCYlpWvqg75x5ASlE6l5vewde9yRin5vi/GVsSAj7nV0TiY8ilrqrecX/tewU7FIEZQ5
k3h+jLszDHUxWTanWW4542q2srkMVtzFRtWMcCmWedWiRXydbcCczKwVxLR7vzCCz41sI+8ZYVbF
LcdEHyo09SQx67odBp06CLtWcLoPRA3+3IGPk9XfpS+AFUZCfOffZr6NNhMq2rv2a1akZp83NRoJ
Jb+UzlpKGMaXRHLrRznDFmVxbj/Kkt7jDmhpmgnGoirYETZ4aSJoQlnqFtOhCPjpfCJMDPnOdQt3
iFnFehFPmgMPdu26JwWHkHAEhpqyuCzDP6R394kMJx8HhcCRGoUwpp5/WhyJ2zTGKSChRISgkJe+
b5n7ER7Lc3VSlgXOmX2uGT5tXaTLYBMrjjY8eWcpbN1iHZ49JeezF1tssFS0HuYkf7iiLPd7qj69
UPT44X3yX6Yp0ZEDIOYwYGm/U3uqD35IWfDzyobmfzJ6OAJKayHmqSH5WXFFpRJ5SoNon1iP+VAx
0q8snTda5+OX2krqQYdPRLdIjgW/2p58btwidktdgakadygM4dT+WBb8H8f51h1jZqQX9FZn5ngr
e2ipOe0A9Ok46lNCMXE3YFY85Yor8iQY7ZDm7XN/8lTj6iMEe6V68dNpTLjt7mawh/EbdRf7W0Ww
rHQ4RBmcWQXmRTSH9YgFn7Qp7UiyYPZXdk+46ptX0IWrGWgtlffttTtPeU3Y1asv99AvN9q8HpHV
SKdM40NStlHI1/CExK5TAno30aRAc5DwZ7YIfjXMf+w7fJg8aUxT6w/HrV9vZGxsOzOq5mFwB+Rm
hVzIx9OlnslbSWchuSI/l/iFyvJz04HoFAQj9yyK3FR5bA48FICVGT4ZROnG0qIynIFmjMe5jczm
kiY8XbkSBwQcO7l0s6zi5WDy2k03kTM4PZcQ2vgxuyNnP4JmBKfBYSJSm7wxnWzOHtDd1udat+cX
duKk8oKUgpeDJn+Qgz8/FjIa3FHdRTSGxyF3TyzkKk+uXDGVQXxy39rT21x4kXpmszvLnfPyb/a4
MnX5n48C09U0j5buuVR5KiazjwD6vO0L2bhTD7CmvOZz265/Z99MULKo8QlOA82wA+6I+Lb4ckdU
hKZFHuZJlKzJNfxw2CmHVZgzxWpGQGc2/8i/HZIjEU3nhk8q8N9SICwNS7yR6yqfVrRZPAeAhrGy
Hk01qsz+15iAZTh6X4kkBB9Z6SFdsty96snNsD7MMekKPDlgCT8mMh7E972pyOxUaNZtdGLjX40B
N9Pq1XgiXKVav+JRrYTQ3A4G4gFPXa8ry2a1S9XVeBpPxcbgTK3yWzizLKBQV1x8SuBeumJj/kJV
iVdy5YVPh8jQrN0HBXCH7MHviiP0ZnJwxdfu5s3Rr+nCx7qZVLTVwkBBCWY/Uy2OPvAq6ob7Np/l
+yKQC4MHr0rdyyfAMI/j8LhNCTIuHJTmL/OUL4bsXb6tjnojz9kLdHMZS46SWv88XnR8VcnFTkzG
91qDnHRoNgJSfzcVQSXfqsgZAi86oR2HTR0at2fxNNult9MTyIjNoT8YyUDmp8Rx8GdAhERZu+1Q
wz5SSvdKNXK2dFOOk52+A2ikKRffxmWaga413NsBt9chpLm1v0Gp9FpKXIUqOKCd02PCIiBW1RM9
a/WGai7esJHwEKlsVK4dLgCXxeb8lzhwusFDUVZQdrPrOtswXXjGKQgHKnyapSFl/BjemzBwRNDy
FCE4jTRcHawjVC0z5DXMLXik2ZCeFou9WtjGpi27iZfP2/Qoe3KxTxv+sc/KQ6yXmMjQ0RPUfN+a
Si0wqt8BdmuufBPrQPiWq8fgIELQ78w6I2CKTivUzYqLBLVTyoAhd8z0ykq1eWG7leOM1gOPMhqw
Nx2lT2m/A48rgjQTvC4F2H5sgpXKxyoD+DXRAK2kZS1yY94PCaxAYgboU8wUZh1CTJG2ZVFkZTUI
zJA/F4JMic5myaZNS5btu+8Qr/2J+fZoSA4spGuEWUAxIrIFBHepvh6WhfBDjgRwiMVGhY8llNDw
yjJF2+u5vI5NZiXjSs8mAVDUIQLmYpkEjVCnKeI6isYOuWz2Is26aPQ9ZUgJn8IcEViBnMhiCa2b
BXqxy/Q6ZCAFS0lkmB88E3YQdq0INy06bo5wfSqP3FGNHrQrsWoWcZ7Xis9C8AixkVawWkXYyC5E
rCqcUpbEQsjJr6bfz2XghigbZesDb3OvltF96Ut3tvwHMmqF0cXCHMQr0VCoz3Y8ROxO/8HAjx42
2No1bdZUxuGQzJpnWHrtmuovdEiMbFSx9lydRbsH8Z3PA3J42Fl3GZhIz9gujG9y5H+AcPGHptgI
6cEOBuwAbbrxm9yy2cKb54YCIu0QaTCP2PkvOnjPqfinezxZlhbqszP7P6VAz0Lv/3F0/vIGJAi6
0g/8tqfZvwyS2UGAqdUAE+oRAjXVVObooBwH+JnOy7fBDW1PQejKOIt9sXz3z6se0XyjKyG8ylVL
4LRIHhI/DwmSWT1+QeCFHjEuOJj3a9ssGU8rxT7Q5gmdBP0C2840VE4jWZRmpPj1Sly45yL9QvYM
qQqlCDP70vVlh97S8NsFTk+Yrho3GQa3tmubUcy82DS/59Mth78dPh34NZ6OM7i4rmivXYulFxXm
8RvwJL2G8lvId8dfbJM5kFnUkDDkNR96W1yRdbo9jlnwc8KKP+Bas+8MffoMyLFhZfJo427t14tX
xG8XNbYx5uGX8KBsW40pda2nskzfUWgvqQeWbrTUS0Ghhjfd+7Vm7FPIXI4NDMQH0VZAchxKa6yn
N6VsOau5EppbB96tsCMwnYBJlzSKGvaBja10XJ+5CyMNmYPEsVr+a55ivoIspCp9lrC6EbcV6EGB
t6sHZOucqvFIxtvYeZBtljoaTFkLtGlHbY12bWI8HsH53mbgWX3smuKmzjlAIy0000qXAjt2mTK7
eqY1kM/auEX2P2ekwxSbCmde9JAyGix6khlJkPfQ7NHNxrsS5dOFAt5JQ1xGNsPloW/urB1Nj+zB
EPX+ThMAIP0dRc4FHu1AVERXTMdPKk7zw+jfSr831roLrEKv/OM5PEKZSq0fYmOEIFfprG+JD2G4
lw2xqEK+G/qVxHU4QhF69pqp+CpX//xs9ycLzJJi+V2D6Lo10kUnEjdmunH4oumP6vHX6bgkWDj0
oLrSBTno/yaHLGDc3Mb1ZH7H8fSJdgiRwyNFpRMLmul5KcPYt5Qt4+fmPlhTCfOhD+5QUkqcxRYl
/O+uz+EAiCQs0124Y6ezex0hMyeG39rm1mZXYGrfrfpYltuTrfnPnH8D7XxJ5XzMLh4i/z3EXs0I
cqwWGcXhhkABdXA34I/q/HIlSeRkW0XKupKb2tVJLRTPvSlJOHXOZAuueDD0Sxq375EJOV7RyuhB
/972wJcNq390IaqyMxcktxKxWTeQfchZ5m1Ht1JOsK6LWEsUnShLKzJbPAovzHU/aA3SHb7rweO9
RQEWKa9LncPoeT/cpGSFLmE3/pXGPMCBSkID08Sw1iV44Qnk9sMeYy8EM7CTXRLbUPKY9pySz3A3
nKig97aQO9Zhbju1FsgLq+rNA+qKRjcVZpf+I4l+tget92FhTeApbQ8rsIrHjxqq7aDuhFGqGWvN
2GUgnfcDlE1UisrG+MdBj92qSU/7nvSdxomuze479M3Qx9rboFGOJCKva/+kUoxYdcR1zkpLCYCj
oeUc+fUbJVWebWa1iQHrq3HfX1gcvRqfL/6DMWSK0evs0tcsMXUzVi0w9BxN1OluxAJ6s78tHoEU
klmD1asId/UFklM0Tm/iiGYGZuAR5q70x4nnoxVUIPjnF5nL6RCKGZ5NlnOoPmvpP2VCCn15o+4b
YMDo/fv6ahkuA2y1TzkIRvBc5pAiTN05ETDVqPv1gaz/ZFB4eAFk3hoNcN5tkRw7fSaOg2ILWSXQ
6gxOzFhttYv+h4VWMooJrppYbazBERdyu2r9efG4qWgAg19dyI1IWmpiPmDeKt2l1q42FrwIklr7
De0+HRKc++RiGUJ9f55LvAMnyJwfMoa4DKtMfKKoV92y4p+oGaOJqkWAw3okiKSA90PPSdJIvWuj
w2gQC7KShTDPvm1Khmrdzh4l0bIozzvSbDytOUtqisWZ+3oj5kK5YYKXv1duFUbyHRZ1M1UsyaV3
ccvr7be5nv73hbHjph+wYBIfmFQi35A4+hM9OG4Voiyytb62xsaV5kEGASRGbgszyNHg0vFfRdGQ
gGk3aPOZqCw/GDFrv/LQxnC4y0otwjPIWfdlEqaYEqreVfGPrFGtuRdeYV8H2uMWFxAJfRFOh00r
LUs8DRnLvR1bykon7ekKbs9MWt/L2NiKjjZS2ZpJBlhisndmuZurRrrrZL+Gpc1gOvpNI81yVvLU
dQ/iYUF4tSp0PzjqH5cXjOM/YnCFkZeAvTFa9dRFUUHHQoxDS7b+4TkjL0WqzAacSiysXUBleVU8
aiDBIaimyX3F0z7qmUAxNFkHsu3SWsD/Qf3v/ZdLXdZqQ/54KkvfjmZsZ4jwDTDd3BrDdo7pmdJf
Bd0el3k/sK3JzU6r7aGDVSJ8DCKyeWN8YflH0LFEX26XcbbjvCpqkco6fFvlFX+S/74GPIv5Tbfs
sazjcS5oqh/7ZRJnFAaC0STy4NLjNDmapfGGRQgDqi657u36NGruE6BRdlifdMgDMkCddXbQVuvw
reRxervUH/ydKf6iYGa4j+t82PHFXcSaRhpOTrMlRnKHIAX61oMQRsU3fOAgrW0rDpfZtRhRimTE
pJADxWMZkOCD6MVUH3eVCEXMk36y2r4lJL0nZz2CwC68zpTAwFR29OVpqTPuZbOFeogIz5Y8w2gh
CwhV7ZgKL9diAB0N1VAXI5WcTrGs99Ob8SqbZ+ISzSN0SuTPsvPbCeS+eaIJSDwkwwX62SHNqxJY
o2madfFRdiNiFwQhbkJz8RTgCFDpazY3Mpn2s5KQpZtX/Hh2YuNSfakxWB8QYszCI6WjoBBwMuds
m5Qy6V+uavgoCstnXfgrimuFLOimHEjx1vbxPBnJ/DT7jStnAJh+JYPrg6MR/l1Gbb/0bGw5OGRl
W+2JCtE7hAkH1g3p94Qx7MqEDOGbv3awwI3rVk65eSiffymLvkF1NYU0b2WCGSxyDL8/2Tg09V8N
aSAxo2W9ywxZJyGOYOaD0BQ5pDdyW4BNDYOTNj0hnDCan9xauRQxJhJreJnpDtCVCwMbNXLUiEKI
k+dY4GNHnfC5zzCqfxBcdkCNY8bLL/ZwMWmVde4wips4pnKPsAPno92gA+6dqW6f+ym5cg8a7RBf
zqGK09JYMPbOZ8COV4hG/SCVF4Ajjngx1svN6rZXW/akSvW7NZ/xkkxiTTl8mw5g8paLQOY6zIKm
xvof1glcvW8nW3uNFmFZloysALBhU3+rTLDfIZcAqFf2fbaRNmfL1u2DjZryOjluCeCrviaT/KaT
oxydRR15YnyST+h5UYlz0P4avjhHMtWZ3BWasPBeLFt+WHNUMcH4Btt/0Wu2zc3JEz9NLvfR1ZnY
71GfKfGZ0yUh/xusUmWjUsGGelQ1m1aVe3Y+b3tloT/mfYCX87ilTuy8NVz97KQsMFlHx4mylhg+
eBVUftfV0EzRfUdK9B3Zppl4bNANMb8ZzWtMUFveetgYdTEx7ZJyREYP52OTb4x0v7RJmxuUvodY
iDUE2Up8SFUVflJYlu3SpAiB9sA3OzHYryp/1sokonwrwftuJG+s76ZifnHZLqTwYweVLq7a8NMC
gGH8WfjHiqjPmGxR6mnvrSfnVcPsIrLXg6UiWQeH7LFUH6QwpyfQ8iFLE4bRA/O0Aag5dsgls2hX
k5CZKaSBq5CEIckmyO/rKXYNZ+XAJDL4vFNSbK2fCFCBcc3Xr173tqQRb7my/Wm7yLcFQBbJPL+r
2PWz6JzxKowRKTMKoNAl9luD8zZ1JlXwf3LFVddQW3r1+pe3EOpJUPWVkVbJQwjRvx95EqSNeE7m
FH6i5xM6V4+PNrO2vuB/+OgpJslVTTMKopEgPlfIUwd/7dL88AoC5haQumCx2Iw7IMTdmF635uXQ
KAl8CHLTPSEXL9vk/XzrkITFb4VVxvpe5xXOOGj1K+RA6WryYfsca2aKBnFqK5KvNuuvbGMaxcJH
tvhb4zykaDK6SOZePIlO8aEoz6wrcgRGbB+hoCP9WXg/Nq6lchdQfJpSVc5hUhsWQphAbhgB28us
60ywcT7847058g4ib96zMW2VWjtnwzO+sNGejqCSiW3rAr586bSXsjlsz8owT6mzR9UvkcM5I+yb
JzBkwxJUyqBXcf+Jeu3HkvnONQrlgW3Mm4/V2QZr8fLhxSMhfK923XVrGqYKftUv3zDbAZ6XKqzV
s3kC4l+4AWLjVCE/bIjhb2hiPcByenkAiUzUCSYk3IXGJRk+brMuPQ44X56020DlVa4eYDo73my5
rThS+3RBXNp8aHe5p0Dz3beFQsryTlOgnK9GF8V8cdFG15jpwpIzuKqxQZAWyuJ/esrcpfKcR9EK
NB1r/J6CWkZQzevXs8hPQ8l4rd80fgc3tZNryBHF4WsXeW1oxXKBLClSXZjsfKJnbNjywiNx1G+y
uWMygqtHc4VGxBSERdw/Rbg1kkMvfRh2zIYI40XGfCe9c62YyyW8VdZ7lWCeb5jbWh/4g82J7jZm
yB62HMG5WCNymY7LEBKQ2gZuGUmqcRrqu2H06oJBURhHKgV7EyvupjkUyuSPL4ukxYYkNc72r6z7
5/cQUOD3QNq3iDkdXaAAX5GazpJZ49Cc9cpS+RmlVe0VUeNujTKDsYZ+CXKV3baPqGfvz1nMSP0R
fIIhGZ1LOM3Q79mucJ6ek4OamfMR/GU8oj48c6E6QtJ2fhuavhv4lXP41IGP4YFTRbhuI8jWJt+F
D0hsXOnEz7i4Mux2k4MQ6IPIhJJT5u8dKK++eI9HI/7n5hWrI/zOg1YP+JIctFTqNSXYB4I6Vdez
JVK1LHtJ3ad5dr5nx9T7JQ3NWB5HOOFK7grSYi2Z7XjmUCPDPIr+A6xGZ+TeXrewn2SmOXUvNHDg
G7d4e1N9DQ86IueYviD7ItodDq1J8x1bkz4B0BEAMS7qRBnQsWMswZejkQ2tyCD4ID1ZHfNJKXv/
rVxBe+aR3cfUaEPldcLf0/AhKjQy6s6umCIOb1AYDzMYgEgZvlTJrzTu+yQUxv5LvXqVCc+GH2qF
A5UR+ke56hXqcEu0yEh6Cyayo+pqx/2R21kIBZFjtNAWC5rU+qeH5yFwP13fqVml3nJTWfcXn2Ew
NfMZFErauCS2MTFHYEUW8W3m/fWEW8FZF0RjF7GGjR6bhlN68CFdJzx1JWn5Cqn6p/Vr3ZEvggaN
XlDSxB4NrRSY+IhShICx++3wc/hUhjca3ih68sbNzN/Pkiqz11GME5Nv4iURANnys4s+i/ggLT2D
nPxyQNuY8nsxbLranit3et2vJy3Vbt9BPlsrT9ayx7F+zLEFzpOhArqkuXaOVhrFgYMwlzq9V1b6
NUBzbreLsdNNBvEwlI0MImjrRNZu4h0c9ZbQ+tCoaxLbhY8HqaYlnhzzh6wCktHXwkXhgzEtC0Jj
8SfIxkg+BJ3DZb+pKwLSx23SmzM2qAk1OAocrcJtxWt2RDIpjngfMG3GgLEsI0ClXEVXfIYNBP/D
V+IBjzXeGFJmXSpGihAnGFk0HVGhkoR//xhvJEdVEx5jY/Fj2BoMlNGEBfRUL2ZeaGytiR0X5ycs
dTc9we6DuGlzKdswpPrGbCV41bO9TGEcry36fXy+VcxvLepf+DJhaF3P7jRgHsOkx8I/FYvG8f06
aLFSyHZqCHPOziLkohjNeHZxHlIw20bXt0snAQGcwZYtU2YpuMvmXh1Sd86ScZRB+QjJTZpo8079
wKqSLutZnYYU7wKlwkelZ1PC3wvAHQN9YAPka3vS/bGlBTmxQIAZ6BZCiyeXtSApmY3ci8OFyVo7
2ZhKXKoWLbMBeqromGZPRK/pCshb51fkY+BTg8pkxL0/BJiD/8Oq+f0WZkhw4bKiqkLqhBHDuSeW
I6vX++ZmYTG62JChZRJ7MaVvuSDfFomQ97YwNlkg2//3Yi0Xtupkc8Q3NlCq/xNE88Q4wUuoqCcg
Wo/TFHzg/w7xA1RWRHmoVXPZpXtXLYsgz6vllBHYdTFYVKr65oUBL8bUchN4yCN4H8v2/a1tY+U8
VCKoC4C+XMWr0RaJ8ID3zOaQy3dkL2Ae8U0rQS5ZSlS3zVGzyin6FMWtudrCrHfCDk1a2wrHBUn1
mh4wdd+lWsj710a1O72Z/QckvHR91aSZqy0T19yDEIP9e6QED5Uvf63yDRATZUtu3BPyZZuTog5A
VnVISKXT61/rY10jOyWC0ryHSfOdTmNEEEN2V74CwFGMSv2KaiqyBDI3QJErYLjdasmvDBwVDhrI
9MmPAKoOwZX/7Bv7TRpP2Pe1+ZwfvOYYc2FCC9vSe5meGgaq+uIfkkF55nHFMzgy+0xECkDEgXix
vZIHziTVpTHNyXbR3UvqhcXEyfKoRVvRTDAENFyfJsK3GZKtAZi79Y/G+V4hx5tZzOY7HpKZJYy2
wNVvpvAA/C/VvWWdQ5YRDrGMVkq81KVzxuJD87DA9q+wDkCyb25ROECfQ6tVQU3CwHP9XDh2xp8j
aMkFsnr65wt0uvi5cFWF11ZWxC+YaL0jydKquYtQffU8zXGNdXDvWoU/uuyFCy9EWImiskN9D5u3
C3HhWn7mvqmnN0P+x2OVmRxqNnV8Upbz0tX6amKoEes/wPx8xWX5Dt86lbzK8lxAK1LIGVturTUr
WDyK8nLcl+TFyQBBtQmTzWOAH+omEhd+KL3chPo+EQew43gB0czRSFmd0odP5YvCWFJheFzyGJVg
jZ3sixW1eREQLUq2mckb4VlfYYgvCFcXTh7db5XjZuhpI1BNWoauD0zVJpC4t5iNnL2COPVoZaAy
8s9uYaretaSqS3bTRK55jg5VDNg1G1jSsbcA7fLXQKKwu1QTLSiZ2aPX+iIARME/RAgYPOD8bOYU
ibmcxuVuCyoTMfK2MA4mqxB/+O/DcgTtf+3/ajtCq8c5VKJmfoF3YPJFs9GOcbCbvZHAWbWa9Ng7
XVxvrWyYw05xKMl71agRjNP+tFfQZVkFnIupVoeBMv38kThZF11HO4OTTCi3G7+UuFlUXRzJLtw3
TWrtPwWpuj8n2aTrCUPWYBf9sod0aIn27EArVCU+UWv5Qvc4KkWt/INPRlGGOU5pL7x/efw+qTKZ
dfKdx8bFl3rSel3vpJ7m40Edl0SqjFhQoOa753SA4cQ9vXDYzTrgfGoODAIRlEooBzDNgjld4jzI
67ctxb9qFt7/EtZaHs7RgXiD4LiQL6A9BnLGJYOwGI4vmP1s6It4e5rWwCRKhxC8pV0W8ADv9dlX
ElcEZYu+RDYoucHHS1X6cjFePBzD90UL7pzN3C1WHYyntggnm/5gU4EB74Wt/6rBpRGLYqhXx5c/
kVxHQ7I8/4PXeFdirLmi5i1JZO8ZYloiNWzM9p7Ihkuh4pMjsX1kq5yH+jqf0u22hO2MRnQaOdNj
01+5/L9nmllLucNLeYlfAxPgOj4NwvUcWg7Ud4w+z13EPflw5fFz2LIRFV6BO+0D5DqU3SiXVw/1
J4OZZcQWzHbEBFjt+lJJeQBWCMhbTzWSwskDOyeCXXbN1ZneVQqvPJN3o8fJJz+MRa1tq4gOLmLW
7FSz+s8d76oNqdjsEDH7FPFUh1VWQjc14LssyoQyenYETyZoNZEsA+6QgYPDYUjbOKanFNQEhCKV
u7INQkDxn9mmS2sqQjUxcD43yj6yW3XJy7qeGmIoT60Isa4pZT3xlKdN2iWgcHQkOlVnrG7/plau
j+Ui8o5yRYK3SpDe/LUvOwe9I58GQE1xRV26cRGA7a2ZpWzMMpM3+N1xMPXero65AHfpfES7x4Th
Yj13m2owqJDsWfcJZoiQP1USpAC7Bmlce7bjgjrlvjoZxwRv5x1OMY4iZXbt0LERoNu/EjGJy+3H
ayLY2w8vZXnd2g2OqO8WGQ4y2bGeSQIWkK2Dm7j1NGB0LEEWNa11KCEnjeXqja2E1fbBs4Kx+C70
3GdPoyYca0IheEJiBuTE7z86Q8V05aMjoIHpRZY/bB+TG4tCHFkTPWgSNMWJb6RPwrCZ4t1MMt4d
Vqm34jFkuHGkq5xGGZOuvVsnt4PRKxsm3jDNDtGBcd0ABECOXi6al+q2z3Wb9o6pfALi4pai18f0
HJjZPRPPnybdwuJEOGm+OWHE3/+T1KHsd5ZqPAbNltWnhgQlaPKxS+PRcFanHwMjmLoknnXlQdC0
9QtUewURkmaZXcq/k13nTDrxEkzg9uji7U8/zj3aD0f/lUZZamKa8mPTebi5ioMfVmLWyUYxqNrE
AuZ8cYXoM6vyALDFM9Iv42sNMIZ5QmFpXt5SDYFV4l3pi65v3+IuvjFRDIbVMSlDeLEQUKiaJn7C
XBeMXgmhigAZZGcOiKzVpBQ6lcHdMMFirn0k8hdXbRyG2g3LV3M6Vgknf/CCYGfJu+CDnC0R+AlF
GPtp0pMQuF5yB6EQFUDxrDG0a6r0tmg1kicIoeY7QNriIiC4ukXO8/3w2g0vzT559wymfQKFQbNN
5rsnI0Fk9//VnptuVb3/zoOgzkVkfmar7teLWeL6O1c23QuL7RqbnfNspq7RnYOdFzcUTVmBlnX7
CWb8GpCjzB3Jp9OW5MsSYZu9vKUtmDfdVLSObsoODSsibxAJ3Nb+CdA6h/Xx3Wy/QHWaan3JHPjP
87sqqZTPJN5Omi69KUIW+vly2ozo82KGmB5IIzrN8qDYFdrG+87oM0EZzBV6EOLnjZ4WZzAFSQue
59jYiTJylVmrAaux/fA6vPA+L/TgIgcJlrZFWkSKQW8aYQ60AC0bgf1pPD3fWZZFJbFHUeDLygUv
2ztsnd7aOBAggL81Q/LDpxGtLVPa847dUQUvsKid8zVYPk+t++JDJHJ/gJIYecvcXbpj8FVznAit
KZzqLKt1BkFoMlmvo0BRzL5CUxuP5aWNsZ08BXX2g3V4052bpKabNz59q7c+ZB5vs/sEKoRBFT/7
wWGnJeRTpMVCPt7NaWDdvSZKVrHx6ODxbaNRqbQAJRIlWj+Id/OnB5iqKU8UrbG0RGyllL7U6pfg
bP35zQNcaMBXbGgCE2R2XiZNa/k6x+yvNTO64g2Rspy9SmwX/bSbhgT/zPqi3lGxr4ZLnREqoGre
DxcmufH25KnS/LTb7a1ybxbvlvu9WFyw/VATSeq0mYID1ptzspQHXbPmjGbbZ1NMQgyG1NlEgsSJ
IM9/ofX1dD3P/+ri9rkO87Re/Sr5R6hCGMXAFudGZaF2sJBWULOwcvTwuVbFoITm5L2H10/UEUzJ
NphCtUNcNuYals0kT96eebySk8AUx5sAoZxYDw1/GXUqTOLlDhXEQE6wcDGYwV6mhJ3WPXy/qV4x
yJKX+GYxzY2tPianB6O8ERTWBkpZhN+PAb2WaG/ne/wj6xOAWiIFLg9PAcQZIpQh5c/QcGKg7cWq
UVNzq7GNRZYfpEWqgVtX8c1m+dd5dhMCmQy0F0weowLH52LjHOyh8L2DHC4ADMVSRcwmeQEPFtBD
imNqGif7uP842lt4m2dHKdx4LVKTR8P1NAw9G8Ugs5JaITty695fqbJVqTI/FfTlKPim1RxVQf7B
tt5EKp4cqrb95/VQs6ZMfew9/qNl7f/qyehnmu+FdFQwoQIlK8FbN0m5OOUJnd4xvYoziHBgU1KF
hxlk4vTnIBNA0hz2JFebJACEtTTMAVXoLtrXj7Tbmo6mg6hL76OrJc1vYsQO5YiAYBIG+VR1cwG8
qV6Q6U1/nq4YTI7+BK7DAlSfSJItshgaPyOndhOXYi59s5QY1AiDUhAWlaurww6oEp14f2wrErgc
sgEkTjsBFzLEhG407Y15Vi2iDxz7D2+bVpaWSYVh1x0gkg6EkRRptfPr8gMKiUPyJEN8QRJ755HT
1/Th2LmsORgJjscKekSfeZpR0Lzh13zPVrGzgqgqgVThITQV7TgwQjjjcVk4L1TNRVwsMslMgI7N
Es6UC9eilGqUYH/wdwtH63MKFWBrvDUW9HazOe/7KECDp1Gugq6SQQbYfhoAg3Y3RU0zSBAWTmc0
YymXcTZTHeqONR13A/34r/EbCqr8KB+fiP83VgZNMR3lMGn7mdl7oDesatse+KLu2zmbnwjCZmSp
eh7nFPH0wVHD8YOURqS9q7uGMpILWa3I9quBvYZ9RegpxhxRw7RbscvdmJ8gubEKqxW6I5oJToni
QPuha/UPRhlyiYap+qNeu1qJCM1TnwUXCEg/HwpC7e8Hxm1HiW0U4qqNPdJwBh+ndBixW35KdGgX
Mf0onNBtACdPE49P3dIERYx7DcmLJepVlpLazowb9QIMS0wNMEUy7ax2Tl6xQlVnoQZCDxRkYFl8
zYEcFu2ndrCAH87WdtVBbSj2/Q4H591duvr96IOdEwJ+hzyDm8f8OeG9zSIPAU0wCH9h0U3yPlod
7hXaj71CW1RtSF0NrBaPuYoUglfxRtdEP6pB5lwQHsC9uFWUrmV2loMBJyNOZZXMXKT6QGMB50Av
z5Iy6jiwski2NTWQbNmweS2HXYuy69soPnLsuAFHOGaxQ6oYGBPmzrSUueg/H0dRuH6lVehkq8ri
tC+ZpLoKa8xXLlkLRpBjATDKmB1LhBoGBYmBJfmgHUitX/o+REx1vR4HSrofVoojBhGtscNg/5Ay
a9jRp+IKL4zpMdwhmbRrbxIUKAqebBug0pox0oUJKUAmTorBlR84jOT+U6vKdKhEz0AxtmNPPZO/
p1nxr7eXJP8IRJXhxV4eddcaoNg0F1d8psPdXp7edg45JlTH/HZKizmrRWEywEEglru6lShsEj9K
/sWz2BGoxiDqoQngVriusTsEFjwZs8gZzsuMmzwU+wiZQPM7uV3dN3DgisvAZIgeSkoBPPrIkYTE
KKj+P6ut13nww9feqoEVzzdaNFn5ElrZy9fzxbhp/N15R3mGylN1qRqQwO/8+/iAHaFQogjlQmd0
FjFKS5lNJq4VM5hZW3k0xweARVOtBlbtdiN2nQcwaWRri0lr68o4ARvkYVro3yFOzs0tHEiTP+0s
8h8JdiNPYAub9oRDFH/dtZhjLCBkwUQ62gGs6k7os5jsrIIgslwTfsAOpexW69rI4ScMReJ2QwUF
NAQulqFL1mv122NQixmIxuh3he8p3n4dEy2a1tlleBuNTNZX7AHysCYsWGLCfjk+F4FVmQCnWrD6
42rz4rlHmigVP0v9KZNjLukcZcIUU0gNE57rFl/pRwS06ImQgteGVXC4JaZM5e7Zt01GMBVobaQ0
oDt08kGH1AHUfv54tWDjaGEWylPQYDW1meb0peMCm1s7YEvgtg5FM2MLtTRrNHEP7E9ZEab+z21I
2G2E9ljjsg6Sm/X0lh/8kV7f4PdEWwelQU7zxY3aqKCiwJgC1hgBLuQPNzO0TkD5H6J7mAhrcoeQ
LzZc3kw3xaO+IzOXjiaytt057yrzuHxtNF5t3kvJGRJNfXEOGF5YBPHfaOSrGzGa14TVXVlnpnkq
9jT+8Oyoy4z+6K9BuR5ap5Q8tV4H1slFRFoD8zh+VBzXuP4jv6hDIHTaD5dVA0qRC0w+FrpXsXxo
CO6SgjZHveBABzLAjy/wLxc2L1HqcPuaooYIadPCPtaIuOPZQJ6lqkO5BtJq8pDlrHfaLwPTzjbj
Ae4sIsNc3DxHekX/QaY9Xe2BmM2JHvlMFk9/Yb66M/6ZDmTggGAn8jbx88jTHzLTxGjJl70q7eQc
97HmSceJMHDKXnspdssoLdOmVG7LfxfdNfJvtbRtK1Dg4JK0QnyjGDhy5Eo0Ako985qH6PQGFy/k
lcA6vzP9k66UTwkRMRRPqtBb26vtahlWFixZeSFAd2PUNP4Std++dErznxr6s8y8cax757usifIK
wI778oiWxAGX1uM3iuDIP7Cs/C+x6g05TADSGJWjvDMthbmGkbpPK0ClCZTqYR7E7QdTGDtNtJoe
IB/evwFDyPjpffsdQzIqS6h0PB6XivgjcjnDluEsniZcf/B8dbApf/apbCBE3P5qOD+1GNOc1oBz
YEiWuCZdP/ruFy4Qn98M5Zv2izWWEz5cCEUaX5SeVKng3f0MlcI4dKMMmWO7rvX4RPXxekQ396iP
c+SbjnQQ6Zdd3+gtS9uJVQlpbSsF9gwt1N5fcJD/Q9X6xsSxpC5WObkS6KPgVkVd57jczpFrp+w7
Lful7e4lOeLFAxO7rpkcJ/zLAxR7eHN9N7A/XgSzv47rMuH9HxZLl/2OEr+Kvvn5jZOWUnHXjXbg
9Kn7GWNGVaJeeVVJk38y2KCdvA8SNnRHGkwFs6mHMjFvOxt4CBWvvxCQDtotmmvtiIqdceeRjD2H
Yne7Ouhw+v7YAvQnqzAfzV0u5RXIYfnMdXox2a7MXwNuaSTti3Fre3DCe//qyzYyxTpIDyP6rAn7
Ml7weowoDtno/HOJbHUt83ONd+YNwX41tYxn1Say73ejWKvOoDarld2VXetepUhNk3mVrEgg41+z
egS9EPwx0sU7IigwuQFK3LoFQpkfL6UG1gsGjhgfIGyu0+05SNvxRGvlxr0bsCmhqLxlMzUAF8nF
bXIKOPRzvRYOqqTvcLQEeCD7TI7RehoLat/pTxUXjMitvilPunIYWrx0LNaKdytmGP+l7IZXgbAm
phh8OMSUI/envx5LM+iHM+RVhu+Ub+bZzu/WL6UIhAT4uCFybi3Wr0LHXbsEhDa2gHQgJEMab9+T
ZtYTS85UsyHiXPv078+Ik/q01E+fjgjjqqTlx7wdvu0zXElgcXbp0aIVJDb+RwzC/+olpt1BDBbN
ynVdEcVsHfFFf06fkvbliPLf0ZkefPnGo+F+9uzs4T8yxN4pvLcUFz6j3RZ8rXle3T+DyYgCuPs+
v9sLMl5eoeiRgMeDSCsgquxnSjsqHrqSA0YfjlM5sUy2uAxKImgQvkdvEjgmn8gY+lXLHpnF0Tqw
U+s1Hx0ydUZZtytlOdsKEUaAhWJoRwtnHkVJ1IHuVeIcx/RWCmW5tUT1tw0RueptGW997beGugVU
Ih63x65ebEmcx2dfpZyAJrDz8TozUc2XmhbazIjN6CzYNmQBkNCtW80AVX7PU/np47sJUiQxCYnj
EbkJYzJp8e7UvaEfKuj6DBXtyYaO71Wu19hnDyCzBBoZQmg+DQtNEIhrsAamIL8zAiMG0MdVC0qM
fdstVPckrKJoi+ycJiX9nSOoiGwoUfIw0W4wN5a4zBqPdgpTdTnTfqfPKCZZtZPP8pt9n9SBDSKq
mUHyO6kspPNpH3oSxDDIYV9bLJFErgUE6xItiotqbRpNp8Xw26ekJZ+TNNkMCp4T22rKp/Xs3NaJ
OqTjZOoCWsbaAVnHybzYCGpCqta/hd/AR9R1U2+J89bs2LuWGrB3po3aJIyW1hVeF1KQjzXyM8NB
PcZdddOgAmZxcaVW1Qlq9nPE+OkmCOxoxTJn35AiUFCxHcoFgPCgqSGKPT+J07Ccj5SbpX4XCpIg
5+0Z2Cs13oQEXntPymF/spP+PIHbFfzu43eqGXf25uLHfuhnJwqkeNfM7eHvgVtok4XdEDd1WcKS
L85glbNMKObFYBmy6Fnlz3gYGOzMZjsEOSczVCDLiBVwtRpnesR5l/wUYX+fa/NOsp3kbp80TKTY
Wl1OdFBy52wFjkvzbzVooBJaMtBw2LJy3Kwx/Hfe+zZx8AG99bs+9+lyI5/pr74qow73ntx5ox1L
PByaEGHpHXol2/H7mkv5c2ex3woLETvqUOCRMoxbsARDzaycnz2BlbSDynwaqwTjusNmpfQyS3UA
ePbg4fM7B0ChGZZRToSrDSH1mubKrGNZc+ADcIXn+X9s4NXqPIiZVTGSCWFC+tdN25RxTw7A3PuP
j/qFYt3gRoLXcSYDZN0FXer5k0MtUOLt+XgcL7AKSdESf6Iclv9QxdF47UqAQq+iM58kbg458QjV
1gUxvwSXB/K8N2b9mU7xO6XY8ttcqt9XMrJlWLCCRvdmY2vmM0I0f57lSc3jlLmhaM7w5+r0GRhz
SpnXipzpC5+JyErTWuiY0zodxls7KwNG/lBn5y/bdK6kVKpsXq4v45YrAo+b4lcDVk9g5ct3upFh
lUubvHVGo47KaejD8Eg5VEm/CSS+IT+XcCLlmW7lQqz851YroA5XH4oCO/W16fMtNX9+TwvFxGMt
z0YxDoKIjzIHTgpYoAJflIwECyCjAXBi2dFS68vVE9/98VlfPD01Pul3XM/Vr9EO2XLzT7BzGXZb
Zm51cC8EDS2Sv4ZNod4Uxb6YRw80R7HkA9sij4M/FEj+1mDQ51DW5szUV8e1wrxa3HeWM70lpgBM
Ucrg+jJxB2tuydBhC/RZsJbLRvXa7mgKwJzEJ8SPN4vrm3xtvmuGCLS4JRN5AToMBjJveeC712vJ
AelAq8voD9AJyYF83bpI3JbAanJ78RktUKSChem0gM3/1PBw+IPOWvCNIiQywQEf9MQFzJjbPOoe
9pzla0wo6F/eLyd+x49PamLtEd8ZnaJlh/DNF8Ewe9LiXorOCqkvsCCb7VeeDOlftBwf0ZviCty0
TCKEAlGMKfIpYlqmWfQQ2BmhLNxx7rJ9PfIMzZ+tQa7yUTTmbvXxA126Cb4E4bw9Ec17KtiVPgr2
C+Y+I+k3vPPrD9pWf8M1ijXBm2jcWz2BJlnrc9WIe71dzzOB+8UOobqy/K4yBEZMUIkefPkOgRm9
HyWMoClc/l/WK2e5TybXoM5EbuJOM8oO8Tq6iGUlJPbJdlxqUACPQu9qI2Ib4Lv5XGKk6ipKnisI
AJ9HuDI8h4STmEoNJo2YBODTtkK42f6hPNa5kSjz6rJ82p37ao44gFfvF+AMMwjatgWmj6GiI3G2
//49AoT1wknDJ9yjlpsMk6jPE0zGk7sc873GbUEpAzuvm9hVA3vp2nvmwlW1duA4WmohUNuct2Re
fLAtDfZsZEEmtgLKJx540mKAOos8v3P3Oc2lymHI9tuMjzFR/USSSkB00UfsM8Onn202bC3G1HNU
T8+cJnBFiDweLqhjyRLzG9YWk0vXHTDzRGeL9Mfii688zBhlEPmrMEmOWyBnLTnokH4kFajSO61G
DcPjokMxgES6rIq7OTzIf+nDjTjKiqALp0CL2+AITNuCy84qIIv+EzBpjocDOJkIGJS+YJecHi31
XckJ4QLCr61NModDtf7KhNSuv9qq9RvG5H6hKNmL0F4dYTsG8s9gB+pyFy73EmWJwOx8FpZLcWc0
oc/IioEaNMwrBOz/rKeuUoOhhTBvOHNBC2QHpxz2yRWibpgBJja/OGNLFOb7u/ujCp4nRMcJjUOW
J8MPFCCug8tKfG8jCeRRtcj8lwy7xyorbu03QJTIHxUe2U6spddh8mYNVFRoDtwmZ5yU/n3Fhulm
PZdyG4AePEJ9qOQUEf/x0hdI2VERWjNZbL/WIU7QzMob3EcSwYrOtUwca4BAzhgX46caNTVmatMW
NUDLME3sDoYGO1I0MG5oUg9E0UDfw7hWsgD6//od0Us/fnsEczhM/IhpUAqsGcTciWPrmAtAagQb
zhxztBlyiNckr9r9kM0gRqT/sC8BikggHaZm5MvQk3pQXM+iA8W1egCwsHWNc9GwU5Jre/ziC2x+
+Nn8rbGSX69CEEsfbLwFHrE260ai0I0pG9jE/XHBv7SX0Xpa9wSkstatmQg0BN5NAEXOhrrvRH8K
gEDT4kJ2k25t8B/610cIU/XjZE5TPx8jaOSZSWDUQ9CwF/Hsa8SLz6CwvliKGyqDao/g+jOGS8W+
linbeVg3g3b9WtKEnYzDnluRzyO6H1Y+IEb15YCdlh7W3ic6z15N8EhTIOdnEN5J7d4R8tATbftH
PGBvYA8tJNX+369oJzj58zDDbgWweZXSRFSKZuJ32wvRs59sdP6IRLOVP+hrKvHvtstP8XKyYe6/
sZy9i7dPuULyYbYBNFGrbxqFkaFkTW80gfnR5hOPacGp48RtnqNVsLSWzH4FajtkHCq39gNMwwV7
HZtlGlA4FRrhXbvDsGOSwrLEXsfSep6xdshv89v3d7UQxaIJ6gu1gi7mTudeILxm4XAwWmnfKZK4
03T8ZPOUZCgg2c6GqDKhRQAdOpW0vvb0UlXp3+sfvdgKmMo5w2Sb5FxyImj3y3SQTyrYjRGRfqMf
g3k2XwfJZf3sqN8CFkBXvFAP7pFTL4NxU8FJL/gekG2YSAiyNqv+iZOJ6uMnzjtViN9E4M3+jSfz
2J+9tqXpQM/7AW3RP5VrMxGpEzs0/0wuPsHujf6Nuui7l9wnfIaEkQHtxEH/fjSEMHaaqj3MHTZv
Sp53LHKP8dQ6LjFJ+OD7u4xksw4sXswq7GpmZeGj2MiFqiPDr0ARqwCK8X1MKKgesUWTq0A25sMi
6vckEt20AdikTo/SAbeiUfZlI1MbdBx3u8tYwUzHFKh0mcWfXWHm1W0hq/re9NEQsLTnr4mYrotv
gck2IFSnGyt1D/L8H5sI2vlELkmR4p9BnTdg/YhkV7W4Py0V7HOmk4u2XRqKOaOfWMguGbjv0Q3n
9wHkwtKjxEQWDDezPOeEcff5BZAE9EMtTLLYu/3XCkCTUOcQdIvY7UTJGwSXIdfmQmJG/Kv+I9zM
fuvzI/D+EFt8Ux33ntWuQbe6v20F4X8HMMI6KJzOgCND/5UM1aNMiwT/OE5ATZDasL6ZOfGf01YO
V8ygMrhYBK3VGGU2YUNrl1uZJljptTwUIed1pkSHxWWXP6Wtu6F51WXRYAqmJ6LvZrc/6A2OkVDI
t0NUcxidnkEc6VJQPfgpjw0Nz2b23EyzHYqqdTBNHlglNmzzauDCT579LyzGFMbqiyIAFmeZ9844
Tmzg5uMMgNirxID0ZX9Ihti6tG6tjk5ZS4EO46KjPQrNJMvPrGbdDFCcr0JcBHnnk5D0zTgFwYVG
xaxbRWSnXx8iQaxJBucmmfjqA7rG0A84fu9g8q5jQB8pqNNfM4I9q/vNkiK6eJGBLOsSsJ7qsXMg
+MthDblkCHtI/0MqWrYpIJapEHV5hBVPWdbhlbLNpXHOnNLjijsFkRvPsaVpT2tcYgU3dQPOP1hE
5KYHHVUXKWumephsQLVwzo8BmU7G1YPK1iCc62iZjOuiVOQx4IKq+lTHPbG/1CxKc/F2W3VzBRJo
w3J4TpqL6HuczmRdnWClITZcbNadI6XPpa3Z3WAFo8EhwMoVtPdlem43e6MdWG/ELSbaDVVOI22A
xmRGAu3UX8QHb3XPG+TLC/jpkQWXJoc3gxfGZ/yitOIZUJwXsPXNhffkU9Xv+C+IIbEJ5L3+tD4Z
sNVOpWPi7AWUhucb0hFHc9o2fWgMrY5MIcrxZh774dlciUvRYnBEe0K4sv93CeSxEgSd0hJp7v3o
H/OGMUwHetEMVjM5nI316O1OTwHd4DTqo25CagR7L1xqmCrC2dBVM/riTVSCfpHVm1pW9vkghGl8
d1WlVcWsVG/DAO04KeJlPqZQ56hIfEFOTD8jmJH0p3G3mFK9TSP3Hc52KBSOiYZ1K33pVmT7BbXf
e96y41gBd1QZSvIZI/JRMBlP83SIMY/xFLP3j1l4Qqxl5ccIo9Gcz0j926QEnlCH5Wlp1Kp0R2iK
IFDB5y5n0rv1BSxKdxZREbB9fwmXUbZIBWRtO4IRunOpFviHlN0nHSnN6qIjgx1aHAW0Ee9NYEkT
B8vlmdnshh2F2Wfc/xR70cFPTlvH5VgMwYTTJsXw4W9S8LK89hm2F5gU96y7rPsDIfAByGO8pKvt
EZ7rfviUbRf4Nl8hyv+mWvVDeLVHceq67WEUR5Cp7FQth7Efb8dgqxblVIt005FZ4VctOcduVP47
V5dXgvjT55+ZubVoTkw1TsJUVcPzWskC0kn/A8KP2Q7uu/S9YhFSqg85ESUddcjCruhN0W8X6yVe
AQviFUllt0wwDCTJoNnGo+XedTUwwWjIjWNZvqa7imIwjy4/RGmjXM2crB2MD+AmSiuhZEw8ZWmO
vfLPaWQD45SBQcBlj0ukIe+8UVvdeKggbXXo0PIUPnoeALL1d0V0k+wunjfAwKAIXgVr/ZSixJ9S
oAxj0i+duznSsVqbYPoJyIHoL94a88mYypJcO/zVb6cG8xbP6PGmgzwEB39zligl1NF0Unna0F2e
EpkZda3ipMYJiuvJREciDdxuxh+28/tT5irDvUcWpVpW6vikzcXDSWqbOr8w4Y73iEG0h1D+PLuJ
OBztWCf9WmHhHIWpyjLDUZyRS3FEIMm7W6aU+Peas2xmTjl0FfluKVSr/s4C0e84RPL4ubGpu+nT
iD8THfuHtwjZJD24vJkWxrv0OJKl7HmCdW7mf40IfymDGS3Ghghvw2CzwMWVwDl1UdrNd/Nfpo7E
Y+V96yvcYKHA+GI6eFxueF1FpbLwGEwhgdDKcCyhNcBLUXxm8aICgY8oJFF3XAxeOTnb3p2To2hq
71cISBNauZf8G+AVwqlffJy+VE8GPD9SownJpKh/gj2wah1BOpCn8k1lXoUdHj9jBERtigd0xh7U
4pIImMpMuM6z4l7bZqgFWPLlyO0zdhD+vr1VB9FrybQqfwxYaGrTPJVSXZQrpoq+MHADdauVewnw
yypwx+jBptuThVXe03vZ2awIBcGpPbR5ijc/vkSEASFwUJC9eREI2IXddmgPq79Iql9gvGfvdo5M
H4agSjPEGhEUeBxwdbS47ZJTtn8Fp9qeHTlvlA4TB28CNg7sybtYBbMtmveYEQP/vOj+t8oxtUT2
8UE2CJqvHclWx5u8csxisr/oXGKKVwVBEFXOEIoiHla0/fRYhhg6Xzq3hKXNYwZeoBHQoUhZcfQM
2L0SKDtPT53LoYbE/pr69jOrgxi+0S9I4dmmpLiOllDX4uk+0maYf6m3Jq0LqdGUJe3FYHHK9Y4D
Q+B3JmdZnc6Xk3z3FVkoPG1HlI4rxRixZ/ErIx4O37Ahltp/HGLHWl8EI0FD9cr+J53HycRTNQML
v+WJSI1/XluK5GcqB/rmuEPPBdatL1VObAJmLUp9uEUrcSKIVI/8KUnhRnHN0nNbVIx6gfPSTRuA
zNQ4IEhB4uU08ZE1n1mOAk9qYeMUo9uw7Q7TvGPpo87A+egbSj2po2vutzab9/KImA+lE0AHOfGR
Poe7NaA9dNGc76oVVpzzWipIDDPPwrw+nwcvHKcUXDyonqyyfEqhSMTjzlt6R2Ze9dcVeKI46eMA
g+XxoQ6K60PdhmhDZQd9SG/f7lenLWUR0Z1EN4NMKHaPNbBJFZ6IKCPUblFUinBvXRyrLnhbDrjV
dI/VSoAYo0ce1WxLwzNiPAxKpgsNNL/7Moq7MNrm1RvIVu3lgXZvPzwxQirFHRkYJT409sKjul9H
rZYoU+FX7TIgvqwFHwBJi0BYzJmDbPR3Y3zynZwLje6uzPA3Rh7hn0XGxF+0RZNSnFRl3FLfDAf8
dazu8iv51wJEbre09efeOedLrhgNvsdBM1jlzX6MDN2/x1r0Hv2jjcYv5hx70RXCWknGZz1kG5Af
lxdIzfwdJTfw18ZY7UN8S/84bVW7YUdUQgRuzHRltKQINZo8HMK2uSWI5ILV4ED1j4emvs5sKQDt
SzJEp+CBR3G1NuHcvx20tTOz4Ax8+i3ZMzngqECwtqthKlysNgygkg6vq2BE8ZT2Wisbqi6BBQnz
jaj47roA/dpjBWizk096q17RQIwI1OeWaBWjoRl2LcEs0uG0i+ZJlzkUVaJGHavPefyNdOAMDLfe
deKPXrvcwBf6tMvYKVQ6ea7X6xsvy31X+zUSGhGTgXzyfLFzRPf9hUQLAjTXmrurFYBpy2d9icw4
7WMeMz91F0WsKS+wQfGvSc2XRCBAiyConM1Yk+Ll8PP80dqDwoiwFIY4MNPT+Kwremb9Yg97hmnj
foe1ufotgOMrISxEOR5XTTP/rd9trIMBZJcL5nyJzdVgkdmLkSRD/eyBuEFK1dzgsPruHRlZ1vvd
Poc0p3yWMITZXd7cTadFMWLUhrdpAF0QYCBds7DKIBoei26/r+cqmLINpArK96DR5nUyNQMtSzon
zNrXtp2gFgHhYJbTi3a/eYD4aiZAUPpDZDSvcwS/NTPhkUPJaX1HsEYbyov+f1Oa+gJDhXbJ95RF
bXgLdFP57y6lsZhAneTVWQg/dKueOIh8WV58Z9ufVujfs0lmwX7Wout0fjuzsX7uSaw0CTfJDuzW
0J6hiB8edH80ZfcSL/LFHHR9gRlxpzOy5ccng0Dyv2h9SbllxhuR/HVai3U5u7dweXXJ1av0wGfr
jXhlRz69y1pZkO6krecPvnEUESIPU6yrhY09RMo2GZYdzeFKBl7s+zubxfoGJDA/AgD1wIV8Myyh
lahR/Dmsq5lWFfzDEfjECiigzFM5QrY353X95GVHUToyBtL0zbsit6Kqs5Cag672gGSWBWpXRlrN
hWqVClb2T1rGfTKGFRk5Yp7hHAttUyPZK+LOr4sDxO4NOtQU/WPze6NuSxSXSYU0MTfv+pGxSgck
B3OSCU9XxVR3VWoLNPiL2UYU+5IxcFltss8+ecWbhCmS0H82IGjCXcB1bQjOOkvB4ROVPvYRPBSR
qFPKr2GgvyYSF8gdpYycQ3i5mdlCjmXZwq1FO0lWjkbyVqd3AGw3w1WrxEkRjOhRgWQP8SW9VBI6
VYotvY3kg6hesRmi/vN0b5e86+23T5/HcoD5Cnp37Hp390eg1E2illUkcjLAI9Q+06YulnNQ0gBb
a3kJn5NEKm/2CfEbyLn4kvbGainHP84jXecWqpaoED46VYFf+of0Z9K4QhMc+4YA/6i3coDZmTxH
+n+rMGiSaCbrY6VDqYGgBpIZ2xdIuUbyjkHSmKVOF3wIdv16d+JjhkcYq96+Vq4v9y/bhJ54EaR3
kjhtdjebucTeyEhBwdKfi/bsY+swU2pEPuECwpk8sE8ZnnQancl1qLo//luNbxP+amUIDzmSLkYW
cJhdqT/u+mWAMPlQ0ZUVJ6sKU8P9jqPRehosBlV1AxeMKKGBGkjXltkDqTWdM5PwWzggsroPtiHR
UVth95X93NN4fL9vKfFlTE1JlGmwojA2KkJPgh97enfH68xRKKiSERFgj41wVTMvdKanVv5UaweY
pFO1qF8ZVQzc4KOfyHB5avIANZL2cfVJ+uvJJmNmHg5PGG6f8T5kEKEPE7JwLEMgwnxbMIKH8MB0
FA8pPhcP9ZUnJTPgrI4GWDpCjaeNeC7hkQMbnDwcsvtkXOllX4pdXMy/KnUEy0zGrQM/zOVJSX+i
J9owW78100Epn4fb21czO6aquC+1NyE35CmT7mg3IHdh1KIu0gdoreD0rX67NIDWpSu+U+hIlzDH
t4CDbw9kzqjReplcBIffIgBU02foeu9L+FvFUecJlCZeIZyzPgDrP00pxjHpjL5GjCHwSohJItAd
7P++kVMG4HL1wt+mqibPH9iAevM9HKL3cp0kpv4jjtj3ecJ9iG+dq3LUeWlZ+xBSNAFxQ4/mJhpo
lC4yNJKxjkEGnhrGBXU3l8lD6DgEqc+klC06bdpCdNlvMDO5ca5tikFtxkBL0fMkRlRDrIUtIOy1
tHp/Zf3F25oj37noPr/pQArezVucv7lPi2VbwRhVi6ufykLyZWsmQt0t0oOhXvvRf7pdOdGt7UCn
M5EJEjXcPUWOUp0ML40W43TCDSi4dftr3JmvKnA3OsJWvkt5tS6EloMu0MAqW3I8hMUi03KqaUDM
Z3N8IyjP5C3ZE99oPST967MR3hmhNKOuxZoatzSQLIJm8FyC1JmywyiWVxytme6U7vLffmq1mfkU
OAfMBYn3wgPsVChBlzcNdbchk49XnHuyIyeW7kG16Ihd27TJq8Xer7oq9U9CHOBzHflVINxNom7I
JEWxfu9DmY6hUNHROhVg+qm1tSaj+JzjkhAzWe8j3WpwaAeqIe2pR0tg54jh8tG6ODy9m4UpxRyI
5Pk/Pezp7Xag42SWzaXZBTfRQ2XVleKAXTbLFzPWMRpQ4MPDPsdlH3Ryc7ygjSMGTdFibwJpWP9V
GrILLqg9tc8tzTcsnqJs/+wpgXXihJZ5viIe03PU35RWsK/l/kAfoiUqXp+4wXmzkOXfiTpac3tz
aXY/diPKm4WRLjG3Yt8K8IDORt9RYbfVf4G0LXm1IKmouIeZbD5BnS2eBF9nIfDvJ6CfCFUAazFJ
f/IXd5SSpY+7p6muYbZgQxPjkYhVZ8LJqoTbXUwmesKGIbBnYH/qCeSiTR51cQ7SmtvBvkCZ9+NQ
n+VOaxAkajJI/hq55/i2qa3oxOYOjpSJJExbq/+nrC4gN8LKt3VwbESXxQK45nEGN/tSNn6B8FXj
s9xgvbw/o0gUtcJAdy8Qhcwv9kvyvBX2J+8Eix4J7fi26ixItBRxLjM0ub1iB5DD5ap0ap8C0fsN
tBX1A0tG/5zYUGAji74x9h7QBq145hDiXy2qwk7YFjYTmuPcyYfCs5D2TCQaQad3cU7qq9jI8ehy
nXWVDfWWNZ3EOPUe5UE8/S9AKWorYdVrHp61Wn9gL86YJCUSs/aEYcvdigV86LXvkELlU7C/OBJi
twHBElT+FAPlnbS2RCeJs6lpyFtV5+lyKJa7q2kz+sTdLQ9brXFKOo2pH62bIfNlkOgKwwVgRM+z
8EIRd/mRbUAgxw6sNCSQyWOEOB/FzEeMjXdQoThZdIqeOPFGmsfeV6tQtj5KbzyRY0oulYm4DCMJ
gCrkMXN92YJh+W84yPYGtE5zW7gMWQl9Lh0ovF6iP8/KS82N+D6PuogAm5cSUoS+MicckJAdTYC2
jbAzNoXuDcgPbpj3PzPO3dON3TRBMOgP5BbLm3he3qJPCnquqqD4n9uTvWhmXXjyI4U0xTWVbuXt
OnSVrk0yJZk/OlDeCASwzHf+k43iAGXOoZ0vTVc29Ij7NiDUtheAltvPFXlUHJx8JRz5uRxMHRzh
zu7kh+20OgQpCNqmP1p8ZprhHkNlwSFvVVaMBQ1wvfrUhnsL+yteM4lLRKbQmh0cS47OahAWo9Bo
Q7YO0LdJCnoMV+I4qTWWxrGC7vy2hvHbpB6Y2lDeu9VJl05dJw4hw3x55Wj0EsDVQetcnnR7dREQ
EbU+KNKjtgDtVblTXj22msZJX0VbJ6IEGXBG2e8HJJoFAOl8DCCWyTpbqUJFhH4lf0kgG9GH2c5g
iw6Wc0G2+n0A5C5UTWbPCQ7YjjOYN7tHjByfp1LpxJZhw0yRTfeVdbOWRO2Kl342+GkTY7/rAaO5
DgqrfVc7p6IkiRd2CW7pfa6LvrRQ9a4B58+xPbQDcXGdRsDXvK0pK8ki2pXFgKZhPMC4D9dqcYSp
nC+F+MiQK8sx9atOCgNKYmzlCVFsLLi0WCFe7k13SJ0IoVAWxixaO5z+QudIft5GWYr7rshYmF3o
EdmO/v4BW3plMAmy8/1z58bBL2qvhZt0rDV4wGkFQSfNwbQgdnN9LRcqg8WOOTWwXSNzSQALDAqT
0/duB+xiEpwWlitM0ZXkrxIcfuMwx72zrSZx+UTqPxgo0nf5J518K1GwxNj/66kt8APDRj403lmY
meJvbBiDPnLSafeta/1xq41KbZ5cn1b0qqiT+onSPWjWW1oFpIHlzeEh629ujN1+Q4IWOaNfnL+M
OpchFoZO8IvtpdaGCZRhJz2I0hqlybJni+iU/2M835KaDWBdghobnGNXrpCQSW76wy6PNVaJJc0/
0DVk0C4WypVUv+P2uIuO8gePROzcFM+j28c7z3MCGrND97P6/0vFVL20aKe2ALH33Cw9ebWEjpqz
3jFd83z2JCgV78c6SKo6j2gF/e4741TVgMWaVRFMkbmZi6vLCEN6lipqNjteAyLsYPEQqlk6IMyn
0g3LOpOmjM5TNBX5hFakE7Ey4CJCSOs7rt+iTVb53pm0HAMwcijwEgFyTWxEmLGH8Lav9ms+dgrH
rVOvJ81zW094OY08zRSIhKwAn+qomKNrdfb0dwjikLbacROUvfQAk4VoH/YHz5OuR4HGY8NX/Smc
8iCtRdmjxuUz+YL18k7CIKvRkcH26+0Sroje+oyk3V0RvSXjKUC9inlZgsLYt9k6szxi7IJDke3j
DdZ/UnOycrl2T72TIcoxawHfPkP8BDl1ILrsiyypkhXjjw9xwZ4MpCF+zeKZZjhhneqUnrPXxV2p
Xs50yNQf3DIH1EJKLUHfg92i+odMnhpJYQoPHUIkBF8qXhWiOBA1FnKjdgPgFYzkxImckxQT5U4z
QxohaombyaopovjNn/uCKn9iY6PywmvZTFM9L+lxpKE/dUwHqElMn5pu0HnmtPr0scl14s+ZgArj
DweKXId/Rw99+CnTpfFgMoPYIfMQ+Ql2UM/FtlmLQ/E1bVwu8rhHpMdGQkCzJGR2J2DonyB634xb
9+uQ1myc/1oY+saoXcviauViYpZ8nEdeN8ESkad64YosHJAY+g2dELfS7rQEq8fycjzyh6aA0yK0
LvMXpPyVAiT/t1tmes2cHhTwq1F1klzqeVlOCtuUBAdxEA77yuxqp1NkWTnZGVF9UL/WoBFMXDLM
Xeu2kiGSDb/E3VR93ERaoyjV+75qGFFiMovM93PSt1IlASmdUXIYxBorcMmgWP3JLynSHMFuEzDy
ohkdYIU8TP4442Ely13sH56o2xVfa8eMEeIN1XgyCQWR8RwkdVIavsPtqAS4odTf/ChZiGCY+vA1
NwmXtBTmL/U5FzaQdwsbS912dx7zz0lC6kTPAmA5SDk8ws6vP4Kqsw56vUs1mmxoodnsCeTk/Lqt
XV0vfDnlP/gPmqQz2V7vADzgGPbO7FShdaUP57znIUGPV1p+BEAEYeR5MTdVRykkY8LRea/KqtPb
/jFdej3i0nnFXs1ZFajzUOkeysdC7PW/0GOmygQKls+O6+P3DhaWIgR7Ia2MsrVpy/rrlD00v+Pg
+i8pQrXuFnDuU29i+xfxC3VuUfvop5XoY6j0EpB57MDwnyB8jPV+RqT0bhqb8PIoNkqIJFlMV2Fx
pxeOpCiDeOgWmytkxr2YEfiPovwHxHfEKcOUm4zfYZWAMFYXZ1EEefkdy4sl7moV/3BvD0a+QEAD
lMc4EUuSdIHymtP8u8l2ohUvYwW0aPmU0bix1a/mLfs8Jzx6Xi1t1mdxlCni5BMr4ZACqm4il09W
IOAOLnZjPRu3u9qV954tOwtTU27PD+DwCdZ/aQKX8CjNL1H0zz5i7idIx+q8rqTMTUd6cfoxwbN9
EbXjgbassoIr6erFF+8YRq0SfXav/ZcZ27b/Bc0iZtjEm2h05HxPRB1EymSOGR1juJJ9iWWovFRt
E5RWqLiIm4xSX5CZQ04O1b674TpKBbJwYILLMZau0T3su+9CnxCaQRJ4jrGB4bIGKaspnqTr30kp
Q1iZ1Qep81ItKhQBmO6dcXRC1YsRrTOgavjF6AJpDQZL4HrhOjVQCoj0w5YzRPH5SkFnow+UJpVg
SUxsebpfHsqiAbr5Og3lETDad7zYGutaB6UHyGAsyYawOIn2HNwmgfBTguZlNV6Rq2NPU2lfjYe+
1B14HKiGPHO4uQv8OVwSvBNoxJ2XOLcQo5GnAPhmGhtsryYUbKQtxy5dYFj25arynUZk6e76LuZU
NM5BOC6YlBTtqT2MYMsGGAMX3uj1MEW/s/kxay7Li0/x2VlSroqcmZTtQdaK+76n5z3P2lZKtea4
QIVxH/wfq5IzmRee28dYyinw7wM0/3QyYVdWPEhI08xx4ubAV76p6Hq2fvmjIUP9RBleVa8mF7Ks
1f4gCHQ9RfnWjCbEagbPBJr9jK3BiVMxngTiTKdzb3cgS9kppvuumTDfoh7gYxE5v72fHb767zg3
k+3iD6YDgB6BbrI8C3b8GST26bdmvN26Mpm54G3zSEcqimPzSNzVUHRLskoCbs/xlG27WuWpW/GI
mXtfXNoI8IB8SFL0ThyhnK6Jyfe+evPrIRZ2XXcJRIT8gb9wxeAmAGigXuYPTw4YwE7okA+jzyGa
wLMp/mXLL4pL2SR7U0fH+jBxOn1qcEHju4sCUW+eyi0QbLcjRzmdYG5PEV/bQloZm+O0HV1wx8Ia
hmNntqqLuGtkuWWvEjVRyP7+BqTWEA/UptIiLePylOsHIyDAcF50MQSlwDCIq11NO5uG5YEhV5Hm
tTakontHoLj62s2krMlWi9snY3z36pYBACN94Uti26r5eubOYyxKojW3vMg3SFMwoTzcGMsBFWQq
8s6z+1Xkcmuj0G5WHanMrmcm9fguFIgkBN3U46UbwQi5XHDB6XIOMwc0d5sRQWJzaTugbrg+ajK8
xgWUDGm5ujuZt7nSCrllO9nfRKtGYhuY1No/iRVQt52f0lM3ZDrzyJX0BIAaRV/yslYCKyOd4y9y
vWRjv+qO1TZKnj0Nb3ppSoyQgk1+nLRBli5F5oHapeGaqXOZC4fU/GZleSuFY3sT/xOCoOTHwgKf
g53FxIKdlNu9aNOkIcXJVgWE55WC80302OJ//A6TCIyRLm7D51VIM/DZltjT2Xfv+yyCbHd3Waal
XH99jktjog6WgZVPl9Lj+791UmifqcuEOsN1q1APzgbi7jusNJfVElYusAsKZdBm3cfm9M/K/7VW
45xX6ekg7oITtEThh2OgeyjAglnjboz4JhNw3G8axbe2zZmwxOdzpFl/VYu9ivetrrIsWPJuGKpB
FG4kSrdnROMOBC5v/D6KQ9FDiDprQ4nsZ6yBfW/w9jAvReSaBGZXmGNgY9MVLjbP01aIiNj98vrR
b+EqJSRtexf3UDoZRKd5F95d48txFflJaj9h8Sa7/6nq40TS0dayY6708CPEisBIgFGKw6CFHiUE
XCLm+1LdqxM8lCklF6YSY+3XATVtfT/DE8Jchtz5GLNThtH5o2K6UMOlJSfOOgD83sH7h9BaXUgZ
ljoRRZ+e3Jc9O0L3SK6uliHID3S+G/OFCp/GKsc91v+/mUOg1YAGTluiJ3E55D6ZqhKGCfNca1kI
YK5IyytKGZ1zRdNxfgE09ce13RyYGeiNmmpc/98qWFxVhJLl9rucRMpZnCI2N3mAraicv0BcvSip
fo6/rkJs6O67MvAlzeKkaDoaT1LL7XP6M2xlTToaF47tcXWv8Era5KjHRww1bY/zKmbMDONavchv
6Fs7KU1o1Gvqx3ajcodxY/uxO37eG15aNIZy+fEGnsiUqxviiWEzSJZNR0sNh13tXy9Fy1lB8jj8
7duo7tGKvXGShJbIdJmquHEA1OQJuxk8xhxIXbFq93xd002/BA9OgK+AyUcr0RM06b0YxVjPi91e
+9Z1UoMDzjNrydIZXQor8YpUFLQWGN8O+IC8NX7FqB1uq3BvK0/tHAuDmRgN7i2qoLURrAyhIrk5
RC/Ry/bOH5Pbumc8uH3L3miT30mLqsNJGflyBe/kytnEJI0u3pCRV4OjIhyy7qiZduaJweEMT0QV
tvJzmh57uiL83FmJ6K+rJ+ktwapaOD2E6gcvSXQLV9Ra+cvr+GFTdfo38SzoSvpdzX1+OP62DIH9
J0y6LzqBxYD+35ivQkLam/zVAuGwrTIg8W6ZrlmvaNkZkWSI0wEg9QZii7EunsBNTCurD6gh9Si2
1Eat7PSgbuVSOD6cnyGwd7FbRL1+sNxACqBImlCKKGqWEo5l9bD8dYxmvvmxYRZwzw7LNp4EMAPO
FKs073RK94fY+tHkFM/thfXa0SOpvf1/A+uy2Dj7IYYkUUX08uMMj8+JrbxjNB7r8n7kgvOwMhpk
YbfSvge8R4BA4qRt6SNwsMb02G0zix3u1G5PNmkZsVyHQukJzsd2Dft+0WWfV9Dg/YqI5n1/DXSO
dtS4rNUc7c46V5hgnJQkle56fNyuWPtQDdSe8cMYEIc53iwqmWnz7dAr2yz/dYEK1LNT6btr/Gl5
AFO9lJ3uZWeZ26HPJsRI6gB/FSxh+j6rGDK6VfSmynJ5KJJPmLzKk9lb0m5sckO+eD4zot/1k8E+
U+vdQDYbPB6MarpE9QbUvMRW1+RyuX08sr7KbM+phZkgPD4710skoDISe9SrWKoEdSc38DI07NKG
2Rp75ka9FUpfBh9dsiLFzHxDWzXlqui8+rWnIUZ/DGrLDsuCfW3kOyu5F8aeaWIvV8EcT7pBnuRg
c6LeD77kmrJrGy/B/aNAMP8RGAEqYQzIOCo4Hyp63yYl5+0IPvGCMvIJ1yVsddHID2HWD15Ah9XZ
PT35v/OcchGSo2eYWuyasACBykwDm+p+MDXLOxRm/iD5kDBVRbzNG7MUlvbmgqIm+OHwUSikun3z
NcMwm4DBUAEow/YBPe7v+deGyFQ0n3D6eW4DZ+hfmHN2CfB05EDL9azzAn9NMywDnJzLEg+Ipdxm
sRsreMBxQ1tUaHXgPCP3nkPhyH5mtiyIRFk9mG8UBTyKaKXflRffe9QGYWhYs7HVENpjSwgafVTc
aqOlBOaUpF++h/nrgtaZbaQOmF0QqGwziSe8v4pYf83SHPhdcYfHMPzGiWexJzi2J4jS1bzB2jHV
T0RI8CxgD6/12+XLwTtI57ZEpcnMz5nM9p2blvwWpTemSgJvVrhbOi90gB5LjiXYhksUyPASgi3U
r8SqFtwlokuiUgOXGFGXvCc8uZeNzFtIh7087M7DkiqdL+95pQ7dhXoSPMH+HDo+3sDlJ89qhERA
xij0Lts/W/ypmGvmsVHbyaPMRjP5Hx1L7AhHIgup4YgDrWInrUEDbtNBHmnrBPQ0G8PzVENd92ez
u2IUvlcJkTJxZBU1aAGa0+Uj1hHhWsL6F4UMqZ1ouOYCRkDMyYZfIoOZ770v/Nx1r3jqe2fIV3v2
HuNpeH1VwpJU6ykRfcOpdXqdBgtzwmTdbQfqlpgI47/ItsAFqfEM1cik1eThd42x8g+5oRHO665c
onEdOEWjYZkoXKZSePju3B6quAKPE2jwFEKqdLcarts/uleUNeQ+PqrxS73n2RRZDjuYdt/3/T/S
pj8AmDeQPwE82ffP1AyIKW4sqqGsJCtYhg8kUOPLFlLB9GLs/fM3KUbG6RpbOuO/aDhOrSckzYSb
wDh3N09PPRWRGton7tF1OUWFdWj5oEgephNWlHSu3cWdVd6aDVD+xLWL4tlSAcFa5/b2qOt5Hsu/
tbZquJ1CHKqE3ZEvMyLxwC74ZFgcswieyAN0rWO6VztdrO93lc3i8K4YzBB2ffOf0wMEda/29O+u
v6ycUWUn1A0bPSNFjDp3xpcB6lYSQG/1+xlJPmEoxakXTSsr4Y7Varb0+6yH5TZZ7WHha0Smg5Vv
4rBKBDfqjWSOXNtg4nh0nIu9iV3n4v9jeB1BPcsSqHwByM85Yt5oC56dV6DkVdQmJAdWDU25NCnV
zhzHFbX/F17CKXGODwB3ivcG4HR/Ph9NU9Cdwre0YfTyfk/lQVty3xeniQk62FSm6xHVy+rmuF5G
ePf26VG74i8A9J5XFoZGKKNrdLWy+aR9kCAFgPHWJdiqknAb0E0zRWIzuwL5rrz2ptY0EMquh/L0
lXU9i+D5bnM25JxpA0EZhOHySATnRc3zAVySCHe3OS+2gxxiDXNjA1UDPDOyBNONnDAH5QHMeHuZ
HN9rjjC6+IKN0MXZ9R/A/BZaA1lqhF3hN2ecVh5tHlAo+TTn67T2kFFf1xDWlCh3jQessgLH/tne
X9gIjxm3Tx8DEZMLIZG1t6q/VXHb9HF+N/a6Jf29djCa++WTehT0zISSbHCSx1DPDCK98ode2JBl
llWWT8uyq8kCfawuOx5k+v8zmRHHuq6CIW7PM2IS+HO/P/vQ0qBtVJzWpY27yzYqgfEPR1XnEpI1
zEbu68n+bhp5DHcn481ixE4qjz7tcIROhJm0Dhk9pEuHTpoS1b7cSMU71HJy5DarbQ0MHHlC9kB/
HX9BlMbIs0f3BmzfgklbehFCawUJOz2POfjvWuq7p91vjABsx73wf92xE5e3ohy4n1+MJInmL07M
CO3xpZI6+seIa1bRVqmjJilAucAIsogQYmcKuLm2YAKmDBt8mQAjdGfzFDm9phubW2FQkHfTVL5Y
pNdi76fbafCdRVMolxkM8CziKLEScLBCxVxDgAXlAGkKsDR795++T/bZalrjYGKOhBZs6u/TDi7/
k78mDFRXMmmCXC72vvBacb2keK66cSpEzuNjhnEmDy7PjkvRXD/Ucn5tbVi2gNmXW+UDJUP3th9l
iEbhDDXjweoZxtJpUcBftgwkEAq4nyX9spb/LuMjfU/uCperiiD5C0Jp0L5XaczFMTIO9YIwtebl
VzpiOSNSNfIfYyZqcGiW39Ox+rqbLoCZvYItNR0IWHx2vVqt0uRtFOXvm8PPGKBEQ83OR+06dy54
aeHlpnmhWl9A7s13VP8STf/qdyB9NpOCs81Er0m7UbhoTlWGb8GoN0SfQpSJRcpnpHwDLcDMj4Y6
BZ6ec8eYiUIVUzJmbel1ivduhDbwreWrQDt1eg6+jTbzACm5RLsEOfxOXbbXYfTJlGWsbm9SSUko
oZ3TM6A/RraoD4fEdaXBW69dMMv5UBAOxYflgkt/scYS0LdaEOtoanssYjPwBLVOwJkvCYRDo3mK
wHN34JcibONq/1AGLfGR4MdcSOttrPl/5BF+eRuQo5x2BTJAO5Dq8vCbD91Ubojo8PFTflzdDjjQ
TSIL3qp1uJ8t0/nov4duFosP9MPDEc4xgTZXCW93ADr5mZJkQV1U3isDv0KsZxVtQxVxsrEXmcOx
F2kZ0jXK1C/1NQt4hY+KnamedsXRH2eyepvQGS9UcpCAs0E7+MVEh+96tuFxwONradrSu+4cahZ5
asmTFalOBDLlXAOCwcqYY4aIzqutZRUJjcL7/6Yc8u0DX/9IhZ1pU5aMrmc6eECYeFtChiafRLP3
kjIUJzUS27XycSRFmOQ4i73EFjjWZfhqroSwH0sGVBC8+mU+yQ2BP8vloSofY72Xok2jMqORz6PB
WpuUb9wpLXNmmQROdpmUGLgzixU7ErSwKfuBqL1ekqwRIKERi9thn98ryNCRq7b+ykl9H4ZQf8Bj
NXnJ21AVgllTF4DydzXOfHEhl70A5WHo3KVooE1pjeqOYQUPTQQPihN8tUdmTIspZ2JhyU81DSG9
gUOh52mFV39jaXSL+wvP6J5af8XVBrZTSt60ozrakOHPH+WlP6Jp2AT5bsbYA3bfllyRVEFXKZCK
U3/E00Jd6+floI9p5F2l98sUB/t3Or7ivAwg1ZSTYy8aWXLHWJL/4q78D0xPDzcBNcCaQHmaU8w2
XMWrHnGPQW/O+uYNT01zjV4/2JjXpmjGTBJNdGOaNvGgOBd0m9faSIppbESszrMzUmKRGHL4O6rx
fn1SV2VpqTFMOdbXD8XEpJVH17+rDSesSaVcuddkLFHM9f46pfVNpXBV0K1efXIiXyvjnU/pit8l
MXEuXXuMA4BGnG4p2XsH8hNgNF6PDX3M5RBSYYIHdLAKVaK2nUZEoiB87adzpCK9nUuo2kuPJYxe
0qaZhMxR4SlzE/0PVZnaUu21mhUpJeV75DgCrdwAPEq4Hi43tVN+Mq1gxWdt6jfiJZEVzBtd03JG
1seaxw8x4Ne5Suzkg31lZju9Qfl8ZeSp3o3jQa1QPWThbootaZHZl01Z1RtJaxoV9gLJWScMfji0
Fjp19k6AcRjcxh5P9ml5o7OIaLgPz5b6g4nCUURDBsM+sDEf2k2RRhsJetpLGEr5YbB9fx5drSkN
b+JvPmJWIYrBCwKsIUaphOeeSurrZCIy4U64p5cjBhUfZv73+IZWO+vuzfEQHFLRUJYWc7xTY8hW
DaU79uTHMjsQsogPVLVHCx2574vsmm+yLmxFUtovmQlb6Ex5v+5tY3w9d0MfMSVq6iwu4MIg8TFu
NwEvBe31URlC0E+RlMJTFB1WZRqZFEOCHMvvWMEgpf6PaGFTsdTNltMz7gEcNAVVEMs5xR5CRZRU
JCyPrQ/L6UlaJidKxJ0WANRGjpZMo3d6hTF2yfhjRJh6wKa8/kCwziOkkM/sm22UcZPFUbjbHGBt
ql5CSoOFH6HOo/yZeUUBBOlIwtLSxLBx+NrjnS/Xrtmf3pVYZrN9AzUOLCcz9lO65eQRpYALGmmD
5Gs4t5pNGeO5zcvz/gasDQT209bDbBvL0haD9WpfqkyrKJRLtBxseIuRXGCJyrpYc7fLU9LWyAeV
hXDlkXLfmnFzEXRwdWMpd8300dQN2LXAjiGe5A41PHo0ylr73K5lHy2cVQ+zoIQs89fRaAvtz5qz
3RVYyTeJoHtg+QtS2xhOCtHSsxV5LQgp0cr1upbXbn+CwPHCqPFKhV+duM7lctIaURgWcEC9+YIA
pGlMePtnT1LJZzXhMgVTv+P3AfZeOuCimwb1/U3QTXsuQeg61YakB+AtpmonwpIBn/+aQq85g2t0
aWcht8rRrYfcELMtj6/fOyOywOhJbKZgH6wC0OVXmtYSNyDssGQmvzZQlKtKmnf8WSSnKg5NrDSI
CgAS3YothuGa42fGJ9+FavrJFYLzimhvDm5FrgN2D5bOAOLF+cmnmyt3iRT/c2CQIXsXdZFp8j6m
umQ1ktJQ+WYurpv+7qQNO2zImIK71VLgv9hbQEE/+lst3T5IZ8BDHekIFlhyBMOFufqKVuF6Q+JS
CBjUzoz3UIbuFw7YOYUi2ZJ9DVdeCI43OJjCCu1Hqx19JqK1BqxIwfYugm51ZUAUrs2sq7t9V818
RNWePYWC++bL7o/LFk0wMbuszsy+jO9H+1PDccpbA0hn1O8VKYm6QfHGOW95hiwXAmYI4aUuJJht
UCtMnDCeGfVK755M+/tYp5aTckOKxtgt/CZCJNGAByFS8v2e2bI8S22WKjc5662Gbiij+0IguqQ1
3Me4jph+IVLPuJmjDIe1yng2iIcLs7T+UHBMuJxkJTjK0eKEnbxxUBU5KvDPNelbMe8eBTL8Nfw7
wcxFk5z+KWfQXvNfbK1c785CkUY6vZxPDxTFR0/4YK/Qcg8p49rUaMouvvKrR/cJ6qK3FxANgdJQ
2w8+mSbdS1Pz/UTaqtRkDgQ8vubtdtwyjmT10eE/XLT/WUu65jyurPegjtA6hrdCSI5Xu8mMJWPF
YsVScfrdfHAohxWzJ3mFrhHFUw58v6lZBDpc6zyP0xTJKnEtttjGuvq4phi2VilDScCQRDpR8P43
XtmutCylIDgwMcDHs/EDZer375481eD2rScxzc074i2OdWp7g+857npZ6v/ZuZRyCbdXlLLv6Jdz
gRkXNLVtVEUpEUYI1CfKRxk79cYtgQlBmdyaZGSkA1odNg6knJj0LKFl7cfboie2qSQqFeUM4hcK
3KH7dlVbRlIy4DLyw/4Ia4MGFQiLxtsn6BzBHBQNRLVE+XnYcmbpoSZHxYj20RcsYYAd1pGWIpxc
Jrp3BacbVmZANoW1C4aexkul+GoOLCYbDMIKGcUdf5ji5f03Qf0dK4QDCDFXQA70M+JU58+gMDrZ
6bRb+/cAnbIIZwt4vADsA+MFw33FIcANwXqrqnzlNmHVG47Rv/YY6wRxJMMpVFA7P3N4q0jhKhX+
hHOWPxz13Ns1nOkoytyP3YkxN/2tNhpXh7pXkmyI6IusieNAZn3UW2aCYvU+fHB9oDMLvDptodtU
mb9PX/EQi9YYa8baAf7uxSI5+3sup+72PUOVKD5QFp2ByVIiXzW9RbC0hZr+aZbTMh+T1CLWWPQ7
gcH3AcHeIgMY52rc+Rn8gkkUNBlUm3//P70kQ/ABN/0qqRb02RbqZOo31gyReTlt8oDaZ604C0n5
cOqoGP7itY+qp1qjz30SPcI82TtwzbpmWR+wDyh0hhykIV0XxMi+4Wbj9Amg4OieBB1WybB2zeyb
hvvAG9LNWG3ukNbqvCk7dtYbDwpu1O7tomTSTJyOfh0iueoOYWX843rI5Azz56wF9fLdr5oKuhbA
4jY9VOiKWXYJ0HIB3HRfgq6WNNZbnyuNqFlXgocPbaEpQ+BWDoLW4gawCmoeoavnJf4jq8nmIcRX
EILrKFfTA6xSV63+RD0FNTjgics8pgGOzu60rzYlP7G2k9SmHwh67XyPDMl5Ta2yLiXTiUfuWe4q
Wa0ztJRl6poiqCqgVLlNJjbVVc+SleNCwWuHejpmll2xo7K5DAw/iUNJzWXQaZ//sKvcplHgnm44
68bqlKqh3cicyCAyY17EHVEEUzTcRKKjSn7m69XLNpTDnalx1AnVbZlSiK145iL9viRi4YkDFrSY
ci0ZtSctryLuisxfyXytdb8C6mvQNst2+sMjinxDrn5C6aX90JpEZW89c+uEj+PiTm6h4D48VnIX
HDzwupK8ov7kuPoWLhPI4h0IpFZ0KiehJvrzSuJVT0ron7a++7zy8bztbvqXaEfwlMDmCfIiHhIV
OoCH30xfsK0o8kWPT2a3sD6Me0RFXZRRghSsvo6NMhDOompYqAxqaesxBxbD7u/P5zL8v5Mmr3OU
wkC/v21iW0Nfd/8/bOJR1yf3R6UP1I/9tcMqHLm5LaBLu5tSQ1gr1VksBS0GS3FCR+XnqS+gsvfQ
3qpxqzMrbv0VZlwE1Nr3xbjFK9aJk/KSCSIJsosU8clFqw/8x3S4II/Xa5mFQm42cdHU9cuLdTS1
IG8aZWZU3gFkKgNZdS9jm8ggP9wEDrz9tuErcRoEyuy6R0EsEfc0Syjk8eNDIbeChQInV6P62EzB
vtyh9qjbEjYaudA3DbxD68k9KR9BarpNHshAnytMOIMKxyTGONWDyT32MzgQIXYfcCypNvcV2mec
S2Y6ql59Tpyi+SfOkzFpejHddyNUgB7MOCXCPAIrcbtHZcebqtwbC6yCmAhJ/iKgYtM37sl7pe+u
0iaNuPH/0M2xNO0q0toLy3pnCUt4wNHWkAS0J9dbyY1FtPxZPztlKgUkj3hfRXWpLAZVMpe8zLrx
dJybn0oh6yXkck4PSXpN7kYe6gAgA0ra+2kq5a7/HazAt2UXM+K9KIe2/J2il+WCTY47ggs7zyvx
vPfvtCm9RGpRvN73UamLsFTOnuPjPmIr7S4M5fXEEa1s/3mXniJxqbSXB6XFyaVzjEJOZR3KTBqX
IIumF4NpWObjOCRd1boZGk2zqW8RET+VAtrDExk/i2FL6RGjR+ja/LPZoHTF/U1f4X8yVS7noqx7
HGjytUHjShUlGxHJ+PGGf6E6ArMsdsfHi/6hozK79wLYuYD/dLwUB9Qw+vgL0ughX2WwF/9Zn4UV
uycodXkQ6+S/BF4eOb7FJRoAXVYHnW/R/QgUx4eI53nei9WH9wR//8EfxTUl6j3yKKZRRDD9dcPn
r/Eit93SN5gU/zHA2QhOTqQ5biypTrNbfks7Sm07An4o9dPDVRh1ErrvcX+0nx+OtcS8QFp/AdGF
9O9sCsCY4pBwAglz7QgCkOHmT0amd7Jd6Dnnz5eRTFBqGO0dhdFat5tWbiRgzVAIwjCKXripuSEw
o84rE7OOIbF74nS+zrgXolkuJ2DDtq70VSMiVBTH1gtUpc9RWxW9AMh3mXws2bmurJsUh+QfjTw2
kb0gFzLgdNRyr87zUewu2Yu9PUBlbY6kMYGI0ky07wGnQlwnZADadqfTVdYE3yxThUtdFPl2RKEF
XwKraKuyO9VpLEOdPknOKcM5CIT2butCFy6H0r7ASXoyQqKk0j/5xKabKPXS/HSkPcGtCdWDjaII
CyZO+wScOXAEmKcXzoK3ckwPA+5KBqY09rygXQ8/yehgglDjYLNccOOBqkVnPYS6NfM7YFZPkjjI
JVrj1DE1L6Q8zQdUJDiWrbBpkNQG3RB2iwqGrYC5uP66S+A9XzJ65sdgN8prfjha1qi5tMHwNgrl
1TRhms5I1qUtCx0AAjTWeQBextEja7Haae/AvKOPg6zAHdKAvrcue82hIP3IHapHiRTiP+6qAfvN
efWPhs3QOP1m45C87IzMx7CFusGxs/oShfpjw9yLPrfAxYgji5N2xn4jXGYRajAKQwclfOiYIT7C
dgHRwXvibhhsVt0xhQIN0J8Enxi8HMEjGcit7RE+vXKOOUqjBTBbgJfF6On9X54Bo1uzm+1FBVRO
MObS9svaJbzb04TEPGvNL3OAc6Fn0QsIVlwudsn7FLqV+/ss+UJIBdmGkHYL1N0wBnoYzybg39qh
6epSPEnMtfdtXE9axtW25OY/oFEoxl1d67YBOXPIW4GtBgaTF4cBtexOnJSJDvSqvyAiNKHNN8so
pjgnk8esdBtFa+M28o2sR+1lD6iziFR9ETQ0kCe/nWTBFW7L0O0lek+5szh5rxJH7p9XaJ0EV7X9
qLgAny/8/HjPSXrLLkCJCyARZxgDAPiEYYbpeYnQnAlzdTaQLqItdValiCfhRLxUZZ5PIo6xE/m6
BvFvQ6FNEMwP74kCPqm8cTyuB1XGGjYZnmXe4K2xrZOg4HfPZ2NJItgbCQ0ZmhXni90ro2qjOch/
NB1QJJ1lO0gNmtXN6INdPLvaQqEZtIqzNuBG7kd82z5XRDBo6iNIx6vFvq33hJfPZlrtqOvyVcDm
4NRcwrr7THsI5bBlEK5nGCFEamyepdaCn1AmcgKVLjKLRgYNcjgdCrC0ENQ5FlNGIJsT1Nh/jD0M
S2oqfM/u6kdzTBjyqXkNAf2ykkHoml1snuZcnkV+PdiSD6XbRiqzcEsJnsAA2ns3LYDE/Q7rGbK0
9KxkiUohRNdR/lMGN5urDTi6wnH9CvwBLGFsFds6SfKubAEqkS2ws5vgebfM0kRLt3nQaCkBtxgT
y+LhiXqmPdjQmeM+RxfP+Jb4e0frYaLtOIJ1Y7bp5QXnZVJvzQcMYEEGIms3RliI6/8iArhpXdaO
ib/yq5ipz8ZTcF61hNqprO7B82LcrQOaXSIQ2Onkv3Xa/WKC3w95bms7loyJMW6iGXsBeP8IYzg5
j1wN9EgxQugyo3VPgjTS5tLywrvLUX0IsdMspUaSFVx5RF9kO+6PY0L55h+TzdYHVPMnM3niKHzV
lByOiUy4Zg8FqzyC10xwOB9pe7jiMqxbkTpJdeP4DtSXg4MejhxKqjGeFvX1GoMWR4J1xeaGBv74
Q4/Pc1yT5kdZyfoe8yCyJ/K4hLGYhmU0Z9NUP+yj7oqqErApuvra/S90P6RjBZ6XEFSFCAJAbKW1
6CosmgfGie41gIrXIODjcpiDzSYmF51BucwscWcodSgsriQwEZ3jxoyqvnYVWmPrMeBKL5QIQpcg
WI6V8UjWnO6dpC/+ksvl9mIvuJIfM88toIFBYlw9SDjP4mDFqr/5SlAiY6yd0pkYHDpToYhJhEpT
yqrmCyx/zWDpMmx7mF5myiiKhovILtzNruPNMKjjReSAzOoRETbOuojq2j0pMw+N30QUmjouZpDG
nLoFIh9304t6aZtN0H5Lt1fufkbKFYhs9PlV68AvsIRW6e10FK4qO9as+1IFuM6LI0WpjHRUMgGb
vK5zihIey7pqHge0knas/R0WfuQo2OXAN0zzliw005edfe/mXTsyF9fxzoZrRPyYzvDC1W+JKp07
kOAN3rdrl8UcZlNAf1hM4TLnwuEzoFEKJaBsGjzmECNT6MmfmnsdsVI8f0masUnTYhCV6nAHIILt
fG+HBp6GWg/4x5arHkXt6GTS0Y4h7b4u7zFBMDskbELCu/ugyAnGbO5hMPPAVAtlgvZjECDvg5YC
DfigLrO6sdmM/1rvSz0DzHkUjk4HFRfsYCc5uzOza0YHWAavRUsj0TMR6OqXRaUvGjI9dZMNyRgt
YbhxAY4EPsdDnBQTzLllPex4yt0M70tE5rA1UseHSp333GiL9/ZSY2IcNTUouBPRiyWO1MsTwn5g
O464acSOoSZCasiq2xdgN1XLAF/iem2EWwBGmPb49QeNCwShvO4Lir6VFdq9SLWCuF0szxF2//CI
lmlh0eCbboRw+ANjFxUx3KeIMYy08pSt/cnEJqT2yPsTAhsM/6JZ6TAxMFxgKQEWztOEP2TyfhxU
ej63EFgbPZZjlimEzBvwQLQD25GZOgz23nvU0R35oKPf5OLcl4mRayH5LKoXCaKYVf0gue+N9ScH
gACi/aYpGNIBQTA6XZYHqbwSMd60X6aNnqMPSXvJWk/eEjYF7mVm6tJYhiiBmjnXnje/XCFLQpxn
ZJH9O4c1cHJ8hKDnhWSGErO7GNsiG9QL2WmBRMTryKYS4xY/g60RlvVqjZsIwtQTMpR0uSEavuqo
LA9B73caf4IPjVUfaQ5F4WsJCczKa41zLEj69juwMef/XVZ79mwPRbUO+jf1RC9kqcBPegpOXp8X
Pd+c5y+yMyDM87uV24YNFBsDnIlsTsMy2sFsaanI30Ocn3cY/bi02WW7wyDEXq4XMC9+hDMbNwWm
SO2YG/I1rXoAxf6mrkT39rBWc3BcsnsEjhRb3wFWfZuX7EnjX7EIhjfuTbUH3iU9PzZsrgnPjcO0
Mx1iVkUAO3fRxxtZq9q4z/i8jdIfwCmCNreHwydFXdjsEFeoE3DTZ2x23QiDtLbTDJsSOlQM/4o3
Bclt7gost6deP4XNo5Od8RrVWMw3ZpEfgTEvg/73Bu04QN3Ihn3U6HqBF6Cro9CxGxXGtuMC+kIs
YLiHzEiNIDoW6QXsPrk3xqcwxQo5j3V/N90Cn0rP+gvw2A9BH/YuTsWc7sruM0rWMXG0zZRfQf+o
XRIXWHKlw2E6xPav47MC9UeZitkSpdAdjPDtg0JR9uXejVPGbRJMustW+IbOd+3/8qxxu3d4mrAX
zBFvufDmAqWw2re5Nl0TrCsUZ/s4c0AQ5MyzVMdQ0rTg8LrWodoqj2KJL+Rg+Ca+Ge/oAjwYUGPN
3Vki2U/39P9llVb4wpFPN7enEtr+Gy+QRjhqCM0bbOG6xyAoU7JzSTsZlhM/yFYYTLCEjegaOK3z
d1uoduCdidZbLRw2q2lR1G3gc3d5lXirjcs5jTPRihOoQysorP/OzZBDA7l0bs+s9MJWyZKZiM6y
tHQyK0rzw+e+l6UHl7yXnVhSpO1qLOZNdQHotnxtU8VYVSa/fAIpJ7sw3SNNxh+i9EGufsz90rt+
d9EVm6Jz4tOXUV+pg8my3uFc2V114+vciND54GCR9jiqGhkKTI+l2peOPm/7VfFGMd1Oq07lQ+gt
+D9EbZFQqkJACmnkIgWxY5uu36qSvS/tzZpBSZKatVsPfeyGU6ah+34tQ9CtKmXhGc9GjTGjjvGL
8ofCDChcyNvm50eiLZjP6SEDYg+gGu35A+TWqxhqdv6gZUqvtx+UXb/bYPiTEuLCyGpfb76uQmdZ
zbCjiS/y5Z/Fxy4NMxRzyCEiG9GuWP4YFN974Ti/vZOhgHrNb9NO0S04OYjdmX6aV3gCYHWsCDaE
d6v77v6kGU87wZLKNXog4nTWYMbsjoBOgVDxGBCi0lVL+jnmxevnCsYMWeuSftNRpFhARXsODbX+
MgbQmkA+et8XDPhHelSEeq+JloCT9ht9QDJKtXsfisH69FWKC4s4hKWpbh6tvzV2irsVNStnL74W
mtArS1p9uvvHoKr8lG8/eo+JdT82slGp6ryuQqDZON9iUwMdbRuyGqyjxk5WKCduroh4WFxkfnTT
qPFPjdRjJ0Ccn4AVyhMR5rUSplT2UQig5gvXCA3192WotYSKOJhtrIcpZoCnhHMpgPqmobpVex5d
vSw3wCG+3SbLCHbYyN3oA/3REGzu+5lZCnik5OSph7wqc2GE2i/lDOJb8h5RRUdQ4k3pjjSikHsD
SjJCEZWTbfkO8xgn28+Jai6dnJHSib0KLtbsQayo48A+exxEtB/qYhwhayL4ix15WgzKCCDT0Wlq
M8KCHf6YPZ/5CUI3V1YT45uqMbFoRLAlEBLbl6mI0XwtzwyTwxp3famVv6FD+nX6U91wN/lkblrq
szDx3i0PodyJlwcvXq82K2vtNX3pVN2TdWiMkRiFatLdJEsgAT5SLoCFIxaMYiOBAwRdtRnRMXoU
qVNO/ALyGGM7LeFHB01yZTJj+iTIMKmwiH17xnDlX3/1v6JGTC+wAyDTfxu7yAsciBdMgoauEw9w
h6gO54MwXlojDCJyzs9CbUl2S2sD2GQrucCDr3UhVwwEDUYxHXMEDygj2i3pG3yAf8T64ZctONC0
Mgy2vcsII0kgf8Kt++60nCU3yEH40/k60b4Z1IeQn6VqBuNPU6ciQaptsCDP0HcQNmrVa7o//jti
T5XvCqKyX0vaAXUKyCtz4rDN6b+s9eV3kE/QqTCXqW2sNe1a/s+Hcj0mPKE3v/NLcaBTKwvZj+Ft
A7VevGY+ukM1+XVZF1Cu4SyzHqDhzz83286mr1osU0rmMiiD5ICZuCnIKfiCSyV1DtI1EyqI1kEQ
GFcd0e+rN/T//mJvcFugp8fk+9xqXzWpgFVnteH4OaruEG04AdnFgJvX6NyFk/O+Ek5vUfFZmjL2
IsoQp+PVvvup6/l6awcm2Sw3xujuI2xcTzUFJJyrllGe6cdwCeNojDM2Sawv+mUSZ23pwrk8SY+D
b4Z5AJF+FLxBGyUIGugome1fTvb32z88eCKpEizJuBrszvuBu83ApQxTnqWuWNweSql+7Fe3xOSZ
vwDCFqTZqopVirY9dWFnjHLrfGRbNB0/BCrPekL1du2KXFBM/if9ys8STG8Nx2CX7kfm7XYKL+hV
V4FbQFNB4caObu9Bi1Nihcyn2GiWETC9tlUFlSQ2Pxdi/xFCQSd4FkJyIT9BhxdFIKgnDCUsqvBN
9pn9H5mwy5fhfdWGN8CJKcYBqugBNy1OrqjMRWPmTlu3Wgep+Ztg++QzkF3bxGDR5gN9o5St6AHP
FclwbYkLj7IiixyN+uiRIM1CyadhEsrGYVZa9gixfRNK9R8xjKyer94Q9vP3TxpUvw15p9HZjhSQ
g1ka3W+7CvA/YyllNFPT1RVPlik8dQZybiUaAn3Jbmd7NYZiTn0MCfhtmBCvHMxuFXALzBMTklrZ
/K6liNO7DIOoV365ugjHN+LQlKbNqUo2T4ubnzzGCFEZ/pCQGxeOXFgSVsDVtiZXRbjEurmXtvxX
g4xKQ6m4zY6KQ8VwTJTANi7+pz6lGkF0OH299jU0aKFLOEdKszWGCfjcTMV5tMtNawGj/4pVdKyA
0ovXk3D3JAl92KLysX7K1XH2q2vsGBZEW8zhdqgjJ5lpi3to9WXetzWDMY6WT0oxVpOVS893O1nZ
qnpPeL2Llu1rq44WmLk14CzstS8hvTuFBcUz2MYPhFFuHCfpJMg+RWtvoAanmHdetLdQkvy3cjMG
vFKax73n9M2iexkd5CQx+CiYMmHQwoqIv1+8eDu96S0kFf/SIYubOVuswmspV3Hni2Ew0OZmp82n
I9DhIVHRbW4Cz7qmT1n16p9P5ELhSnIdLH3ExBfDwYkLz0f2VKBAPnjWPhFxRJRYjyMAo/qW4rYl
tDCe4xmKIZUpAGcdogStRNn1aoXMRFJDGpHrWw+/dU7qGGuZ8uS9MRayLaT6ElzYxQnwGeItKs2N
wX1DAP0HFiyjWUyZxv9iWpOXLrisL7FX+FHHsK15adm3LWIBtTQPykV6ihrOZSzKgOYPANsV5WNA
KylCtEBcppDQcPxsf0zdpnddTEcXzN5VS1jHVnMwu7i3KfYKvMNL0qIlw37BJP7jDRwSSKd5Kc3c
RFEwDo0DB1hthSrohttGvBqXSXxaLlydSQcSaMhP/TTsxipj1awN310myDopZc1Rw7B6uorfByY1
BnKPUkgQlRCqdD5IByNrnIcIXFb2ec4iFwQ2wAUSFT/c1pqDnKCn53H3GJ+NN/tzHSG8dQ2JQZD0
8E105OZQ7LMkweWFjzV8tVnPe4VX7S5qWkDqVwsiPVF77in56T3OZD5Svco+Re9plkZ8PUQZmKpF
8ruWvVytdSdBt1wwJj3s6nsY9Fc7BbmJe49haSonHwvxnOsOwaFzM+c/I/5v2j2Ug5M28mHCsBNx
T6fEQJ7R3Xh/wC3D6RBloLXfOCQ/7UtavGgXzOBKpxx0YGFRkk5zJm0hQYmGXvNcc0FC11TV8A/P
PwSynqV9xf1GgFovgQ7AzmeB0FqYUhzoGCXmvZDOk4MYsMfa4wDOlumMbQ8o0br1BIS3VbYHXHv6
hz7uPZ2mFK1+V3I8dEypnxj7sRnNYyS9T/R2wE3XwgcEXkeXBf16qiXUWXRB1bdgkHZqhxEvTNTC
hhz1XsBe4wKoxg7rZ0UClPHrlr6G1XaGfwq+EmMUN/IQyPWLI+Jd+B9ugFuyVQrbaLoEr1JOO7JD
92bk6zJX2HwUtDQmHxpDHpGERkeZJXe2r/Gr+RxrLNQbx4aDO2+G3kpAldmFWdyN6dDn5mSHB4ll
zPrZ5yGigm35HdAPO+hLVL0Iwpyyvw99MNBJXgHrkCDN5SsmNBh39xdGhlYChbxfbB1xA+7Ne+FJ
Gb8uB6YEv/xQa/8zqGGcIHcEriTGzsRA8NHG8YdqmRLEuiJCA4BwigCjc2w28ZX4+KE+IEIOr0Ur
Mzycjzc5A4DuMyEImrU7DzmXBBkFNLcyy37Id0fL+I9UlQeuTxbmRWLSdBaoCrsf+cEIzt7rFAd+
a/l+ESbV3XVjP/ODKJSO1uXPhYm8EmXR0/QqdLvjEIQpgSUSx3lDE+rehmTBjGf2xnalu7uAxD6p
Chv+BalmtDkUi6XQLBW10QBrK4nmLsM+UkYnQc1XjE7H1rFtVbiAmkacPIPFKsVSwEaaP/vT3qdA
JBXPV6KvAQFd+cg1TEttRdkP4MTnt9rIgYvZdFhRS6CcuIaPIPr2fLkcLosQ+aSR+5amBQ0SMLmq
qCrvWBWHTMXYowQQVBVEPmoQGQhiIebUbjJdtXBOYdZY44CtJEJZy81IadiBYi+zxBWKSaeS8axN
DdQ7/O+Yikff8wq+u8y/8rZW0m7Sl0R7DUODuazBSPRqry7eTF1PgGKhTAqTK10mLnI5Ih8AKY4k
wt6qIAv/znNqVNNScz31I6YhXyMjPGPTWdXxkLFya1Xqq3sGODtkcQwoCeZp+xhLEVKck6S/xUAT
+iZAOhawVUp9mwUHp0toJoQpg4j8VJKiV65b8WDzSp60XLH2KwGm2I45k0VRgXPgz93a0r6hFJxW
gLPlpKuJjMA1jXKWLgbzzMu9wU7O+X8FITdBi9KB0EpkVlxY5fMX45zOoVZCNtiesCZuDbKTRpZe
34j3Y6qfKBQ6tRjEuGZ7Jvu8YX4B2aWST9DcjCOCA0FvxrnSnINjdQ71mUJQwzlz7cm/1fJyhKsr
TpiBs4U+5at6SvCLz28Vv32kPX7p6od8rCqKxmTCQUguY5j3piCUpezMQMBKgWbgaFbSl0BWucXE
S/mAw75F4CvrZsP41i8sifuy2BGJd+ncMn587PsyuclWRb4t+xPg0AKMnxbSGiT742QYDxY/QNTr
Ua5T/1s6tUUtP4vHno+/iBdAsEwLEnoIsaqh3OpsnHQTDUwtdBYD3ddbNqWGjmDhkUZiJ3UvGHGO
CeaoiZO7v81Xi4xdAb7lhSKkPk7rJ/S3p36u6Rs6Wcllk3zydm+QyfKlA32fjtgtsGJNl275udlF
jQaCf/9zXoIvxd6RGvoSxkSjbfkWW+Fo6N30cVLdvgs3uuApvc0Gyc0WmjT9sJ7HnPmHj4kij0wS
oxVQeAw4NVGyPUPbA4YtkIMcWdngqI2CP1aZA3dLq2sH8JHCzTpliZnf9AXYBJ7IFBE46Jvm91y+
0gftZLCJxSXN4XP3GPv0y+QgJ4SI3h7RqHVRZ9pKvJmCzFzngRyxCt4VixDQr9ZygAMIqteioW5T
lWwc2rIU3NH7fAgMb4z/LFeaMGgFjwB1ZMu9Xsy6aUHk3OShAOvgWj2K8ntNKI6q7xXy8e+PuYX3
EXiS4Xi+oSfZIYSKiVbAxCXQUCnK+zoDgS8l+ir3Xe+iRKCvDKfMbffv+ejFX1lOkxfrSaynHU9z
BJRhuTUePXS5E63SXdextQBgh0tTrBHM12uM3FjZcpFjXhXzM0K0RsqE8e9kNtAri9KePfHlE90R
6G4ThS0Hu8gpwboTfKMfUHy/seZOnYXdPBkp+8W4cqTJYbtnZ5zjhu4OSjpuaINQ20l+FLyMYRk+
kML1AlTekyefOCwNhJgUqvI3hMHGFPgIqqZVbaSKKXUzI28jVUbmuoP5oLP44eutY5Ph1V9Opzmy
AzWeCIP348ezHqvyBwvw9YRRCsu+2eTfb5i9ejpIQXyHssUcxUUdrJxSsTHiDsQ21VZWgzhUdPaV
goXILDtOzyVNDJgjpNsp8t2o2TCppP0SWIgcHKF+3K5UZesbgZ/gAnhbe+iRidCYHOi1HjSDAVeg
g3ULu8g2ghdyA9iukJrRwx1NNujjurkewhdk9Na4IXf2/D5RzaKXuGXRFQX3O+cW7ebfUlz+GSs2
9JVqDBFuGPFCekUj6lvA5dvCvv7d6e33dezDhiIKEOa1DVr0/bx7r5ey1bOxPel2VYO2BixRhVcz
rngHnY/+OirevEhSpSB1qTZFK49l9RN7r7Y6PQeXCDTRPqf0MubtVBsGzc6USlT+xLPESDGHcyNC
xLqeW6SaDQaAK/TAOjmcGJMYXPkpLcZTrZtq2xQNaAPaX4c+6LXWCWd85DPOTKQKOhfJJ2VXZFIy
OVyCYITc5IHkr8blyIsyrrt8j9rVDo90k9+7js7kQjpKSwFM/khXMl5H1v8wXNzNS4vFasSh0Ok2
M0AgC4olLEf9oOD7lu/3nZqnBil/iU2oQ3CtrruGHpOzFyrNX7v7aYHbXaw43m6Ja1OnT6nh6BBQ
8Tu7M9Vp8plvLfT+7XT1bBw4L5cJuzfcSN2dEOixxu4C6rPyFPbkt0WixKQcqchvanBLv1sSOIc3
D4J5XiHFxy2v0oFUkgmRJLad4+PpKBf+OmhVM4FeFP9Lkf4AQbOMw8QtXnLqbMjR4HWuJM4ELoov
CtMntMRWi7yOP8oSebTUDiLob+ip4DLhJ7c3HKhWoRX+xL+YSVxfqVHg89f9S9rCoCgZFV+YYuzf
LBABMnWejSdMXEeqB2yNix4kOYuSju3iE1toZhs+upqJ3vn4LUoy2ZibPPeXYaoIGcViICtDZE6B
pP0r7Ik07KcxRz+DC6NRUq/OvN0TL11i7j8yS/a2NO6fk3HtpDzYVmM4O9vikzFDgrxCi+jMdoPb
lTy4VYb/1SQGd1pjmhQaKe1szpuZzVTroWNWm93bcP7qFemFsjTpW5ETSL6XIyfyT42buPhLLyeY
Eplt7T7EuBXtD70ROp1GuE9PUoTzND/pM0e6x+NHfB2Cz8YaFR0rf6HSuyQVZ8wO8qyjshgiqstl
y42UjsB07jVqgCruCbYia2oDJmsydu9OjY9D4zW8DC8T35GALsoIFpTiu99ObNHIvdzLq6MDOoj8
tqs56b6ifeLig/eZo4lkE4/YjiebylMGMCNf6lDUmhWbRebBbIa4pILm75isQPS4uY4pI3sg43Qv
hz2UODkwFn0OhBdqUPVYD+Y+aDwBbjxUEvHrddnxmYw3UC1yh7pz8ABT/MM8D+8eqBy0kVoMInbL
zaY+UAGaJdRQLhdxzPOhPu+vQMeJ3BsILQywYAOwv52E0ncWT42+N3xLQr4FV3z6MGjVVVPDJLNi
bfADIqJbCx+Bp0+SJqZbQl95cCR/zy9c/GIz8u3EkUF+4uKPWZxkMeonJ0RPZot0SQRk0P3B5L76
WhUmsesgYSbhau/1Fj8u+ElNdB5e8K7NIPu+TOx2H2J+FGkWFSPD+ExyBJ0rUX5w9lpq4yS08YXf
zmliRymS294azkTAxYddYpuNA3Un3aTJlLohTT9OSiKr3VPRg3K+Qa9t9IIY4G/pN00aRhBCNlZ4
ikIXHAjgymQ4h185LB1yzS35F29X4UIacbGos9M8Bgu/VNzLaU5ElTad+ImEe+RI1kvv5vJLRHZO
1rQCRCEJcBojVnv4jfGEA8W8MoW6OTRo+ICPjTZ6kQj9ZuH8MPz/8ymddYSoqOmzd9zW0YDPwK3N
y1rP6ZB5SZ4N3Bo7A5kgL3qeJV0fRm9wy4d/EXDvXJxBDkRwm8iu+X7g7VsQ30U3Gb6WwqZbAyfh
HIVA5njJcu79cHr5u17QcALbO435hfvGIBZJSlajXvMb4JTjUEkKptmplZr2Tsz0iFQkJwf2DQvz
QGGwYXgrEc6Fhaj1mcmwArgSxj6/On1xtShzluayEvgn/+cPDMv6pg/WohTdVtL/JdIfsvXNcyZF
dWQCbUhyJqqRNWmxd7sFqO33/W3eeY4VtKW5Q+aiV1vFcC25W1VS5vHDXtTy1pkg9P2PBABNPbo8
b69oEKWF7LPbvU4Ek3os3xyLb5jz6xok518HgZSvTphPuWZOA9U+BaZGgf3pW+RdZOQGnkug8KdU
4jjxGiknN9n05zUzoYmG74gdducYapNGcngp0paLw+SBftIZ1hexTKaOpnXnYFNGWbN4iMUS7M/F
ge0IoPPhFU5gSk6Ar9jNK6YjH3RxVC4FrYZIq3VvmDprdBxqgxa8zmItGMH+qiFIU9qgBQqp/XMO
spxVVQ7z1Zg4tmyxfEN8+slQqEK7slCw4YiOEiajJkkHJMTd0ltexVG4FeV4625Tfp+AGnzqFE68
4s32tGNh+jGiNf3cjI27+mYIqPoar+MME7vKTYrjADA/fX/8QvSvHbaj5NSd+OGj/2zJYPMPVX1p
7XVJzAvzw69lZIjC9gPMEfbW7Fa17Q404FqY2skJFwQu67dcglnAbBji3sVJF4vqTJGlRXV40HYJ
p6VvDC1SxHlYx4I8CpE/vNn9D5CuuW1BtWIqQ4rxARBBvjhuhOi+1DVgYviPTRhF0FbyOom4z6k7
xHMS8wYFl8CBZFSE2ULMOO8Jjnmf3r96KNJbLTtzdJTGU+C+mcdNPicAlQRwlWEREjmFRBoHA8If
Dhuks/44FTqPbouGO2xzF9ZzOYqK567P3kMBgJh5TymuWVI1oTF4yeOZMOktgxnm6Y0m6h/WfYMY
DcmuttDc3+vKCof+4xCkuVnLX2cIDL5yELzUEwoqQfiuyVQFLzEa6BKfqpuF0xVHvLvQvJ4TuOYi
UUY0k4FNofZTu9wbiDTNOw95XnVwqir5ZBM94k6REs6VQdqMerDeWK04uwUAgsko9ZiVSHKsh8AJ
hffPPBkKJHRMcRIV5UT9a3jpNFRgEDkiu9K7SUykwMCSS/ITNW/yH9d2RR6cDmti4ruIERwQFU4F
ZrLvUbwNuZUdasvl2l0uSHVB4WnEA6nENab9uQqm+cEcrm4kg3YcbtF62jq4o0o/xqvl4vLdoaoC
ElR3eCYlQ7C3uD4lYAHRzz+LQRkLvpzr5WpyXjZPCpIO2UvW6CAUe+C5MyW+4pGU3QXxb3qvVZ6l
vdK/xRyEbUkZ4GY4RjSI0bR9eqMv3jgbrTrpW7MTn54yOT4FVX4e9+Reo1whJGaZqaBnNzr2emUa
sosS/rDBbsHCy3mwWa7yGPLDhdlsSjqmRGw1Dv7U+JflvVCR0I6i8LRpUUErsPMu918COZnxfZma
U54VQuhkmTcRqIf4Vm8X332ziSr64w0uFyVpV5lS5UOsQZN+avXeGe2nAyVd9ndvas/M7mjOHonX
yMfdqV6Bb1HI/xhQox6u3k1AWzTdzuCOdC1XIDE7gIMsarqNy5xzQz1+avoRzdwh9N1QD8K6Wy0g
s68tGccVWNDvTKw/svfjYwKW4GdL/8XVorQjm+QCfKsDG/KReFFhHuf/qhXc4OmHciE4NtEeKO2E
oiKjOJGWE2nl03Lu78q/WUmHOm/jqoqKqyoAtxJp25H/EgilasdXauJcmdWAvUOOJU2vydVbb++/
Lu1H+nt3HTRfG6i7viF9igIbtCh8e55Hjst2u2N2Zy6bmN1U4vnN7vBOzS8LM/tifk90Ffu7eomf
3cTtR2QlufhEYoNHs647qnGEvmIOmRgZyhSLGaD0L0oOUgY6FOcHX5nzEdIVIMaIvsJzm8B/dGYW
szUNj7Nju8e8rQMU/W2+2R5Kpp+2liEpz7JmU4/eZLVYQ5HE1d2UHQfc0xr75eFdGTkBVzAGce+7
OrgnbixzfQP6utPF0BAdjGhriFfAkkrJKoWkh28gmwcBMLUqnw6Yzsk4MdTm5NmLdbcJ5ukB00BM
nVkaK18sNmScBI4KLynh6/noxbsGS0LjTumAhGz53mE4GOAnKNr8ScfaRlNP6LOYUGQ1C0CFmNU1
esmW46g1OCnaqK5jHJF/W8mSDrKR4Rj4qDGEJRTTOr+Dv7WU9Ks9qKY9f1/VeuEtzYV4AU/77guk
/6kjdrBzjo6ibRCSRsr8OF0lrKF0N/n56KRC77NaR09V2T+afBHY/ebWe/UxO4Gfv7h8EJNcqY3Q
NufyJNHY4cvASSHOUPxyWvIFYk/0GCIFokcRtVfEhzv59gkWzKqvHSalL37yjE++p5fyG4XLS92i
G6RE95eIQ+l0RZ7vzbBAoJqpncaf5ltOGo1HdEoXCyGutS5Oi3Tih0CxpsEAQPOk0ranQ//Ov95n
kFX2T9WxiGhETQKH/4J6ZbEhYi6ASiom6NUEYzrV6eJ7pBg8mQv8n0He+7dF0oNzwD2QsAYZ5ZFb
QrBtlf97Zra2G+N25oAE0MzY9kEYpSdiL5coAVblpiiS1us3Rm+vnLTV3wubH8s5BqWlakJJw7uG
tnnFLe2NTz0oCc0e77JyIy17gqJJkJBShbMjUtLNgEespJnFFbu/yAiUZ9Azr0p8N9rUrQo0HCem
4sIauoo0NlLckHcRAz3myvUqd5DE6ZcoUTRFX3CWERtAOj/zFiw/WBRaEytBHRL5oMF3diJ3KQYL
Lv7Zz29aphXVNuvHOiJTA4ADNTD9LPj6mU1fAlA32LGPrTwFd5VtOaSHlrTV6dYA5kejObay/vLe
drQCxXEFbn4XwQ1DfoleX6qBrQkWYk9jnjyoM0tKCnX0peOcoPkA7VnaNIMWgE1A8ymS9haVWU1j
SDqOO7Q+LcRW7Zv7P8z8JqNOwLU748ub4XsQGIrhggHhXMdmT9Skran1oFbHdBrNXbRAZ9y0lgTb
PLvaAerEy/5l8JveCMPEItTDmEb7yzYUaRUQDD+im5ALHtebF0sM+4eg2holvRpfRsm0GH4gxv8Q
JnUVM9xEDajzsp9OvSfiOsQzChMkNqvI8H6BtrT1URHvkuaTt/Z6d5ws1pnCGwMPEApsyIsAlLTg
jI+sbZxSSxo2Cea7yJtJL+GPinZEMQ0p0R9q8MWmw5+Lg7+IpQVWvpmIQjF5g95GV66HwmjUS8o3
pUJAJlgJlmwPi9ybbyim0sXaD0HVJaKIkd9su/qecAJYfakR2st5O56aFMvAvY5yMW42PyMngRbw
qWQL+oQcxXlHgit6HFwv2lPyN1oRGtMMEKPxOivwB1gH0GyPjxUT0WUjC6fv8wUV+5gdJT5dA9cK
zYzWKjqFFpXLpn5We9f+KSVBNpmLQbJNWba/Z9jT9GD3wnd5rP3T6m2bJI6oPex75WtayT7t8GaD
7g3JXNCuAdJcdRL0Ew1qRs8efMgAGw6xKgYarA9SKVEpZAtXzwvD1929zp5zTy7FD2OiGMoVUsqp
7LTtAPUI0kW0lEhBb1QA/9Qw4/Lc1AGZ71nOUpUdmbTSjoxM3HlXajG4zehVf+6Ym5GHYAAiD431
qNjjvCpYMqDOa3ODrkL6D7qusOgkSZoEx9h93WN1WxajfyJ4dZpCo55bw0f4iMTV0xhSZO0S974m
kwKoBKhXRO5F1NKZ67ofKFsdE7LSsGuQ5vrKxFoPWIIpTcL2dh9qG9oer4wTOHK/9PgPad8dJwq0
mTBYGzcQdRL5azSzHZcoPDdOqv03spKP2/On/U6ECwB0hizAFCuERzCrtLJY8Y/OVrEKjw4dGMrg
RY3/CPzyL3V/TyeBZZNeG8+u2zDZdu21c02qShUHPx8DBLdIYEYCwXM+3g8BDWXIrh9vR2KkEd2w
Xn5bNEPh9PyJn2EdKiSKvhUZ+VfZUd4fXvWUF2zC1NiAzoMTqav6pL7pjgJbMV5FmTRs4KfICO2V
+8B3jchf436D9P6NzPRsYkzsahPvPmWt7mywC6rxYE9iGPp4KCEjn5xlsTjzX9GDbFpUAdxiMlHp
zrHxtV2vVZqkXC0Cquudy804LvNgiBZCUtUEwBzMqQkwo9kivnAex3RtpZT2kXpLEQMdjK2mjJ3X
kNh7d0AY67tRsgHPCf1B3RWYcTZwhh/A6qCVMNcOPcSDYdgg2kkW4ka6FO8T+hStp+HYt/8o8z+w
PR3uVTw4iokqxP0aQQIJHXkRxc+vpERBrsBbaudmR5M9vSfo0Ya+ekxMMDtunmH1OLNNWCgT5IZF
z5KNlcW9QvZtWm8EI5D7jP/kCllOaJMPv8pBCEgeUbi5o5lR5QECqQbWGLjiJ2jRA71C9UvLuNIr
wn/VWDenouIiyw637jH7ecksQ4RlaQ8vUwHnUXwinRWpITt/xvpOfHa+jX/+Iy32RIjyDhHG4nx6
wKiO8lHYKyCa+HKB/BlugHuJ3vt/18rQlb+eG8pzPxABmWWIwplE4mCTd9YOvXkCfw9AqrJDPa9a
QBpSnD10V5IVvv4OWSK9xnhctJZZgspTO4pNP0InLGtjjZLaUdt4ogLfxuzxrJPtDZ6EeOTQjVBY
fEJNRqbi/wCkALPbxB4ftQk26bgH9KJOfHx06Sk/Ch63VVrtuqzci27ewT+v9sk9VrM5QVgEvgrF
iCnzzpf4VYYfL4HSCfdnBaMkh7W2GoA/s3w8QUTdTljF97L+BrCH1Ezv+ue6iPz1bfIiOJ74Khl6
dJyjRmfvcCUV043N9sOQ1Ux1sadYgCyH0mTtn6wq0VApvrfPwIRcbEpwNLSjHBGUbiCs6nMKuUeF
pzGNS+yOp0UjNQRuJkDeYNaIPs5DfnQm2/IT47LDXVFSD7qhlho3hqtFIzumAU4oOFT1aFgT7zuM
JG9xusHGzfh/sFFblQHaGEZH2cPNMRI6VdNG1JA83b/9o3uO76GMRBG9imioY50P91/MRh0tf2/Y
QpXtVUZRT4oucrUD2gSKNH2g+fV6pn5+PAfD9fW4iJ63j9TmLrVRAboiDoBToofAG96J8fGEe0YW
HoiOo78b2A7fIAyx6fa6FT2pHkS36JPiFzD3UkycHCIVnKYBSTl5CLkcK2HPfEylEjNn6UFLBQoM
IamEjFIhcGBuOLtn5sIaErZDL0UbebBfq9LSbXxeVNtySpugVPem66GeMaZh3/RSo1XcK4DoBWt7
4ushO10RSfsOaWFSywhTSTbfWJJi6Ec55PJl+pZgqS16IK0JSlR6kTsd480Z0HXMU/OVQaQJM5f5
oVr/He3ew68mOrNEpXdwPxwvKlliIroB0WxHBjTVXl3a2KKb9hR4YIpIDrw8TsU+PK93CjmHjo5f
yQ/lYP3V/gn1W297CKRQDk3ZAZgh2zZmTWi6Oov2npKYdejXifKXYVJSRACIzpoLt7vUqgQw4zIE
rLnvP90JY32H8LZCZrS0H1npzl0YfzlyCNxGBcDLuYJsMmIQg+k1/pL6cjtOW/O0c/2+BX1yc6qx
Mfwec5OoWvcNJFKZpWvj+tcOzON0WGZ2Yo+r2UxNa92lN05SQH3liCfMlKDHgz782gOzwNHxB4B5
DAQ435e4W+rKc987kZp5h3u6ib56VIwvrgFDD3OYtvWUnGQdipy6L442X8R+a+NCZUMxdc40AK5L
fT2wsqZhldLHrl7WAxTHWLBMYZjl7GoaiD1WsrAW6w/O7rQPTxsgLgOaebSvwViCNlQQy7hkp++I
JCmdGNkByFKPsC1hvuo5b1U2dx7lfMaJUDHKakOAG8TfnMQvKnHzAv9niVI0p1GJjzmxhRNYTtHg
ghzi9T6cCFvQLTIo45XVILJeMDCoX4PjuOZR0Zg4HRNeeGrEapQ/yi2an90So9NPpGms1ieYmIW1
TN/cAu8rbfMisRRHZ26ZbJqbtitMr8eYZ8+rcg/vv6MRpzufm2zKOVL6rJmDF35YYw3z+QtmZGFh
KlHri/Atb1ovWntVOqneaRrDjUj8thvWU2n65OTG4t7BcGJBocpnVaZ0DMMQq5aFMjj1oSm6xddd
onEiq0+Zje9aFS2M+bWvKGhPj0LHSX1zyXfGUGlbrZ0IY9Wp7tMfofgppVxZyEV2cWM0gQwgYoNm
aAiAHBHt8W9cA13OG0pay//IyBNpykCjzVSQO0YsyhaNQHwDlJlcNsQNr80KpMtahfCLiJ9sSzWa
QQlYpiG47VoowfIEertuulZrGt7xuXMfedn/VwFwq8NqpgN5iwakvf6Yq02OHyvHjv2rRVjQgVIa
1xiFrObFzy7IfDj2gN25unv7T3qkamwRM7qgQrdzI7V88EQ2sGT/3JHNn3A5oegcUeBHp5TIB6uc
1sNA65Rk0St3XyABwddBdejoNr3SnoNyj7+MCKSkB0f7zmFxUzJazkNpnwAkwvTZOB77IpHiuCZy
f/7zm1sT/XAiLNsI6pL1xOk5yhit7uiNEvcpu16NpJwYGsDZz8CAZkkbVHZq1OkdZRlYoOGaZQfn
uguCIaTfCdmtDh5SHIJHfPKc57BbJNHTG1xmSNJy5HjqOuYa7ZKU8l4x12SAAPzL4pkrZ2+kfMvS
0NdFhUA2OV5EqYs/0iM9QoiBxaThv7bzbmHS35Lca3P/JcqSUKITKlLR145qYhaJoAyNhAobPWX/
CHqD9x9O+BduAZzp/m1Ry6QQHjM/3wfamRPskbwv+kxcuz8zEtt3B+AbcoHKRFCLrNB9yAcUrdm1
O/JzS+UkZLfpHl0yFTtK4uz33c7uOYpHnk6M5CHM+MEnaHXu1IvGkMdVjGJRkQe5YDQb0dHkhEYf
GSnAUUDU9tOhieMb0B9GDRycS3XbLeveJaCgDVjvJ6vJW065+E8KMj1JUZNcc088J7kE7z5dxh+Y
3fXIZzU5ENOijXJxsOnt7UkqtOk+D53O9X98IRZU0l35PDNFS3v/mt0tfYqpYoxIpy1mfYr9oZgr
b8oHrZmIp2MyqDDv6xiCzuPsEO27prSdl7tCs+VaGMiZj34k+pAbhqGPYMyLgf100vLYP+lbzoZI
RA0QvkJsuEJ1vbwjlaEi8W/E1Q9GffDrmt4noQPPl9yMVU6lFXFV5CpbBQHsKKa5S5y9cYNbNRB3
2zZQEcvvt+MPKY4guQUA6QplQEQg68o1xCczknoelp4hyU1EUMm9SSRMlQppdtHM5tjR3EQ6mlpM
CFIGERttdSwjhXWJ4wDzgDLe+O1c4wc9dqVkzGImKBYBTo/oHliKYW54brEWaaDzula3YholgKSr
G7FTFioBHDkbE5CImtHNpZrZKxLHKaChwUSqlNl3q/u10TWXg+v7top3EfpDyIC7O4a2OlyCl/J4
6+mu9R9N+BPabwqw4rIhJxBqelLnoXt9Feg3Yiy7joQWKizOXOiiN8DZ4fQegg/T+NmOiRiGkdu8
ocaU19o/l+b233Lsvse9C0K8U69pc2yrS6MGiiFMEbQzmXSP8s0p0YUAKIT2J0AG+PSvoqUGAMVW
8wZS4sbBRUYQwFUGJjhirVlRCL2GNZcewcyWDrwpINW7DZdxu3m6VtI7rSNWoZggfvvxhSV+vc8E
8vzlJw4EzK/6XxtDfS7Gzinjwe1RO0F0d9MzVfN0T+2zWj34quHL8cFQVEIwuWcIA05BbChHDnIk
V/RPSrztvEQAFK1G49g6ZVoprlCVarkZA4ZJaz5ghZUJ0OJnXqpRBjIb2E+DUHE6q92b5PwOQDRO
/n19xHgeNK+XSsB3rOmxMT0XPWIOzaNbK6WWEmJn2kH42xREJ/AZVSuCoXEmLSgYs1eZSyiqffEQ
7LxOW1kav9+7500yGe50Ssc6FBzf+mQztG+f+pile0NEZCMcQMDfXUAyjT4YD4revLRkq3ZD/gzW
BnKPmI7ERLytdRRfZjtgTlAom8MhTKAyppB8Pl2DjMre/bJuevZGcXMRf/nvZEvWSaKvnkWSOAAo
tQeGueaqw4qPjmEemOVSsKfUSL4cb348ktPUg02QHOgTyLKb4BiH0D8NEiUMikZZZo+vywzByvD4
bYrzvC6Fp5+hR6Qn4AOW/tXmq3x1WcTQnCFhBimTu8Nv+ZKBqsX65baCtbfNCgW57FMI7xDbZm2g
jfczpHdG7iFqIyN9Sj/CmcxHO5JbpHHeIzBTTIORuWoF08QG4y2DTc1H1Y6yudBsNv8IMNmjjAgY
RxxvcG5LsEWf2wygEwsbPN4V193PRnTv0gAJ9WP6vLuIfJg6czA/ZyHM/1vdTS8cr754zm4jc8z9
N/3GC20y8j4p3htlBXHGYueQP23tVIyEa3XKNb9u2slKO1PeSY+S6bBPTwaoAuQOHqZiuKn2h4rx
DB0MKVkVu3fNDAgvf039WvbJQRmD8nIA2RsfEfzn+c91EMF8BNkQG4w/aE8hvJHreBDZ3ZeEe0HW
59U83sT7m4G3Jd4H/CMgxwaxKtHCjZYR8sREJEDzpvoxheIRMQxu1R+qI5U1swWufP0IiFX5U8WV
5eIdQQsuqCNZkU26ikxp5mYPflZQ1Bq1u5bvrlkOrrOxFotzHa5uHS7fGsGrzoNV2TBLzVnBivo1
xuYwS9ojEGdVJ+xhbrUTUeSgk4WzmMl+IzFN9oS+kKTmh1q6P/3qpmXGgwQaaVwK0OWd6hKHNgiM
7vfygFUA8jvCQqlV08ySrOnCua7AgHj9aRpi9AOLYvQuOoN1EX4erPEL6wYQB5/YcELu0aVxlRm3
moMM5evlBsF+1AGDabphI9GDdh3xpngxSoFeFxiKh0TmNt0NC4fm+HAgbWh76Np0S2cLxhmZ9+4a
aAfppti/eTD2VK6sSRADzBajIFjoMWmkX0yxwI4OhbA3uWtBKK1+xEIJKa5moGqFf4HzxRZFH3aQ
/G+opZikjI8agvTceDjHK4PMsLxvzgYuusP0YtGzwbU27lvqepAVJYb5d13WTKjDgtdfdSnmFWWx
MxbDh+7vGl4bRuRf6AhKjfOG/yVsms2KBdJEjGj+m+RC4gvN/MvZVS1ifaXeiW5SZrO3aq5Qlqkb
cTQPLwCVGzJMlKGcN7kcrGfLYJjmJ9C4Kg8IRX1ksUq1zHJiDNabhGjqSGLiik8EJ1CnQ0taETUV
UkxaE/sI0seri7hU0rhpR1/FBwyhtmCjfzF8+yZQ9gZAlaynGiiRpcNVdDvIWG9kwQwRPaoKkzyU
RAvD+LUMRQngrGFeVjsq9H9xZWLQAltj+uarc8TOtY7Sxb8ebd8+fJ16vAUrRPkr20kG7Yd0/SD9
WxStXuF20/25BLEiBxWwUeCGryG369yoiB570gpjLl+dl1QsCyZg/mvv/EFR99hIyTOjYB16W764
dq2/uHLPh1aiOyY4/imTcifKbQ3y03WIm5Bgs4aResQGxmuDE/aSNE/orZdzYMGz808a+6+vYJYD
4/Z7Vm9/zpb/+w7ylC7gAEanZNxunSrAf9qtIbo7vff/nosUEifT3pWDRSc7pVOn3LyFVaiFqC0W
yGHn3r5uGdCsk6oa60DjVqDLJUM0m9vfRx6AoVtYGNEqFRD1kdHUIyjSPL5yNabsydy8a3n5pikL
h+kBXS0ZlAK1kDgWBlkZ7T96PDfypHcnPZE3vkDXuGO2DhJMGV4ndXVNdgmptilc8L4DOyIjNqap
p9TH43eWrAZ+HIxllw4S1EMHz9ypOHeCjF94zpfl3bF69JRtJ9RrgtCqHUlSUjfql1VT3u+9QPFc
q67dPj1saLKUQcaqY8HAuqH5k1LKAL21vMhVZc6w/TbcPUN8cZglol3Lf9hGGySwj+GWLWzYVRu8
+/YN3HHR4RJgd/cZGpF4Yl1HYqzbMhS+RYUWgqr4emxtznHQLwLxQQ2/5ZVmpnw+BfW15WCGCxSb
+QbbvEIs+AxwbKyJ3X/Z2fsDdXpdzl8E0Qyqgsu715VaHGxLNA3FsDmNLJnEk+A6CjYOnjYOQueb
UjWPFRUQCAqKFX/qopA1VIxrPCXkoMlbN2jKw4c34borIauPw7XjdCL2VB2OmFmI8L9dcdmw1WeX
77IICr1DShxZ9DKlrdqD8A+8RlCz1h2E6zylYriY2qlWZQr4E52gEBxG0IL2BSJKQM7Rb1/iipgr
Lwues6eXGDe3Gh/btoGHNl4DyL1weG1eKunmzPHYQnZXkukReVt6aKPJ60IdSmgFYjlPip1a2hO2
oijnLBKM+P3KuB1gRI3Wr3JzBqCP+eoy/6NePftdPdIwdRBbPzkHkyGZ9g0fpeVasNOuSRXQf/mc
eIRdCOkH86DkjMrIO+OK5PC5FX1GITGPqDi6pB+LEqEwQXS2cy78oNl8yMV5BT0KFSPVNCq/3wIZ
JikWHj43yGLjm9RTDaD2lFA/pc+UH2RRosL1l40Tx09Wxf3HaSCU7UH7tFBZDDBuV9ToFOLq/l56
bynJVs0e78AJ9amt8M1aLL9XraMULBwxLW0zr3t2w9HH3v303C5gWmG5AtXdfvD9dCwbK0O9chC9
FJwmVgXA0aemshzm8sMjoCGeRuNx9+wo6bT6KdjwLikDEMu2buib8QGAEbz9Ic7VCjVj1TwizFey
17Yg1/xYwEeJO/mxJl1nH4xwRP2vV7CFGiyGcSEa8lzJpwa/uD7nllbU+ZGWYN5o95VkqkhiEExl
eWNAGeuWuP/9YUqBcyMxY7LmWoqz8R8ANaUmbmQLlSbxWNd/zTlSMXz6gjShpTfLSSEWZx5AsKq1
CUrgLzhiFpktGw+GmyxfhvXbmGiG/hxyXvDq5SKXtesWFrQnJMKoH5a7igVdlVXDuNiJMv7Tr/T+
ksAQGSeC+FakjTk2G81ICBf+ax5M6SNkqefVg2G8NXhdZTormVYNhUEzBjBG/X9ucMTTaQJLwz8P
VLY9xsTAEYQW96vX9sjNTmijvIuGrH1+8+ckA4kaeGO1TZoAoJ1pRNZQd5taeOIHd8ENLd71jp4e
e+JIQx5y2emrTyrzPbNhoRyfWiBxt5xZmz46QcJ2tgxL9vVucfEx7Eg+ZBOfvWl3hvSsyIn0ArJf
uleyEE66x97QlIt4/kiqHrjOFNtF6ib3nADjBhDsR4yfefqWnCQPcYn1pcK0yKcJb7GmZI3BgGwN
M+lnvi+J7CO7WNxmqQF9vm9SvN1kLqaD6/21u18Yq7uRRYgP+EupFWO1GWnFfSTg48gR2ngU4BFc
eSXO2CgcaWklBX8QeDJ5yAQJxKRjNvSvM278NuKIZwBw5cPLBMnwjB/6Pq+A5wZ0/LTAr0ZlLiF1
z31299RDtttVlGQzRNx+tRgO5ySltMn4ikBivcmu+HZ5EwMViZTR5zIbO9K88mZFQTbcp3fx02cS
ykCnAWbl+6QH0aNwhY+jxuO4lUVUQhQ2yWHWERs6NaOvOnDgGdwzFwBDFoZ0duRM8GF1A6AwHwf7
BnXk/RKyZOGvfpu6xRkodLqFJ/B+Hkl4mu7fTlLQTxcxEcQMieNRcp8hwydZ+0cvKdo7arTkIvfY
Typ3cmQJA4RFgoycKhlHs8cGui2dy9JVhdOqa/G0o8cs/VLWhp+SC3px0Wsj0xnQv4exL05/u+ZA
c21xwzwW0owmVcKFjBTangSjNOWFA33f+gwGGm58mPMY0sh19kSgTuB3xtROdMYWm5f/0KiLdXvJ
JOiS/inl3XDKrQ2/4Ikoi5LbBfZrnu5AKG0yO9f8mtVixfJA57ZBRWqIemEIt6EgSex8paIF4DOd
aLK31UGfPP1QqGZZr1DQag+FTf5GMHucba2wucs6nRuIz04neuscEsjxiIoiKbliBajHtIg94fzC
QB9/T2d/VPc3AgGAKAUcJTe9S6ldra2892jO/Prli5n8Eezy+EpX/d5BMiLib9fr/Q5WGiN7RsRP
Ew2X35hW8nsaO6x4g027se6HyIDUwX2+7RoM9v+rz3j4pCNMRyqiuFaMhbsmBB7KeKC8j/zV5NXK
aEqAkKqiqz3qDk89YuXH6DUi999y2kIGduaFLsJeLWCQXG1UTbm1U0FVCDHOdPjhQsqvlph72KLK
sY+5wscBVqVtfdWRW/k71OCBTaer0IFjsJRtIDS0QX2VeUoxjAs57Q/0fHHDBQkBiznU6tz9CGDG
cxxkh7Z+1R+nLEaV2EfR1RXDgioTuvNWLClSdH6Oie4D5ApNHfhoNzUurqwzp7DsNmQZzOPM6fVC
IieZgXoOBSBQhICnDwuqKAJii5o73SKSEM6qC5fgNM8jlBJAgq8SwqbfJnxjCvmzsb0tc8UaUGvV
LcQlhZohecfryKpDw/nQF8Cej25Ba6+pb1JuDuL0ocPgua7IGog0sASlKH/MiaMSLa6hp6oJFIO+
aRrGphMbABBJAnfQak72fYuukpKCi7q/JPO+QFbJNyugdvyakmob6GDI2czPAHnb4Cq2uIrRdNIx
TyORO/TK5mtqaN/ad0UqHPbQePDLMYTNb2E/j/qjs6Al5VNP0XV6JGp63nGIEqTxXCJdRJiNBIZt
OqQtijrKnbxEd7kNWIMkxtGlxqM1srnqH6FGV32TxMnkzHBz2yvnyKXX3FzPJh+cL3J3va3ey3BW
RYmXaWzeun2FL8TqVZsbNyXBS9HWzxZS5a9yNNFzXDnGSARiHbq3icY2D1wS7ZxLDOdcmcUjIbs0
5g3rrjl2mZ+f9WHWMJcWCM8WDgvNyisvOTYAZ6DJZAFtLGg9am0oH3MJh2pvYfTElDMjQUxFh9+i
hTJbVCwjz6g+Fe63jF5AVVkP1iqrT8nQp2v7YuFVwgPNKrM+8Ge68Klu/Rvsf6/8Sw5QgYTdFAiE
pbucZg1KsDoDQGdGOrQ5ArTDZhtN+S7xT1zNRTjgJUxTdw0zIUuMWJPB7JrIKLb2YZymw4hpcR7Q
C5QZ5DeLRFoc1S9H+6PXz56E6r83hlQ60X1X7fcYRhIPp2jGETGwG2P2Ll73rQ/53NbnTSkniAPj
YIfOaGFIiTb2elAG4XyNba5xbwxxRQV8/mxr7YCilYvWFPahEF9wvcheMQGW5Zu2ZJXCLroDClkN
0dOR+3+6xrzWJtRpTNJZXBzazHLSaVCeyFpvHgHkR8ZUI5PKHb17Vyse5RGG78xrbv2xuEQuskiL
H4AVuz5+ckMF0Psc6Z2AZRWdEqX8aXStFzB0Ez7UI+TfG1c1ywUMRaUt4ZgP8aC64cQdJtYKvrQM
+uu2rBpjzDVD2wasoMpMuIo/UUMSOjXRWaMVt0W0m5ucF+soLv6C3pE9c/9bXkuxNd1EDUcNC194
e3N+ZeTg4bo9gpQkzYn7hrypv7kALhCJNLRnFElSZjju+G45CwgV8l5l5SKR6tX2j+N6661OBvWK
/5UXD7/JU+hd50ncSzBKbmGyZ5sLTt8Z8brdJMoieVw7AaMqT2dft6ytMorsEF+IXT6L2E5CBN/q
EaWjHZ5UVF2b9SsuUaw2dq78pgOZUvf9DoSMWu//mhgD5tMZHEx0Jvb1dAkGa1QAI/NM3y2FGlCM
TVAibVPjv/n8Z1dZKGuZ7J6bxVYJBoATmVgorXAzx9ufm+4m6jSlAFXfMdFtejiwAS79FVn5yUc8
BxCMe8A9e8TOHVvrZp4IR99vf5re0qy8ynQFSOX7h9Pa/RrfFjhLqQ7oRetf8fumyYU4KhfPBjq4
/wabRCZOiByFdBGmn2mclEHuhRAyG6arojTGeCBCeCCFuxDevKYAfRzbiZUbM3LyBc0/FXckcI+Q
uU8VfsKSk3YUZNedoC+EgclFgva6m4nUIMz19qU13TqQG47eGo1BLd1nWkDoF4+pSYfRXUdIN5rk
PFoVbtlJ041gtz73RXPx2bMfFSCTvrZkdd7bOQXhduwflLhcJIHqtB1T4lMGZ+uwmAGOu63p9eBS
VDX2mrbrzHD6hp+lUbzWLK5kh1n/neZeKyCEZRZvwixz/TiONnH63nvHbSSjUDjFzghvYRd9e9lq
E0eB8OjtrbHqtcRvBcUu1OGXttf5M9FNGhpg2igmDFeLfjJKwMb7PBwAF6cGqnBHzh73K3RLFOtf
2XgMAbJVa5ttuAL/XTL9IE4aNBXsye5b4rfwsdYkIwh67SS3JDcJpxpeb2/GulwEwEVguzjG9FMI
rXn7FvTgC9sgBB6KNzMyhtsY9oNF3DQ4+D/+Iip58wV2sgbR2ua+mc7sjz4QmsVUDs7LUp1dliCB
zslb551bU3tXXqGztQ1yNo+C1rx62YATPXzI0CCXcKje4qCSGT+Yee/bhLgKtchVYgMSB7etoDXJ
z27kjIs3AErCFrgR44U7o7kpkIoEKz3K4zBZ+lWqTDPmYd0qXll6yzTpck4sfgGAekknJ0HVedhF
F+cP4LcCHF3pVHuw5fhg8467GdF7BazaOP+50K5qXAGzqKzcfeSf8s1Bme/qNyaI08XzK+OAT/Ft
f9kYumgeam7ZAi2dcZ109cfrtfZ1QhgtGFTNk4slMjl40bZZgGCIruZkM6aeesq+eGpkt4/8tXzH
y9/yxl8Jyifkre/L7kFc4i8z/2IdqhCCzJ/eLmnOhkNpJVjZZ3z6yklfqJ6ZOjBD2d1Me+BEc8Wd
EBoCbnkS2LFCnZiI/qgSmQr0vQOrG/fCbOYe6jih1trqU0rJi/JsBmEd8gkiVQIHH12wDK9LgoB/
uHOrhfqhPp++jG7WFUc/tI9YClCedZMIz7LcQ8L3Cjm2r5MYQRr+/rYR1m5X51+xn8+qRKfMSIYg
ZhuKJbsXZK+1X9EVxs2AkpQolBTtr0UGBGsiF1Y9aH744ROu37ZZsnP2U3MPI1pJAARg1NcnvMMQ
sLbY3DCQ1WPKwgk7rZMRlFxtd/TIDTV3EjvdIRBqdpycLkNVU5cmKo/AAM/zjaFyddU+ZjTErJha
aC8NjJ0Jyp868WVdEpr3PpXotPCY/2ce8d7sVpDSwPC00NVg2aATkGZsEh8OUgi4yQ4MYGAd//o9
6p5tbHZY1YfYuXqB0E0ZYPguR/jacCX0LQ7Vw49FFfaD+Pa7kCh568XLknB+1gK2vOdw4SyHH0Kb
TLDIHuKlilbv6m6W+4a2FpDyiCdcyIhnUM525V6ZzUmHiVcu2J4plgBuzrxrt2ReelchrdoL3cpD
x6cFGKp98LRUHMs+SkiC33srNBhpainJQi69HIUFu075YS1nJySu5rA4Olcn7jL5tYE9l1Owd7iu
rEthyWPSEgsvafm/pA+puGWAgNGcJQw9H3O0gI8VUg1ZiOm844y2ojeZfyrY9FajfZJkQjsdkblM
tqA2on2C0jWU+msFHijBTDd0CM5R/Z6pQr9uiHDVtAE21uB8wDQuDAUptY/t8/FojLsxm+ZZLbTq
sU2XC9gS+NkgiUP4lTaF0jlfL2CLV+qIc2uaHK1s6JovE3z8ROiOZqbq8QyXCB5xxe5azHM+yUnI
FhKVmv37aYc5MGUmbaGaUt70xTB09021Wpn/gIbbSmkEawRfC3O0QK02DMgVtA/ppD37I3eDegvO
ZrtaQskAML0q8+BmGSD26ZqNycVHGiSDYvzekA5mbsmtnJQwrvjiOm0FGF9k9sSuEH0DXQHK0QUe
j9V9OoTEp6tFZBHrb67ZyA+4AnjwRgFxILIPdu0MLc/v8bqcOJYZj4UjJGvVAG//+XbM//AMl8hV
Bv4596fLz98e8E5s32xIJJMJ6YVStpm/cG0NrNzUx9Az+a7BhYYTG/nd2bk34t3ZJiqEhR36vokl
/xC6sFFIFwAxxwzdxYzpzZHCcMEZ0kfoA6fFX2X33L8aoS+x16OITBzVdjnofCXJUMlR9TSnIt6B
g3LdIVrhKufCBCnt9j+aD74ur/VG2R8jrC0rsFWgTwowKHLmh3atBGAVt4JGkMXFjRhc/K0MWqUD
ZbPplh1AkWfOwWfF2dKiNLs9AKeyHMHYvUy7TGWRwb00hripjrNO9q6a1/Tet4ilv8DCpoj/8p6P
bD16L2nlYbCw9nLZbVxEmlPx1srzldrS/ep/xQ1kMgKyW5MAMx0StS3j9+25iMw2/i1SOklnJI8r
FOqPx/6wPoCCVanQ3e+z7lpXO0oSMAIbP1Jl74QDhqE5VICWRBVwxqYtgi4weCeRvw5eV6ab/bk0
r5KTuvOyCPJwXi2JnQy2ai4YO7eJ0/LUFQxzNzSbF0fuuhBIzko+NeQwssEJxIQsztUWAVAVoEZO
QD4kQcqee4KgHvMJSnF0iwWUfh5t7BBhGBVz2K3zQ86yBO1y71GW9bhfHOfxEd1wiOH3Rg/qabKN
kAF7L0Xz2kEs9sKV4fNsbIBQ2RBiQzURPR+y1MBv4WLeA+nGUCW1tHE08kjkMrFyXwPu1oBVUHqN
yqE+HOjJs+QLGhzEv40JZAb9MwgX4dof/raXapDCPlywzwPYUCT6UJGfKmb1z9d3Q9BDVWYYaCr0
/cz/RV7nfSeC4mG0nZ0/GxjrtM5Nn7KkJnnNVRBqpsGBuB2rEiwQVviPpcL6r82EZsCJIYcRJY8e
jaLSiClnn//cp/q07ZKD7keEGt6F6JMSF2ElEebb5LvWn195hfYYL7Q/r0hpG2I0Zmn2g9rNbb9K
9TwH4QU/qzeFEC1JmuoHg1zSV/3/WBgD3nxVufPkskgeAsS5QvyC3wS8SRA/OoZMSqURzraE7ilh
ijvtQPeKItnnzq/+6nbaud/6A/RhLHOYdyGU80gecAJmAijxoV6ZucJH/Zar8sVTdrsGCPev7u3A
fRIoUySr9o8sWg3XfnJdkyuhB1lJrnXhMpFDRV9DR4Iwl/1M0k9FJxx/j5I+eQtOs0e3YkUnN7Sv
YBbfcXjgpvs0CG/g1A6mRk1psxOMxN8uiiM/oTeoDXw8ym2l2enQjeJpEfLbHZ11XoZ7ogrlDn6E
QnMIgWMRv3ovFlbWajGziyrArmlHFC15ZAH1ii39ViFj3hslG5W63CRPgqkTU3Rap6wZ3fCHSkqO
4+utgIOum/9Y6uALdVdIz3uhjMB0QPMxJmgCjtgx3eSxYpgvmSboGuGEgAW4LTaRVa55nvWHKGPS
0E+61mageOA+uqazpw9Q2ZDOesLoZqFzzZtxjHgj/h2bI+jRDdIlRIfbP0qr/vIYLGIzn+MblphS
Zm5uekKdtOCRybQhGuOwtr0Q3sCCoP8uXucC5Y1WKgpZ8x1dvzwIZQgBjfnA2dQlRasA1Ijyf7/N
tYeRCrPJhoWgFJ/bdK18YT2RFihnu81IIo8n1VXwA80X/cmHfk5DBxb52h7mJ4VomuzgqdGc2m/+
Ix1ntHm5XIY4LFfgVk2qbnavDdFGTiGbQmpj7Y0ScwYYkY15qZIZDrf5C+nmQ31zymzJSqF8gWVi
LWncQ1T+1Wd6PKiHl1ByllX+3R172Tyep/KMihNehv0iiXfx82sj/xMSimT7UfcQcMT9PG8xK9S9
xXZbBpnTHxpafldPstb67MBbWQP8kh1uRYjnxzRZrcgCH2w6CgeHaZVv8g7WN18NHfBoaECXlUgC
3IcSjtY5BzH8NBxvbOHR5yRlGT/4xdI9ulKoRYl5i5TVKrQ6FjYiY2kkcTWCD0svP8Dr/pkF6R0O
r/+F8yF9GuKg6cBJQBTuD+4pORiaqzNwPODB+1DH4jTz3oGk2SNyHopKdlUDz9WdbF5gMg7JGalZ
W+dwAiYZrV7rx2Lo2L1g8nJ/o9gCm4m7+SqGrz9kTj3tlAVU0Ds48g30JpR2RWqsVweoGiJarAA9
oay7zGoj/KxK9Yc8zkqRRGNt1wboU7jiAXRbBRw86/JYAktKcetQtGMHVYKg/dEPmUzGwcDB463y
HfSwdf2BEAC59e06/81X+hWiCX0V9arPnEy0lJTYm+Q2y1cQ3S8rNoPTQ0L/BelJYuc6W8AgykVl
21aYX+GBkWedA4KbX8BFDLuFdWMCL5h7tiADxA0JxA60lCnZLuBFDfMDcPCWZLuxRqwEoXbXrFtl
bOOd5Tf8VR5KTzN53xMoej+V3du01455yUBY1Sj/n0G5fiKVcK2QKyuFdJoHGzS8xVLJ5Zc9Rfyp
TEl4iEiKA7SN4dAgjmDI/hJu694RIBLeUoQrLVidXrU78FDLdjB91qf5cCwm0QmGoM+3w8KlnovF
zNRA9jzF0nD0sGswDIBsmKqA95OoNKjS6XLju7uWsJJdqBuUK3NUY+VJAuhgB1DW2GYyw7aXs+2S
Kd4rlRlKMzQ2xuArkSkZYSRuvo77X7TbKcelGhOuwxsCRP0DOZKDznMuSxfyyq8zjb23ZF63gf3i
tJSOODw2zqCAGI6aCf3F3cE0RXxGVZb5KmzZKmMMUOyFhPinTyUu0I0J/zVfajF4BDsXMebVG0PQ
LrKGeh6N1VfGqeux0XFEtmnDs5U5vZ7QMi//O7Okuefjrl1OjDudNUTmu5SCeCBq4bWXQA6wZqPx
CS4d81UgBYQoG2F7UdW9076Ys4yLUVrShpig2fUAe0Kf5MzXVFMMd5q6Hn4HzONAiDH7yun9H2F3
7Rnx06Rtc8ZOWneI/7JsqXWDuNizYvBjm0B1neSzITOtWdGJKrHZ4bCSugZs2YaqB0vAh0uGkQoL
p1X3gQbCvTgyTZxT3OFrOrNtVLC3s9hr/89g6vwkhaHfzjNV+/uK7YpoYqSXeaWgzXrdJGYNv7GP
c3lM8qJtJwRwiG2nEHXKt04ZZW/6v4d9KCJHlzIMKvS33z2JpuY4n4qU5RPUCFhp2J9UxSeZZiES
Toe4CJvTzcIUhBf3gZWuk/+u8bTVl7YKR1BmljPhvtIgfizgX7F5iNO+NasfaYvwx3bbYvQ2yD7v
34xXqMPR7g4TC46MDH4/fRiuE6SJHlwkluGPfWR5shwAPhEW5cVy5/xpg05nTaAkL3pJiwrY91Dh
X7k8yvMTsI7BlU5ADiFBhQ9vjd/KPK2GMQhjdBTl/REZ/jr92bJxcqHCbMXOCmfLfs5gDw6uF9Vd
dXnIum/h/E1LdiM9IYh26Qf0xOozsJWt/24YhbdawhIm82f2gbeYXhY4Srd6mmOd3DCA4kOXL9Lw
s8AEI71Bck4XwXkXXTFj1Tt/WWlq7kplAqzDmeQ8WwrCPHnm22el037YihhVDjYm5yfZgnnjObXi
bbCiVJ7Kd13KEukvgatFO5sPMX4PiZxvYf1IjvCnYS8IHkJWISB5ikBv/gthE0/w7wKuasTaEIE6
zKIU0FxK0BhfR+w8hzCw/TN5z+MdtH0+ozYrrCedlWqdlFWcb9COJpGsB49o7h7XRxmr/zXbKc51
4E1W86qh2v34nZn1AXLz4JJZP4uMlinm+QGlAceGmvtUuKHN6FQJ8qm/MmRcuI8wN6cBdstwKaWU
FOWLUtxgY34CXGyYNQX5J+ou3vJ7+jKuLwHCVi0jfkPHgLppks8MnkLsbSRZFR+aZIUEXxXvuRvK
7SMJHxjLIOFC9JPHa0vffDE8wVFqsq3c/EfZSfdEYrD1QxS1xEy47pg4Cj1s0EqXUphx4n0GMjzG
BvKRAaCHVkvoa41DmWuXnOeUDMax9tuUyLCPrTMcs9M911Qxa56aySg5g0w4YEfkW3Nulshw0zf5
ltYGurXYLmq53kFRDGwW1ycIal2G4iND85pvi30I1sYrq4PMogDae8AWCqH8JXoWl7kgTdVKRF3s
BgI/xQ3MuKZOECCoDdWFYIjnFTXb1sWdeMNx7DcweBht/bNnZafxyTwVyKHC2pgMKsY+IAyPHear
8q4xIjxjhrfnIO7Jx39d1LjusEolY9xte0lzvHYKs1QpxnHRgDaui95WoJwuUdmE3RTCAFJDFxH4
h9P2OyGyrT00WTuh6e5VRMH8bDd7IYlc3tK3G0Iyxcn0HjRafhX7IfqSGZN921EmSd9VWoMFtDMf
ZxBqvxuk88RDZGbBu5wpF2hy1LerI/zBdnJNs0/54TOaodPkhNesFQuIWPyi3qDScHaV81csIYGP
484sHyV/wvUrmqpXHjb9oXOMx5SKi7x7lg4Q6X9Yv9s2We85dzLIF8q83kuNDupXtGAwQjkE0rOZ
Lv2UeXS+QvBHmF9Bl1W2nPFl8a70KPA30/9liDv6mwYv+/p+qSv3tmh9aOfjkAqjpzHq4EkK6f2I
V/oN2tOmV1kkuWi+i9zQ5IrtSYdenSastc856sjkdbdXeBSgz1ABYs3yshzxIahUCwCo9gN5eLdE
KTL8qXaTBU0Y+T9o9RTabbfzMWGwpkLfr0GAIy6UlE4HcQ2lEdJR2+ERZCN5fDZI3Arwtj8dZ4GD
ZVaCXjDlTwSlY5C6lGU6Ndk+2PHyq67lIjd2IpokZXrRwnQBsjJdQS8x5czHNWao2dOHrp7u1cW0
cS1J917rV/5mQkTokDcGBK0N3+r3HbotxwNW4JodX6rVOodEJNRJtX37e/uNIyWp8FEdRUmylEGZ
Mow1+c4ao8DVfZYI5Iv+/CfPtdKkb+FlpwcfKZAZQK96gWzGfeKrXN2D1JSwwDqziNLudexp6BHa
QwXXpXXv7T9zNaBg6v1QkLszJqFerEYn77pV4xJi0uw1DMu8olXCufdOF7lKJCqRDsscJuuttY+L
7u/H++4UHeQ0g78Uh2CMfTCVFtQMHcphUYAs+hJmfdkLNTLTIsaGD3QTmJ63anX9RmyFOBi+oDA2
pRGVScWTxZSMpfYBATA1rtEZrPrk4v0RKtyoh/saEOSZt2D7X5p0jO4kMzc8oJekunN9AayBdfLM
xxIAcsgzucd8g0d7biJLV7Z+bNkUFBBzvnkyUdfbHu6XB3y+EXbru09OA0p4VpULiVaim2xhbDVI
b5E5N2Pm6N6NxEgiYYFgkC3BC4j9bbPs21Re82Ln2+HHusIBLXWd3c6qoza4h629Pfm1nKYZHU2z
fHer8VljEzfdO+5WAVsQ58TnrghB4JZzgCBjHpau/2G/YatelHSz9WjU+MFJZpTnj4E+nyfZH3zp
S/7KPwahYNF3OjVGJ4dZXaEfA8PGYTrd4ibHdcsYcN2DjMXGvabpJ8WgyFFxq/pB85udE+/GRZml
DUaOqU9Gyj+HK6nwfB7aB/PTkG7Iqm5cR9LDtavPjDDmDV7/uJUotO97iZ/go2mCtcM1XdcwSGuN
seQq5H5ujp26ibQOcHzcW2uwXj6YMf3USImz0Z1jMFXylkQRrcB49Ffsr3Fz6vjyxgLFmHH2DiXo
07g3+BvlSUf1SRy7JYoqic8OB6jHt29F0sUWrbxpWdO3jGu2jAFLqcwXel/M97OISW6DVEQdwPnh
F4iREVDzIY6AovbKCUl1hAN4hMSXvNSiVB+97Q0su0syPKKQvgC58ig3tZXG3z9A91PplJaWwGzt
rnVQNDQDU0SR1xlzdm715O14z1uq7XFngeGWF7iVvydeMg97DhW8aXLJtQbJY6/BdcKEz9dlrHh6
N+uPGKKHXkXRd4c4eFw5Qc3yQbsauUaudvKZUz18JGAKHMy9GtXigrSgoQL67rnsewhkTL2RSyBn
xHsJBqp7K0WnjXxeusxAoJOqXY5AvVC4MQmRAdzbnBThzbgyHLtVQkf7MBpuBDdSkaYUNg+cyNgr
gSeSndgdCLpKpt5aDbU8rfsaNHV5vKs8CsydlsXZzkXFZulCFkJ9NO+nS77Qsl7NydPMI6j/goA/
2KVhk1fzUy4bQn8NcUCSLPHEgJ6NZ5/1RDTA8txsjUEK2gFEja8LvN13Jgv9kSffdjyg9gx5FuoX
9Je5nLrH7cY/7ebMZPVc0SIiz7ITfugmM7k9BytRYmqiTlVMgEPdbR4WkDrJuHFvdRZgw8D4Co6o
InLhEWweTAAMisB43FoE/wCRggh8dfDt7osuME0rvEr9IJmXjbM7MbZYtwCGnQ+htHIkeWSQjnHv
+BPM2uyXwSrULp5q5hqWPs172hjOK9O69vNKako8wHVip4iJD9MY0Gia/Ef9yseXdL0MRpj+NlB2
F9F2K09qickUx7FsDuurR8ov3g7AH6+FPxC63Qhoe0bmXQKEDsLjgs1mruFVQFfO34OVLNIgTUdh
uUMlV9n2IE2BMJTNVnffT8BtyB1twj4QYm2SgLZcqH3eyiV2v5iP73dgJxTimV4vJaV4VITSRoxw
J+sQwZIcIx5FKg8azK8jpKVKto8H9X6eu7u70hcDMkIQ4pzbDM4CV86+IIu6+yNPUQTY0duEy04/
fYn5yOyRL+x4T0LemTP6H0Hs6FENITxKQHVfpM8FzhYC7fafnBOs67/kqXc29THIw2EtZi75/lf0
O1LJIWcI+omiG2eQJK5TKW4p4Ux9SQy0DwOd5gSjuWuVn2jIfFZSb8P0Cl0L99ewG9KfMej/pT2+
egl2hRL1Mqzno+QdfU2oeInvT05URHDpCLYJEdedA4A0pq84L+uyTDl41h16R8xkkniMBGW73u5R
p4kb8O5pEH1Sg7XUF9Xcd7iIB4LfJGepPsDb9l7iidu23JJc8/jgo5YIDxtQLVXWjXXpr97K6r+U
hGje+3VKlYL4JxhYrWHribz5VzQoFTEliCcqN5749UvVAcLMlqpWho4uIRvEHqfSTLmV4sMr7HsF
jc/Xihm6wCEJaxb3wJ2r2ghs7jv6oGH4ysaFOJkOtC8VdiE2rU8xVExI9SojSu2nbJlpwHcUb/+7
0+at2zslw7+iZntZMk8/0MNInf2UCIFi634BiP2j6K5Od2+HniJoKWFw7cA63D5MLX1NsRbbv3P2
9u+IJxAWM9ohp12XxN5XLhHo6THAFHcWcBHP/MBfSvBkUzQcxIVrW5ZR+vHcT61ItnHpE0Giw287
POtfzKsgmZXn0OJoXdVVPSIJUJGCwxaXv6E5yFYZLunD5uFxJbCDIQxMwzTLJ2x8ssBtaC8EMJS/
jMuMkjbOtPf96k7hOmlDviC3laAMf4WE2XFINZqMRLsC0YLU07uKZp3Rj4FU9+k0QQG/kYfhznUe
LuHYzoB/pHs8i39wvDP/C89aPFJD5k7pFpNg8jTKBMMapWC5uTn2Hg3sjIUzNZMF+UqmcX90j12n
BF/6/Wg3OHewhKVkHZ8UzKI3wmIprFhAmiQQkLEw0fWlHBul4Xg7VA4nVoCQylf1UoVH1QeK0z1+
SM55xlcmndHS4wdHg5dgCVBI3+tArHsqK950iVg6tiB0OJfa08oQo+2jEzmgyQwaOgdnuJVPkIyc
Igs1V3+c7p07damcoGWwRvdbwSGS8CZT8B12fU2Gl+bICMtilQwXgQwCfClHmVrgFe6n9cZJWBdR
YOk6VkutPneW5f0v+UzX2QCubQ/OO0KyqFLvs98TN/b+hNCv/ohznn7Y+CkF1Xp8awzGEzjPOJff
1AM8T8fyBE95Fpldt95GQztzr51SimVT+Gt06je26m5nljHex8qFzSuw1zhBKdQ92wbUufmqWdEB
TATLLaPGR+LoxPmYskFVvOd5LrIiP/lCwqY+z7mMMSAmXQt6PuuEXGdwTsl2445uMTTl3PV8roji
FlXcWjhvrK5oQnh2sdX+pHRfD5IQFiwORAfirfHGetUKCFkSRMVPNi88SBSNTyz24DOKblAfQJmU
fj5Vkl2cxwyxC8on6/mD6s3a015SWhZqtXMQLtM7seDdxz03b5S0FjvG5tQ8LG/8Tbh5kSNBgxfT
wDor3kF5i9w1IdcxKiHi9SUFWugDj/PIPL2max2R+SMBXZgrcsBZFfY+/2bCDOQSUDSSnoCymQP7
YA1tUHK2gkMXlGcMBXCPGOwL3aMtCCxYPD3zMU/gl8+Q/ZfiGXQb53mHsBbyPgbHphMU/uFkRRW1
H/8DZ4lGCgyUR0G3yWQAmuDwUR+20Nv+WXlRabWJ6HbIwF3tpGfG+xLARaGaQ/uTYRyKQa1S8Nkd
fHKLXYHS+N31Hi34z8WsKqSlsvurEEuC+6+Nf4aUT31oZw4ZIFTc8AoZuVGN2IdczHXutWORKBkv
J9qDErnxbB4tkrARR/DtQsLEF6jJModvDoSQCb5+pLEL9c4pJjtcfkfSUJKaYP9E56ChAqqJc3Kn
ZagXNWyWwFeFU/6sQYCkcySuawiBrwqosSHuUVClU7vBaBZnYQoSmfMCas7CT93P/xLunDFKFDny
qhrF+ceDJkym2qBUex1GtqDYcrgRH1skHO10hWKJsbOXQx3fHqBJHbK7xXIKmmvwMYmbLe/DZ6oG
Hr6WEwDjz4Z09HyJuTlaZrLWHnF2gH04f5Ra9zuNqU6777fkyWZO67oCw8E9zpzODzDq16AWIDIu
HlJyu02Tm/zRHSlzfZJ0GUZ5HDSMzx/bXybe9AFBioniRGrtH5HKcInLKrdzFUfy10M7O5xhhmxR
qLIKxqfy/H5vekoaUAeVFdeFpwi2hjv204jQumcIIYcksM/5H5sZlf7gvhgphgPBcbWh8ptpMh7P
ul0Ulxh4w8IVgS2e3IgTsW7pny1wEzlkVbAWLQJdHgXxl9PGwK+xUZ+b+uVSZpB0EyNacxbGS31z
inY8Mi4jBumKiGlymATtDltf22fvkOileS8rp7q30shx1BkCAthf7JxM9LOI2aa8Mm5k7OubRQfS
S38RPoUiDotLH+c19slULZY8LvJp5/uXKiA6OkZnWwZJja6hyAKkNugyiO+EEMEDRg57mnsGbR1r
WBawW7+ts7Azu2uEYGXmDOv7oLqQbX6eXfXmsLqAq9x/Rl/nZsROM9Fo0efHhcSlEEJcuMnqbCyn
btrxe06VAl5A+BKYYZ77q8BeWx/Nx2pBHgCjWpQ8QOHsBhzJUEpUnt2hUgnZ91Csu+BvCYK25C0X
zDffrGPtuaqzQnu2D76wZUNNVxtmoPTLIg5qoy75UOU5YRsiRyVEjAqEtlh6RNxnyL8k/KcaCOfZ
CjcLLHx90iXrH05ddX/0VTIZAeuSZSng0BlaIQnwSs2690ibsFu+7QHEKqlotuQceOJCJjBbz/05
nmxj0QOSuzl9xuVkeb3KAaUTj8tCYQtlglACuGNy7SXPabEeQ7lH8Wo1TZ1vE6vpE++dKVWr6O68
A7SXM6Fh+rskLj7L5PupQCYkCqe7DIlPcVZu891q2xnMXGMiw6cb2X4zzQPzE/yE4nSFnC5ejh83
y0u6i5bgjGIrPz3f+2UzwZn5n6YBe5wp2wAX440VznDI1JwIUPdOz/tMCAeuiDgEjqtObkZpgpK7
7c5LVCG3EvvP/tpeZntaQwynz955FzhFXafYQupDLciF39GdgykNQQRhOPa6jXLCKi0q5qGVuYDO
tlW2WY53tZFH4diZ1ZR9oreNZw9evnGYKmfksWoZhCOMvQiBO3+zEogIXvBaoXqdYIb0GBxEeV0y
lvkwrgDIWtTxJlCF2yq3QU+OhYDkHHKLYC0ncir7tdIvjbsG//LT7iiQtGn25MMGj+8WZnffsWTv
y+N/oMGb4qdcjElGD1Jn2N3BfIyeZGxajRVreMr2wNMLBb7Sm6icj8/CxEHOElLpIGDHRBTbxZkN
Lyl7rIV7ubrD9bO/MIudaKBVEt9JGUzWwwEieLwCa33fXtlimJuKcbuuvfzFYBaOmN0EwA+Z3gf5
rAGuHZDLnEJ7hJqKkke/wgq+jaqFhHH637xnbvRKHxLJMnQ9yV982PZiDVKFNlAOpeidVlWt7kc8
/T+8ThwL2rrCkRdkPCqVS6cWuzG9mfPDjCIEALA6s+x07DsPeDOYJSIjsLdTR1tj5Co5sab2N9uf
o6HbGa3ZNMBR4Xyk2FwhDnLhZ/f5IgEt9SS9ylYPzDFMAKIqtvAOiTG3238VpGNR16qFeaT+XUNr
wM48DV4hja0I33T0qJBIhAYuQ9y+0riz4gAsvQ1niL5fl+7i7kY9KR3vr6FsnHojpVT4RaVq/+GN
oy2EGiEqnCAEza5wqTHMrH1zC08YWoo4Db+UcxiNdsbRKy3dP071b2fxf62ZtjGqPKxZ0mhwdnPn
Zt7vCKo+RcLi4iPfHgd7xlNjixEAkrGOB+1jPRTAAUaunD+SwklWr7hYII6QAzjWMBVWYQCWkG2a
iWeyXaFRCW85zHiY935A3oYcot9dQRWuLQ1+w6QFAwpzsfhWkyuozN7UTt1tWj0OZMROqgt2Y1y/
5dKfDWoQ/WdBXu3ELddRi/UdOFWAOV//Hfm0n29EPPHK4bM+3dBZ1NLlUIZ475pNZcHv5dp67SgQ
DBCWHOTAlupYkgldaipu8ZH2ty1vxTsNAmYPdK7S6vWk2VnKvhR46Fhk1DcJyBu2en05nOnjLEdZ
6o/42i5XJgFBM2vNHSYAHVyJnW3uVmqtrp+rIFqyrESieIukfEMlT8hg14NgpJ99ycGd4yfjboPN
CgixZs78cVlmaJLcRHgJT3+w4ckJfWtkGZuPDb2vVMupB4TzVgpYydnwRTtB3JIgN9rngKYtjGIq
5Z/HIFGApP6dpO+mEnr/AOIh8/iPQagnETi5j28VTyv5z1FsxkOxbYarr8GEkEmg06ch3tk2ICjA
ZmWgOdWuYM7wK8/FFpyZdl8TAtCg2m0V5I92a5hdDEz1m2cwD+KsWgxHSKB2fVbUjsukAQJow3vh
DspBUEGAf4a6FiOf6/Tq64G5Mekq7XSOQd6LjbIgxp4fs/cWabTiibR2QQbaKqcxURimY7buN6De
DFiXYbxcwb8T52XLJN8CDeWCTwWinWn1uckTwkqyQV1V0nqNcYzKn6H2fCmkQBauf1BhDxdUdDJD
6N2W9a5SU0nrlbmVKROwrzdqGofUXdowEWINnO7jgsYVRRGFNa/fz45II3Jz1e0yH1Z9pI5Kamle
O5nlCyc9a95IsABhu3yEfhOIOnIVvU88wiDK9N+5A+e0kkRApavjkhBQQVgD9THWHNLGjR5dq+pQ
c9ZeAqrrOgDlsTxgIaOusR8YWzawahGSMH3KuF+xVs9GawTBcVV7cc9tQet/Zb5dEeIW6jx3+lwR
2Jr1XzP7Dez3+4A8y/Rz2mWJtkktomIiDCGnB8FpKKFvFvg7GrOr/KuCda15JG96CBQHV4vsOdij
mt5en10Uk6scORZLwHg+A5uurK8F0PAp9VJ4KepXW+CBa1V6ELPw3zPmFXMLSOcTGPySoeEbAlmK
Bri5KJyIJgIUzO5VxUC8ZuhzDtdpBHC4rfl/XJ+i1FEqMbMECgsVaCU5QQUdUf1mzBwMHo4kqjyB
46F8+27R8ZIYdIeJvcuNoEbjUQLDCaOMia/vaI8sRiSnNkKYya0kQAjkYQFaTwbAcKxv+ndrogq3
Qh9bUtZ/HB6X84mqF99OMxZrcNGbyiwhBwk7RQtvaH+Nd+MG7hcQ/zQnqrfBadE7l3BDiq/wTUju
TEXPqBFYR96oT6uveFqrD2jPjHr5BaJvuIFVviFYIRPoibIa8TyDaAeAsQI9EIN5I6+JRPbVrIGo
3MOYlbO59DcfouaPYNJI0dDVPKoXawmeaL9tKOf8ENb+ilulsIacD76AZRQtlR5kl6c82HXnwX+H
DFO9A4d4j/D1eH3VNwd4kN1pzViEzVPQmmyENfCxG3FeohBpNAk+NR8bRqL1s+ph20qF3d9Grthl
Iy9+PZP0B4fb3I0+kcsIl0fCenCmkJ7OHwWopuOpMoQe29E8Y+ISImoiJ1khC32mEzXfEU6Tfruy
+Ia713xzfCa5A8lwY47AxBOLXMzCmCa2YnVY55j9aMA+cH4RWNMvYnNKji3mryD7VZbz9UMMD4a7
t6eFQkIWmXNgzRQpsDPApz2SSLoK3JRJrskj7VODnRcEwvZphw3BFiuvsWiE+f7wcySitX/Gq58K
BmgH5UC65j+q6k45MVKpXd78fyPFIuwURoASWH0gmteUo69N1wWBKcFS1/6B6Io84EYEQsMhRA/B
IwI0mpPpizykG8VfSZu78molygw59Urv6Y447sJFz49oodknu9HmB4mxG5xXtu1V4Lvv3WffGwyw
un9SzJhADsLmovzgW8Ej2Tw5NTVrBp45NCbGRfFl2fd+U+/rPO6GAR8SShgkqBZ1JhPOEmEIIjd0
jrxr7c+7/ZrpzwMDFcSl4lnXUmE+CCjTAg+AxNylJwNUhjAWwJ9VcHYtNKdMrnExBAjq+wbLegWT
q21oDf1KlrPB1K7I9u6LfB+HLcLO902xJRifwV9kVJ3eNG4R4hFB6DIpv6TFmhMMaOeC+IuYS1Yd
aBBiNQABLqP5Cv3q/6AHZvtszPiApfU2YyezYO7rCwkNtK2/SYJlrq9HfD8/FZRKPrfUMecfkMsx
A1qWsLS5aFkyxd6UpZDCDomGRfadcCp1hOiqbJQHJlHrPDKc0wGIHZgDajNTn/yDLqHZ7t/W9Osq
awkqBRU023XwyKjp6AV43nAQAaAaU4Zo1vPx7uQd1Z/bfUwVY84zoosUcfILMiQ9IQ5NuLXMLzjj
/xI+VTVvow9FLfGn0yU5pH0OS6zLKUr2e2HMhvMi6xFSOsi8ysG1vNcioiTZGuBv6+OHJujlK2oR
Vq5fInF2Pm08TJy0YWuV7OjouxsD0SWb49GLCpGoHZCzVoZYY/1ChgjBkRCKxUC/xWH8d5cvXhHZ
EGaSI4HWIbGNn4HOhqq7Or/RDiXvmUNOxZinTsrlvaMS9/udALACfzeoq8+sTFTJ9nly5QQQL0Rd
pX9x4WIC+bU3vW1DpXWrk/SMJDirrJzYhAVRdQVjwqDm6U8SpQqY2V3c1ctwpT703AnQvuT7ArEp
/UqS8EXnaDoq1CknqW3zXCbP09aZUA6gvkIhg7xjV0EV0KhJvkiYe0WEpIaPNi2Wyj0Kx3h37X5P
4HAWlHXgRtvKPds5HPZdPdGVf2+nxe491DYFW9FLn8iivrgBX/RsurnfvQk8vAJS7XjILt/611u0
2ITKlZHEM3k8+EkF33sd+p1X+XB8dAIDyhZtW2xlVU2rC5IABEqfuJc0KPXl+AHH/lb8foTDo5nz
SP8amLX8zCT4Bfcalwq9nYdgVfCYqDI1zsckVns+n7NSuUteEe99ejONYdIP3XhJp9uda1OvYfj/
Who+6k2TZ4FTR8KMkLOsNDxG7J3HXMupRebyy1LobLBfjduuz0ptd1+8lG/ar5O0jLCOGml3kBr6
C63f40Hw3OH61McFQTwN5+bMRn/KQGh+IA8Bx38b2ujVP4/JYUQkw4amwYXS0HbnUDcQ5ejNdGZW
eH22bGHRmgBHdkF/Q2GYsRS29L19l7jc1qiTA9OIgp889Pc71GkGTiuJ0RUPd8OoC4Dqsg28nhwH
mLFLN2bggBEA6bnpTu/nYWR8QjDoDqFVwnpc2LNbVjzfp1UYbFlJHEk1Q9c+AJ8cwukeJXzkcc9q
Q7znPnUWHXz57A06pR9FLd53iGbT59s1g+fZHyI3ZWOHIH50d9agt5JZ196x90z5O21Y9KpWzOcO
EIajYWdeDrlKx1EO7XfYv/yO28pskoNJ/f8jFxFN8fLD0tpBg3kzER4yiyfvXnaln28Ib3WPfBbo
DbjN4GLVkGuSg3coVzwmZ1a5RG3IVzKAtZNqWLIIctI8fzGRMs9q2yh4H4Kk4/Yvqb8m2noa/EBF
fQ0IydNM3RZwK04Uavy3xxQz07oyptavPymcrmDnY5U+YwKk1H34qJhcFY41RwC3vIDRlu4pNDVh
taJyGMnxejyR4UbUrfI5gWwwbQ+ufIL62/AqwSEXtfpryKCDAXHJRz9SO+6LqorBNTHmNtKTUxen
cY32HIpVkMt8d99rffF/pOIc1PCx/A/QXCtAN35ihuVRc5+TDXzBdpaN323IWs5iosv1ytyZl/9Y
h1arL9CFXMOjKBlfagEMI1cdPvASGCK2B7P7EBRmyvumVMBybEiHd0w1Bcm+0VnWlChhCZNY4Oom
6YxMHCdqN6i2kRAHNbRSY6uRy8AnE9gdFPCfQPbwIHX+H6jwXIr29DSO52tosNPX1+pEgC9SJrU4
dsOSwEfKN5T6ZTCEcUO2pwrRaCBadzed82GlgKGlW8+P9qoXfLOJmYCiFBTgiBVGSRDDKoAxlEz/
LlI3l0q4VuqjR8GyzQKDDAOHNNbfsHrCjukI1niVIcPVhm8ktxocB+twZ/AwezSM/f3gu3sRL5ML
/Dk0W0T/U7cvMJ5RRVgw57rQ8SdQONZ0X8gSo4OdF62se+W9dGSXCbkXVYz3+OpdjZy4Hbb1LJhM
F0e7vTB35UqPsujUxz8vLxSOPQrzJHiDp9plGk9Uk15ugHceWcAPd4+gxlm5nJxGnCUT6CVv5FlX
DHzmlPB9PWhvNfnmIGMSFbvH+ND5cu39SLjQ8pUh26fOlrfCa9b8mnuKpvT375W6M+9BtzAbywhy
xD2u8lD0Y5nxoAWyLld5qhg98iS9mxM13tI/GIgpoqgTYg0PYwoZlBjd1oHBdXGL0xtL0tlmQ2WT
E6Dd8huoXQNtP44SdUuQ0T25hoNa+g711HudDoJtVxBarMme71IGorUVuqAj2aITO0boPJJyg9me
WuZVDqJ1vBYM605jdYA6pBOdlG5aG1Kf6F+zhwqXuoktwpOZEcahdFZf7nQ+lQdCKChvtp75MiCF
b+4voaAS087/yZk8tzY8EdB/RX0UF9cg34O6IVb4jtTTAcgMJLzxn7uE8ZkE3pe4G4DriPvh0wvd
G9KrsGUUJhksZd2Mxf+d+aF1YowZRVQNCCLkTLCjlLLuVNdZNB3M3rm10KsOS07i6kwEpI/1VWxI
ojHV+pNF4GALplKfzH6p90p8p2S+uQ96RXuqEcsWpu547biRrs4fWQxMt/aiQhcjWtfjpVyAhuzr
r1JQqUDBC5yu5MQQ9N335flxczhwqxrI8G5I+zWbs5vdWZbrw+edUS/0Ae3n4MErfHtFFfAGGFSc
/Op2WPRiSzzPY0GPxKBuYmT0k7UNOzTXYCyBUfQ8coD7fXOLOb83NBo/5YkgfZiF0WVPtVcklMN+
V+MQZ1NjHaWMHSbPe7qm+mNfhw8ucGTU4lvGCBvaWykPo/7WuLNrd7rOkxVcI5mqE7xprgl1yTw1
c8C9Wd2jeQ+2keabrlc41vNicvzpd1iukFdDZAqUQhqwOF/S6KNjbjUODnwz/Y4zaNp+I8853zwE
kafSr0n96/mumurexDm9lrYKE41NQ7RdS0vvrtMNG7MXL26hSZCiAsaHk0KIIwr899+GIi6XGIXS
ReBRKNkHisGq9+0iURdH0eL1VMz7V/bjZugJuTwWvpJ+UqQf7j4BEtC7sXCAkhSW+Iq0Sltdjwig
pGqXLnPaFELDJqTg8X5X65svDezrX+UMZ5AtyFqx8ChLU1jA0ewXufZ7L18InEiEOHZm1IRFGM48
JJvEzsxSAW3DMBoqdulP7onElVhm0tDiE+qW6e7p64YsBQnIyGoDVDHO6mxV3JBF19DlchRCDk9T
3LzPuYDuJGo6WKkU2vmuur2H8lJ79V6IL9PdmpsMVAsUdfFfhJMC5CT2kJ5/UDeG4gP0iU2g/SuB
oL4vjuJsAvYVP8BcSz6kH1wL9MleDIxQP/3xLsManLBywENFhjqFt7tcSNiuOG5Z8mqytNbC6NsW
u1t7xk6YnIX4+GQC7CyyrwbZfOtTv75ApHaIWDd7dkdme+1UW8tn/IFFAg+q3kIAFQBeJYrQrqqC
dH4orqH7gMKLUHUeaEDBMchRpIQTZrCvK9UZbSk+M8K8otTl7YoIGCILgmYGtsRjk6WGWzvgHQqz
G++FbLkwd6qbItCnC/zwykLH7wlW5/zozF7nQ/DsKOpI6ztIuBwA7KoAR0kTYhhDFGfEfr2UcD67
04+SUvGnJP/dS9B2r37Sm5Xjof9LYVB/bFXGNok6RYIL2jfPudk6pwgCoDL2O1tW6sdY34LP/DwP
5N3c1i34VHZC+0aZINVCOcVUoY64ZkO8Vf4TXWkcB3nC9oGY6Sq+nGE8dODuQWygJWH+sshU2Rjy
uLec9Ju/UpW16HxTd/Hy9H8L+5eckbOSZEiPRbFokdKszup63fxADAykdjGdiWKTS5RY3Qv0i8zi
2NrsO/fH2UT7Tch1oVS+rmQbGjJqSEFYOVaxzS8lugFNb2t/4Ixw+OBwjKCkLbGo7w6sf7xVkwSK
DPDXLBZjkRiv96E60tpfc6cQcO/9IsjvVq2ffxQ1sPOe2zQyG2LmcWEa2chGpB61mJcvvq6q4pXn
PmdXog1ENnnGzzFpdbUj7YcwAEXabDzz4rhP5AmGEL4dNb7TFNXPUixJXH2zN6MwuI6pDjRZD0Cr
jqiFwmcjanuv4lxq0ejz06XHCJoy9DHovCHdGU/m5SvnoB69gEadpwg3LPwLJoG+t6XDbEfhwu2z
cFI7S5/jCUbYADp1+ScZbXnZYiyh6Py7CyiG/G7pF7rOpY5N/8g28IPut4QCf8t2c4IjMX7C1CJ6
TNj8zjjzJ6I2tV0OOMjz0Ckab7U0c0UPAuKWkwsi1O7brFgierOkg4QMhj6c0COwhIkcoJNuP6WD
R+LCH+Gtr6aRqA0/wDntGwTLz1kWD0c3xHWU5urj6oUgcB9byW+9Tpv7WIJ6wpm5SX4l48JU8J3T
SRh+jA8K3YCCYgrFAZ8JTVvvYaADSgCT3bzGkktEEgFtRwB2/VhwMSDiqJwR7xxfa+qpOZh3z3Ig
u6/ERSoFZNUgNvcovmT86aX7vb3swj4aBDFgW4AWgENnyd1L7APbkWigdghBRp0Dutul44BOUrrA
K3cPYChSAidRn64sDQLYehNUSyGzgflNwjJf6FdwCr8WNadxDogtslAm3AlOKqLYlqs3/tibZ9hP
CVzmc+DOcgmS1vyY2zbCAp4o0Epiz0ubPEfJX8nGGaotXAG8YtL78xodIfqBKDWVvs711FzDjyf4
cxV3u2GMA0dAdG2+hHIV+tkiTR//EruGuhDjIL2i7XgE4jOk9bLGKnD2Kfl2OIFJzIPnplj2cyEO
btVXZCHnwyjlSpNMM05HUWA4OBYPSaBiPO28b+RFYp+Eu7gtdYuX3BXz77LR+P9IosM1WqP121kv
4A1G1Jqv2GITolbyZuPWTVTjBIt53a/RLBmZgv4Xz2vFY7mV87qcAUUIZpWpka1T0iqjLFf6s9SF
J7vez4gw3D2OlhytkBMNEyGtHtvsPjOxljd34kF91D835Nj1YUK5sNASXoR+bh8122btDrNNZgIr
W/x4BORTCRaDsxeR/mPfsXez8xJGk7+vxDcwwpS9JbkA9vpWY4z20MggyaFEolBX2ceNH1HUlMd0
+/uBhwoiBY9FS2u1RGJBqCxtByCr9faKstawV08a1u41LYG6rNmbKGARVosoTpPx5EbVNLugOshi
cEy2JHLGDot7r9aLRRZ+3ENMBryHRae1pTpcw3GjrOzbmC2t4xJaFgOS6c0xNaAxb1HuY5VoGWU+
qPuc4klL6yOYOP89CS1y8RDzIYrWlB9ZY085iUf2beuVpA6ojvF36H2vXLByE0z2y0B+2WLSKq/h
kXgB+tmuXQOqiliPqgl1bgjEAfr5tgtiB6pSqpn/31hGw6bl/cwe+xBSznQvOW0UQNqoptB20sOj
0amUrwcs4psUt/radeEdms1MNSTMuNHlI5cVVMxOGj5ChTpp1TgwrlI6IwcFXV9HJNKjDUIFbJ79
sh07qrVIhQQi8Z95os2IbmWHkZVR8aBnv25l7KTXOPBcNIRztMbDkQmEGFQCk0JvcMZOGfe91/bt
cQY11twXWv+bSiXnUBrGBcGU83GM9Si3rU29K8WmI3n6Z6SkdlsLVzvhEI7Efa6MNLBTy1LNis+z
FKl3xLV4+eadZbGAth2VG5ofFqFL9jD6hOEbfKb7QGnOmHR1feB8KFxH1/JTh88UQM95rsYKmgP0
mqQHPuzH+X+xG4OvFSs4bfWxYc40bro2mRSiuwTi8W0DDzxgeuIyTfzR+lSYdzxKqDfPhWRxWh+m
apTDz+kQDPB4Ow0Vighuf/TYdR0x/t4ISPhwZohKMfsA73LHMqrCOw+Tj5iA4hHldjzuJ9cDFWL6
JZSs6erEOFGZXPtc7yIvH0CaQEJH5o+TxhfTuXnDvZlWmQzusTU2qqToOjF+TXVcKe3zocR5nkrx
kA3Qwg+ACUZ8tLwtA806wfMmNBkoKrDKPP+dX9AGSOOm/PJS++4HP+sq4Ehqv9xKW/sroMFdnIKS
+fJlPaKF91hznYNhmJmTHL/NM1ueRYUJsP6omnOD2md+PsjImXz1k1Hp4fX5RlUCB+O0Mw20luVi
ZNJo2zkidOs2SsbTCS81VI6qn5o03iKCzLKimy0ZHQxsGI9yU/WewHz9tz8WAnVxLNj0xgDuRHPJ
5fbWQ28aszRYH81epxTxusQoJIqejMUcRWXrJZu+z2CFpW6nE9DCJ0LMIMRvP5NFoAAo2rgsHnRu
8eizgY1RUgCxpSJxenNF1Tt+WZFsT2gS1mTdRfJsnSMEyWKg6+sdmKO3C4/Gz5wR4DjZ5jHRqFpW
cgJN0GL2XX2vSnZC4dl654hFl2BXDKyvOlkJeZqdhYAf6UQNkhyvroKE3hW2q+FMfks70UCXeu16
Tl8VKBHxoSrWMKHZK5gZTOj3M+yToWJTODRf5F8CjJ94O3aiGbA2Hw8jG1pRLdJA+rpR2cYbPd1i
40mvUgu0d6WuPJsB+eXMLhX1LuUjthTtjm27Egpjvu2if8tXsXCJmQQ44d7YTEcZVQ7KPHfEjauJ
S9WWJdDGnv5j8usU7NKrHOhELCLMswQXJWc/c2xvtXjuhLxqDjPNCHURdFOnGEj5Sear+zldbKXI
JDrH8Ta4dyun9YdjzOjAl7VXYT0N3FVJDVfd8sevX8wHwsIiq3AcrrJI68CUP2aupMNnnrcxJoTn
tnvsqIcPdGQUJn/fZec6XX4NoK/2R5k8ghMQUbYsaxQXD44y9QiykrFf6fTyrKEOiNBQiYUOwdJo
zmzDpwMG4gh++oo9GcOdBnUyqpqQuwN2adauV+cyaYZ1KL8i1WKn6UdHdFXwoepZA5b2x52lUTo8
Gv3Ze1GwAdTvLh1f07g+a1vgUc0l4Xf48s4/NYAw6OSkttEGT06wb35WhoR6pBAUKBpKsr8rTMFZ
rcdY0bEHn/udY+7F0szgbS6UGZEK7JtDssTbTy5qGvV1Cao8k8j6F1se9aB+7Yzzer5weybCj+6d
1MNhNlVDFBvjMPkQCWfU4Dya87ZA7I/jKJ/AMu2DxtQVQMUNw/2FwvSLvQR5uNovk74kf7VQZxYR
+/HjOTxeKVl/87CKbW3zaxHKXjINtfMnzhJB5sGAEWiBA0+LGTjmhMR8K/otgvUjP/TQeCCw6xmF
rjO0vWAJIMqdgBot3AGLtQFNhxESkYtZoeCe+jrlmnmLY0lKd6FqOxT/NJuuoimrzK/8PzIl0gAF
Fa7p4STGkaxtDMZ40chSlIq/sWfuh3dgzDUsodicMYEM+O4FP+zSOVdqYRZfQ7nSDH2dPOz1dqiX
iX4PY47HRi5uq+Tu20mnpfPwDC110iY6eYqjyYmOlSBrx3NkHNuXSDDAWcskqw7ctU+6lV4FXAmE
RKlR/Fz6alWR0lIohC4nSvVf7Q/vSaBHxGRn9ohdDbkDivjs/AObRoenUJWrcJKriQp6gows/rry
/oUyGwn2ErmE4/2yZyr9V1NeUkRbMP2EG2zSYds2gh+iUvVY/nYiI1Fyj7/45c2U77Lh4URHHgoW
xQGiAaCaUtWo56wdfuZ3sSEhEfgypBp1QtYocJ1CZGx4YUGM7fMY+TG82mBMqhBjQXshZAGAkhmG
zUXHtD9wA5/FroAhGkdrdmyDVXaaVsKMsGUEJq0+xy4qXdcMOH553Va1oPpprG6zP4i4hv5C5jqS
B15IXfP4ADVd2nQiyGgsqcbfTrAW6sCw+IoyuG5AmKjfNE+QLTPPELwRNY6vnrLK86oerqlElFOg
RwOMeoohP+l8+8AzKW9GVxW4/ZLEnTiC8dU7x5D/D1F6eBfzzfA1PvdpfjPfdSlnDKPt8BKs1P+t
rXhqC/hKrbO5ms55AOyd1cp7V5S4WblGKsClbp8K7UGVaFfBTVIEMMgi1uKdquLt94QrHhLSlyAh
S3AzQjqGTbo64gpfY/yC2soSvKAyelprzGNuVcwqs+lofiNZ5uKCZ9Y5XLyB4XbQcV9gLZHHavUb
1iyOtjthliB6GjYa06eM6rNqfD3uIM/+fpDmmVr3KuSTJ6jR6PFyhwrpxdsxEQwb+XtVXiIZ7hP8
a/T42ixIEBYVphqdVb6pZT95ovtf8o0/8SMenjTBUiGBD0+4+ns03eajz/FNqFkqPvR40crgGg1/
F0xUJHy01HbuXRT4Zl9y9QX5knk+hAUWny+ZVvQRZiVjIyLv1jFwU8dydwfsEbYQv5HQVkdvk2/I
zinOweVT0VbYc8dpYotyvZrKAXclRcLCu8K5Zh0+q7FmvtJPLrMtWEfPlzNkXjU+7jljFLUvGTp2
Wr+DrHdhGnFrZVS9iPvwrAwk03c9S6daYTn1TOFegzGXdEovh1iQo68IYv8t1sr8nj5Zi+hqFQyG
l6P8UvxM5gt83UR4Y6zhm7jorjnwvaFtDKjM70ATLPIW7fsyOsB39qa4i0wk8uaFfpBqPyPYTwUn
SYiyvJ4M7/E5v0mhPu24UdI/tNDu6SudFvCPr0SrlY29DRY6X2SRc9uW+gmg0VRPQgiy0es57R77
2uSYBDF0gXndHZojz+KTfbsHg0GLxu7ALZLBS1av++Ph+gnoy5RbJkV+8lcHHDZIqKi87HO+uE4Z
fEa3QrHzzu+2ogUWz4+8/gNWrYx7ff0/z0zMgnNzDnTb7hFKuHZpdD1FFv0pGJTobxxVtURzo+wx
+wtxs6/awb6yjMXfc/xufMLue9A20vdvj1lBPM5lJIn9FzHq3yTVUtHhh9Xj+cafcr9NAjEEWq8Q
Fv/9IzMDG+F4BP5QK4hAdkporDMf4v7XuzPnkGc7pbtz7iXkuHprnFVxnki6vsQUyb0jID0VKZLl
US4r1cbzvjbwGJz1IDouhOzFO1GUHE3n5/e0nil36Mbu1cfSxZAIYYR804hs1SiEDikCmROGqXJv
KfsUPOS/cd8oqGTs56nXAP2osFuhcL4/cAcOsj6Smcn3SUcgvP6xMexavy7A28bL5+d4P+nIsPVz
4aBowtFDtqS4GaVpzITiiUbsrVYaox2+m0eH6EDWUDK+rcaSiJVhJIfH6xEfqIEA71mwxiKx646y
cH65oenZ32f12c1tu1Icx3HRyIu6Nfj7I2gpg7H6j3Ham1DpJGnyNwHkVBdDUnMzSKLgtQqCt70z
IJ4YnZM7qtMAGAe9MQr8MHC355V1sFZpJZux0BIE7yCSgrQ8Ck+Vm0zDCTn1OxuzlWSI3auqWXdv
2PqlaqcBCpwcyyc6wzwP8kbKS65DrDGAi+u0VttP1MZRGeYKoApQLGhESgZkxVdiayED6vllvhrP
0fcjntHVFBz+okjI9lNyQccFYRXwkdii5kszasraub1Pk+DkiW30raqZDl76kWddPsyFXxhWTNJ8
y5R8bAuxvGqSpQbZrI7jgoSjwdGg+gkyU6X60BG6Q7K/CkiQWM5DuQ99WZlsITyM/c3NOJ5cLrfY
Qty7BCTu4C4T5GZ8FN3QN/rwYlrWRDaWFekgVtRDCuQx7Dk1powPEdk+IxUsWxa1kDgqq4xcyaYd
B2R8k9fSXzPiafgDPeQHqxYrTiqIDO84ulKKQHSAiwAL9w9d5C+0lqdeNxWmCosV9ou3fAhOPfe9
UdY+uEr1VLtp2YL3M7k21njfIj4J2T/hoVGqemSH0WKstcHvoI2LTDBauCMA5zoVyfukmyI0bPFp
Ym5IAO3tetXGB/URinAPATNY6kb8TB1GXFKPpt5kaQS0kvTgmvBecn4+Zp38tb5Wd3UUF7eZmLA5
z5JJz7TTIN4UQxGi/hJDMb4XtLDJ8RWzdql+8t3bMAy2Snzcclu2jSMhKS1d8MpQvVtaSol8mjB7
hVh7wut7RrzSiOtYYUhQIl7lG58lG3JjgpfMyj4SQdQayw/QxmyxnBn0sN9nsnCRUZ4Ar85+Joem
/sJAUnEDQ0fxhStbXZ5/xaxgrfRL1jM9cEjdmZEUIfTtPOdGKbTIcxr0Z9Exw1pBGcw0wwT93I/d
a2g9Zi+VaKMZEP2EJ8mTgmBl0q6RbFtP+/o80AWoi/cKzo8CSc30ZX7LSq+YQj0NhnusXey520dT
OJl2n6a5wCQJErof4i/1ovghOYmmifCNEUUrpRSo9dLBhFMul2C90RtWa6EbIpLE777CjcJCnQ/n
HAjy/xKN+mTwyCKtdmdDZ5zpp2IWMLlPTFG3xmaPfCQ0q/TQnaxn8+y8WZ1jyWXEZGSCjS0Vnkrh
yOSqRkIEoZgCj03v7rCusyjX4r3o8gTFQiiYccI5krXEA0zvP2FzQlOw2CY22xL32TUlmcXcLZXQ
mLdhefQgMa2mQuYFmM+JAQTk2lDVT7AzmT3Xhs1t4lO4SKReel7gfeOj1I+wszlRAZVxbYTM33Pq
ISBBsuGUOQWn9mKHMmgoCA66UDgt0xi64moh9ynIJCRyZ/nT9tBKIejDecJ6wmL0CecEotY+/xPg
3OgO1RFpNZUigMs2QbZ8bi9k+pApeFzb7eqVDa5YkLf/an62SuSRw7MAeuP5ZWn2ladRNCps73gz
3hoCb4mjT0TMXpq6w8gPfw0EZc68jgqGhNmRq6YvgsMPUDyiYFr2u5XOdQC6D47P2FtcWrSMbJd7
90hyV2c/9a89MSLnEEglZtRm1RyLASJUGc5/XKszBsC+xA687bT2db1jvCHIT83pwkRi9ctp1aFD
zRu/2vF8ZXJTMWMT0XroRVftw+clQRDuE+YzziGE7Kwat5Gegz1jx76LPom4j38JcWBzClVEoICn
9imh3VvtHfnqiCOyTf9SA5u3rkEaePCLjTD+QmlcipMbimU/tHCMEaOAh53tQHhMSsDwoXxbCKMW
xaVWMB5UzbWD6HykQKT21elkr08IzfWYhDWwQJA1fFyoSJ/4P6DehscQj1AFPi3wgfdsX++uZwQY
MtjZHMrVQTF20452stQOIxyrPlnEXcehr0JWOeju3CyPuw0EoINqCsOny7+FBSHul5bu0v8DRnOA
mC77dp2S6xwG08N9FZgBuE2HTWxpyJWKJuPd68HRdCYdJJJIjHcHSVccfh8e3RCgZOCgZsIwRR4v
sBUFxHwPamgUhaEpJ4K3WgBnIVACk5y8HlXlCNNmEZSEnTkjjK6TAf1i/lCo9v9XcrQFiPE53gOF
TV9qDNUqLJkK0q6TibtX8D4J2m4BTrI86Jz7TOZuWq5srwl4I1li/tRcSqQ3iUKHtso/1F+LMm/D
SU0Tc/lB0cPPGvsr6Kg6Hin5oDWzBZZ/DH9PE3rOJQeu2qD1qHRnLIv9Awi1Mr+86ip3T2CnBxXe
ZE4aThgr60eEeaXKKdsQk8fUbKBaz9BemeTeQFzYH6AfPNd2msqfLrR8InOD8bToohGllh7cb19H
TSVsj/J9OErFTmnGfkYbFqzekYaFCxAzNMQK/Vrb3DReZKUF5GDjFD0PKCghoJ3Ofhgk7+wF+ni5
dM/FoaGjknSXgNqYlmI4d0bU7c+gAvHSNUbgE8HGwYRg7pIEmhhd1ZZmptIlV2uiz8n/sHDGjT8i
fuDHdo1W2ogq41+QOn+CxJxlYvnv6Dp41S0y+9/pzGBJJiO9c6w7EghE0uyGpgeNLIU8eUt6URjN
G/7mnnBsaEODH7G/Kkb2E7NArjGQdHLD9ik603J99wxEPou8epRSkFACkvn6kjt/cn4AutwTds9Y
lGuw6xA1TjSZvGnpf6L2yAi7bSrbvuzi61AJZzveQiLWz9XwKgZNfBZGY7o8ST14byZZMnc5r7xr
e7/7AnYnScg7YN/Qxsb4OD28AktlHqanX2pDhI6sc/5Ffxv4GX/W6g3pdbvsapYKv7X8jg2ddxYI
yxuQwK4H95sVHx0QCiybGm7h5rhCjCVI07btwRlevW6K7+fdzRuENi4yZMux0DHBz2/3KD6Zn4UF
OmAvDTRgT74DR3m6KhgycpP707bRqjeyyBFbVXGh8mX/RUD7W+AIkKREH2IYt4M/9+lgGsxp+QXw
iL0ra8piFQ6/irCgsg7XqbIjccL4OpkDVKf6rTtk1BTRJ5EPTY/Mo1KB9csblj1lD0lAaacRmm5H
DRNcBeRaE8Qzzyj39LELgkeSZy2e3wGXa0tvyt8rFaq4g4AZgGOizXWliJquMdiXMsKP7AVFrvrU
sQDeoSl8CFsT+wtgy0jmROM+uzwJRwMdu+n0fQKQT8TTu4I9jIIy7gI8DwrC4UagH7Kd5vrUzuIb
fTAhNoZud1aT11plQ6edAXkuYjilh+lbI6DMSAgqYian78VC1Z0wXDNPIZEzAUnUqDTBoY0J/g5r
kM7Zk/ErhKLMdfNPip3NK6kWlmDQ/elmzghJNt4xgMemCCC72dEWTCgFd3Sjxt8NP9ZZoTmA+FQR
9q/gzUonxJlvzIstD6VYBNNvfVufmR6sVHLk4e2N8hVTewRNwYYfwjodCY4Int9sp8ieNDyfVICM
taGLu7SUKgOFgABVrRG5a2b3GSW9nFC1yDY0Asr1BUGmbFJP7UoSAchrT+phSTFAyOx284FTBIq/
iEA6UPv99xjxSIt9IcAmAjX3Z7D8EDiqJZwcAa+JmsJDvCYNOwIGs2uskuU6nAZO1iA7E0UHJugF
3GvvfaH25HvhoELVR8PYHEsKQvDGPrgaKMS/Y8W4JctlN847jrGoxuAuJ0N18Pfza6HvTyjvk8k/
Z4ZdAJhDtIz5TRLAlh0pnPwg2Ayyd8FIqpOvxU6uEEfz7OJnq+kahkFWYoIRIboN7ZJ/WLINLrkE
TMnxrIY6y2VHyA0OXCxn3Cyg5mHnt2If4RR0PwaLYKYpsm6sPYKMmoXgYuJbGdNNcuQnz9H+ZOum
4tQw7yDjkTaGX4jkd50muThA0qUo18jsStkvBz1kNNLR1GGD5JdSozc/uSPQgqIi+ONLBbGZwFzp
mTWgVb4v0MDVzFNBDP9xs/q1y2iPL1vT41DdQ1JaxBL2zrHDX7xCJVhKiShxiR0xBIelNVCORLFP
OYsprJQcqRg8HEWpWvSNTQrrH6QheiDExOaQiv+93fQTPFX7r29YozirgkXfDq+emOJqBwCCUBD8
iU43fw7T0TeATY8/d/uFMjhCxRLaXTX05xdCnE6uHV3fHx9BN9zZTlEhzUAygUod3jIue6lntCIu
nWuVkTS6/eRw5f9rNavvs3I6b8T5Pq0xch83U0XI/FWaZATTkqtnkNq/CsoMWXgwuDbksmWanBAL
TpvuEoMB6CeEQ8PYJYKA5IXtz0+Upf6iGLsvLxaozt01+dhr8ftc3vSVYQ3HyDcib5/4xBw2SsIW
AhPeqcg+JeVKtbCb5um/i2cKf7m2zWk9l+kuKtI9/7OeSQ7mkQrzI8eClENsEhICGDgGSzJD2gHe
XDQPoqsGqtQzWVWea6XYnjYlsjHSuJAzyv050+KC9xM/DiCjDTYoWd1W0I/yzSKARNAfZDhJffGp
3sZT1L9x9GpuW+jyJV8+I3P6AGFxDCHzdUB4NoLc91ZQ4tkTQmzBBAJ1kWQW195+qnBrl7yXJviZ
yIXK3uQWEjgamqr2GfdIkAVfVSMNdb3ua7J62SbUTC/e5ayV1D+Y5KtjLYW22Ovn0qZtvMFQCt34
rpHkU8C2xKYDdNCzFDr/F3qs8Qv+8hQTkkm8VCyrBDdMtu7fKoTeTwFm1m4baPgIU6RDY9Zcd3+h
cN4yb8p+gLkQsIa8H/USAICuoNrtWOsmFQ0zfcqrV06VkEjWHIZB1rw0EsZh8MA7RayhTR+Hx51H
rnsjJ5bJcn5CyRnCz4nk4wRytZd/YmYnvbwzgtcOMOj0hTKDEgpVKdmNQZI5dPDbd6wRwEhyjzpR
KOzH6JJEalCFcBXn72vFgFhQ2u2+X59BpaGepOahRgxe/EcW/EwudLI3p/EHN1NZgCJbBL1nlOG5
oiQ1n9p+1kTLAac2+PkmXN7m1KhNxKjv9bxQ3aOsVLX7zaf9RREfE5IKHoder2bzYR1cki8JvjmR
S9dygNNQPDm4kqDizLMvfZGeQ1opMHn2yCsEuz6/bm6VZpmeA/zRRP88Iu33WqSU8hCd4enUWxWk
R57qqN+HTZqhra2aO5Oy2x8P0sD5UWDRLLPVyClSG9uEpnxMgLcCRUsRJ94nElH7A4/kjKT8QgbA
InHvKbFqolHYQfldO7SiMQpNRFWANJD7AWCIs6dBEotM7gvopCIC/6DPd8cvNW9liTZi/TRUzVD/
FGSs/Ggc/KkZeb2cOs2YO5B/Kjo+YhS1HtaYB/w3vV8Uubt68V9V22NGuzLN6f46u1iLWseP9NkQ
hBVAfILHLyncX3QdV5iXlFN62rOInogycPXzEVbrBCGXCJo5J+UVtOgxzRxGwhBeUBG+qXEODuqB
SUL8l90CcEE6yaxnBMCFyetOw/jqrN8TCgcXlytQkSYAoCqGrMQDiDa8ULet6ZF3rJ7Xha3HdwHn
cGXisvgkssUIvGzy92G1ObXFJFWT3pyfehrjkePxFtpT2uUYuQeEUARBgaqvD4dspeQgb77oBRJs
Ey4tmeedlD209rr4hJ3MmqDIecrAjK09B7px2Wi8ATtSEM970v5W4ocyUiS9MCqxEbCBUAVrlCSQ
i9ZyR7aVXDsrGzNNDl9zs2373PXORCrUEUcn6ltGE0IuQHRSYK0+/UDvY7//QW5NmVtW3CziAcfn
Vs7CT7C6slMjO5N0f6yFE3L/OrRe4kKTtsdikeTV2Sa7RT8i0zL6wioPvc7/rEenLbLJOpUTqvVD
tssJPd9lqOk0/Fi0tHc1rC5ZW9MSbtSvmNo9Aj960U5nDUgjtXCCp3SrqMzNddHIJeVM5KAJJGEH
KwSB9rZgjYxGbx3TGM1QqpwRJ8Krhk6kanJ7AyS0Et/iF8ZMCGEyiwlHyn3XpWI1vFMA8oAwXq7q
ekrv+MKdRl65FOONFx1RQWNs6d9yErb7ov2VT0QxwTRZq2uJmaG1wrFFn5zqqWiFqwfhWh2kNEN+
EzrKt6+yM5n2wT9W6ySdde3h7mmg4cfw/qDyLUQdAJgo2srYQwzP0+AxQkq5Ru07/xGEBq0SenIL
Fbe+KO4Tn33yaLyKpR4mEDb1bjzhHjursBsDM4dD65I5iRPc0Hkm1kFVj0JfWfda50RX67u9b0+i
w8YpHHH6YyBZiUHwy83/1Og+OB1oxXDLb409wOzX5dccE+bGsXyG8UF2t5TkLoWdUM8mPVok2KJz
9ed66fwUFqjS1yuB0NB6vNj/n7D4mycyodUjTG1p8RyCOy4cwCA68dvgdNybqZSUyc25dw3uT6Bt
Z/qPQoQ0PqI2jU1L7DtpdtUb9FlJG79clZmOBHFh7m7ONLbBORkId15ZwQrGrAIthk9KM0C14amD
B3cBMIW5efAHvd3JgdgN3jHkThxIvU8LK5tmpp0/KPqiC3TTW2Frwmc5k4iHxhIGhUKU10Yd0Cjb
7jW1v6DxtoeCxKqrrhynbOq4zVkP0tz8vbPFOKvKS5+hucHUpJVW9H9VELr9QI1/nazyBYMT7NgU
xJqIFc6AG/vT49QlGu+tsgQTJZSLk6GuvwKuI12JVIq2T4UPqCg2xYTMm88rH+hY/WFrQuk2A4YC
NyxSEljsrPmzDHXsz35eKG8Fh4C7mSEXGcpzLCfW/YoOcDHAJZNddHwIknwyjDBEXChWEiVb7sT6
4vj8NVwwWMkl6ynTASLH3OzcutSXI1ecCwLmzo/UDao1v5OBUh3HO6q7Vapg+Ef/jr/ID1KN3j0D
acMxcllClYCP4SlCSNGkoUkNpDm1SGF8PuvgQLP5IaxjD301JFNnWaZpxXDN0nLjWB5e1uNii86r
6n3ZzojakktkVbFFccv24pnWvuAP6cAWYB9TwVjXKq+ITfVI2XISMuvxB/oK9LL0s5JGl+SaLUF8
w+g8zvzxADoc23rtDYOklSDUl3+ffiWoc1n88/qZzMh3gUYCE1ifFUsdsZFb+Mc71dQgdcWKwEge
NzaThNQcC+IaXooQuntP0ecCIcyk6I2U/vTBi1zVZYGEwjPkqBbj5IfIycZvYZNnpuUd3tYDpKQN
elmOu8J/CTBXj+WurAWvct/wqCYTvB5iTJvJbfsY0kp3UrDbzyOM+XWlz0FWs4oqreR7zk2dOMsa
22XWwyaovif1eHDwH/VGjVFJLcJzQfdCy/npvSBzovnqOlpTOKL+YT00nPs4TJ4E/zl5QhEKcyJq
YtF1DrW8INawX5lpgbLC3LePrP2sLQDZpqMMPUX+OWLCg/eC/qU2gt5Z+NAwGHrH7xUqT+bHSOxM
GvUQ8jZFWurJ/Q7byaHs9gfdzWFV6od74SFM8LaBKoZCRPSiNE395ShdnAQ+/gBGkY4/yJHDABkO
OQ1zjB9QVJMYJ8mRb+pbXgCKWIw08xtC2X4BcpoiAVbYGPbotwSb1DiCUyKT9yVcHADhKiegwcq1
HF93yQG4+aTGuhb7GsezUfglV8SSuzyAXb7LNL4PWix+fuxfo4V5KguoXBDNA/I/dfIkvBy5FqeJ
g9xPj6LDRUs5l/8iJfairXnvc6ou6YwOBgrhA2kprjXnsWpA4hAu2MCNENK6K1DpHNVA/AhgmhDz
gDbpujfE1R3Die8iY67iIQfensTz6DOUDAIuLpPpephTngQkmsL0OmIGg/Eyv/I4wye7BXkF5DQ4
BEY6rb/L3c/N9WX+cMsV91QeIYiuiaCtqz8vDzHlxc2f+nxXxRZUqLdZKjmil3qBYW03YmrveF1s
AeIzd++d99EP58gHQx9NQesD5a+FbORRTRlivcLLkXxtNGiEGWQ2ez/uuEmXvKCiyhLwG5I/M+LO
RTTxIqMWT9WlL/Px7q2WHpv0gQUM4Jw0iJhbi8zhKgVFH14A4GNmIflEO/yQPpYN6FxquVbOuPzc
P/zJb+xHXuEPqE+8+T+SK4WJuNkKvXffo60/wBrFZ1TAo0Hd3rzl+RlsByPY7Ble44o+Eq3B+vqe
SHRbZXkCIhwF2Zqmm4izXI8+XlSr2pQ44xjiWEsXkhR9Cggmm+4D54cfi+ngn5+ZuKPU2S8ChbSl
7IRt4m1aMdViVRFDjpd67fv4/tAsGSVeiZeQe+XAa7OvKZJ5Yiam/VCNC5CfDvHKLapnHFY6NL0b
E5g3JPRAUjuKZluZugt+BO1CChBdHYKrScefB7UidpuqvbWKugEDWpEOlUzFyuQSGX/U4tKrQtw6
oK6TrNfuetpBKfMsoSn7S/s3nXA4oxLGVd063Ew3sg6O/W5mJc95OPi29X3TR5BiwWBUy3ixM7wi
+qoEQ+htvIaDq7Y+xaOVzJohc1xRCqSXzrs86AaehpAi0CaAm8f7UashCm2sgcyCj2AjatmNBKQH
L8lTnyMuTdTt3XJBwJUuifB0HS2wkHS0PW1RhyjRcuOlArEYPtp3ofSahLL/uNDbF+u55hndExPI
FK+m0d+OCHG/5UWGwl+bK8QVsTmZThZW1paJucWtKT4DCZFny+kh/R4Zp4J1WwrcqGAMqcAFXjr4
WKaGGK2qpMZS844TufTymO1JFNnaqc80IfTE2r9czq5oIakjJWhA9a9e8fbjKVWloRMZbHjZ1Zqo
aa+l70yPauwh7JvvyFOuzyrARgrIr2FJA3hT0aemW9YBUDWgzE/Fr36gT5XnApGeYr9OVd/9LX2S
+VLV633vxDF2XF+kNTdqWaSuJjU2hH2DzZshdnqDtSpsgSb4uNs71MSDLDKOQgYCSUx/g3DrtsRM
KbpatFPsGH87bZdGTwfsJmPsifaViDnNDlS8cDzAN6VmcoI/gWqZTM7FO/pWRfsORUiRObCCkrV/
XqUFS2Qkr2Py5THX0bKvv0jFiBf7UbTL//e+cN6JMgzbF/hMZXkSxtHnbRRK8YcAnUJQ/x+62uFD
G6bXm7Qj19QKgIwfmqv3o5nDeKxGj8REzYJeSdaRajs8l/E84vsKaiPsMYDfyb8gunnw+BTKCAZX
WXUikgzaVU/KwtV6JCG+j76j/K2Ue6E08Ae6KtPltWzy0JAaxXMzojWJUhUM2JA2E/AhpPAWixNX
5QlFgErgmjImuFt0szb2bO/7MxPYNsnl9+m+kFn3m/vnZaNu1w7z7e0r6rxHnA2Ty98c4JKlYhBa
v9p3Ip3+DMkzWSH4Kyk9SX3mQrLfHdW0vJEqtpMyCNgy+KTWsU4S3pKRsthRXvVmgBnmJggCPVU3
7BHrFy4aaMm9l5jlS0uw+BQH85srD6HH595bS7g2yaHZMAHTLIg6jjlm4o0jV+To5sUfyPeCAW1T
uWvn2IB65JDUfIVCnI04G+2dBfhGeMEX2hiMrBnl2z7E7zDnqm9lC1Dxy2G0LlVsiI1QQqZkTSXX
5NxE4tkRYZiFLQtXzIQelBBDKHu45cqxT7MI5VrfXh0Tk9e8/1LGEu/w3n47XPX+Q8007Vu9Igv1
lFI1qIGzcxVxCpg+cLbq2/e+NDBYaEfMfkscKPPIFgkh/lcY/vEyrEWGlAZcX0J1JTaqRgox4A7j
BX2bmMVkTL70pLsde8//+orHt0EMhSs2nLDJqf7tOkxb2cbasX+jkQXuS0TDamW9Ff2hTbwkWBnp
HWgZdU8pF/vjFnCxqqmm+1Ts4Oi0K3tskgKiJOTvNlCgN6q0Zfyx4KpcD4MnqKzZAGjuEoMKXbTA
ti4I7hZUtL/SksnxcuwpDC9CV9gjnuRdKuyJwSYMFE2/R8Y+vVS5uDS/u6k/Q1aIzaKcmowmoTf/
PGYiw04wxn6sTnNaAbDA2gZVv+d0G0ZvcD09e8gYL63x7jvaUi24fX9XWa2CbnfS1yr9aFdpQP2D
pwHpbemiiiUy64/8kgoTug7trJIMD84Q84SQLm0+KTIFmr0AZReKpNCY9BzZi5k4ivvXd3ymc9A1
ZwpMrzN9jCYjUzucyy3QzbKoOPFNd+5IT3susnqGijSVC9OChil8kAwpOX6yIJo9Z/eg0payXof7
tXqRaS9ZUPU41/ud6Xj2F+Lli1oSG6zxvdut3kgGMaK64FcAyN913quwZd1sqMzbn7RYVjgZbdws
9W2R1hzslKB5U8icVpI+tKG0uYuzh0flqTjWHDzuT856+Y8/ERPrHKlrBrHPRd69wpFJ5Btt68Uf
lwYqytByrmJb8dw3QYXGfG2aVNUjwfuZiCFwSs0PKNdLAcqerE057ftfVZH4IWXoGq1mIZNzTdWd
7eBg+FiNy1PmQUZiNipdIsPrMARuzXF1H8nHWeVtR44yy2ZsTDXal+nGzW0p3t4VxW1NC1GRtOWx
KulYEFfROHOUxlKutDWMTyxPz2Ac+bMmFQ0ZU5tVt/uOQ8dWXpyXqcC3ZwV+HokeTUsu6f9TfWF5
p6bidpHcJygtqxK2UXBx8cwgLvtFJqf79sYiDc827aYpL1ZSTM3v3kP1IuiVdXD0+MYze50CWAlH
vKm8En/WwAVUX2KfDuYF1IxNlXKhZQS+PUAKfWmp3I4g/ETtaS79SrWtJIJSaMYwtT1GDNHtLcmq
NfH3nKWKoxBxh8Zm3pLmL8CJo0EZWDzsEHM1wkNNJHfmwj3FrS8O21uoJOdL7jWa0OBrklFMwQoU
rU7NFi6pEPKal5+K458VSZDCylQDl4sRPsEf/zXtz55AcFBuVWrZz3B69ban7n/PtdB0pgboQZgC
w0ZhJl/BTFL/OPIR46OwQrCE3iil4kGvwfcJceAQKxXwF5MXCd2dQ3wSTwvAg9fhccHhViC2Nj6D
LJ4H1W3fadHSpI9Bh4MAG6seMI9AlxgpDc8CFHIDDvR63d1uS+Vq+c4aRFTdGOqdiHxbzVV65I58
Lp4q8SCHtPIfsdC1AJcXf1Cwr0KKTZhWeAds3/1bfa9dIDTrwzMmhkDZB2RhC/z2V4b2STUvnZyC
13JAQepveosUyHWFdqtpcO2WRxOnzhjab0zCYhb8tVpr1eylryA0k448Vr5t0XFWQtKcmJWwbqOE
MaXcXOMDN4f5JJPZO03s7dk1U1FrhoNT2SLKsviYuVjHMMIddPtMDyqYA9cfifpN7MSNEiwxqIm8
YQTZm1vjQY2QsAYb8k6tfkCac2D7cyVtucnTomqdHkq2mTZkTVIBJdI8nlAANOaQ74+AO+8twSxH
MyMY+NuwtjwWe21sqSg4feiL+ihMGQyzN8cHlCKl8iuPu+LspdfjFmaaXIbJ8hwNMhPU1VgOZ0u/
jyT4bmpeys7TeHGerjgLu6cpEdfXx0ewqM6ym3DKGToGhU9Vp/CdQEdFL6r5F7wgLBv2xb+Mqj2X
l9oN5Lo2zcXF0zexp+FE0CmVSYo7DmXr6DlJhN651fbF5PLvod9yLiaeAbYPizdQteOtunlH4ww/
qqD6AqTHoSg0GFgFGwq6tjBZR4E3blcZYMF3pQwcPkDCReHvH08hz1ucc+NM+OuiVyXDnhyb4tuN
TMYC9SyuA3ySprvXxpxM9ZvqN3F+EM3FkXFMZlFEJx7MwzN4/NxNqp7o//HSRr6scm1wXKpPly3w
gUuJY2eDBAiSRcy4UOocgjTzKbH37EStik3cy3Q7Gc3Do2fnoByUIEXRlcUvNKU2pHs+eyrlKy9g
TTn2RgUoMJtkwdYFwlWOYIcuSRVV31rHeX9Pl5V2C0iY7nTEDv8inKAuCYE0S4CaLKdVUWMiC5kn
jUGdhvDWW7lmng/t7Ufsn0+FcdB5gq6QEocBtsqptM7vRW4CNzsdEw3y+OMFeWv3bHqCj78Yx39t
XsdtJC2FMG/1/bWHzk/xAuae+bKpITGMlMF3Vaixx5hmzdfIufUiBBZuE4t8RNDTW4WV5imxMHbh
P6HYOyNzXa1dOb0XZEP7hNeF6Bfz627Po9j5V348Ceo5ZPkq0B5ztFZMTKHXAtrX0678hiD6oD0b
wQod70876z5ftqjfWskf2plVYmh/FAwMisn/gYjCVkuOdD8IxQ/mRiVDmrgHOR5c6UJMEUDXRDnr
658+C5JVMSjbXjc55JnE+uYMCwv2E+J2pLwWkmuMcA8jEK69ATDBevwFqL7a0fwmZUliNY6a8J9d
pDY6+x9zRKpqR8kpkkmIKI6g7QQM01M7bQUJIOokYAgh9/i1KnUsJ8ZLMx2iovE6+PqR01XQpLPy
K09wgFqZfzry8mgD84rg3DXSLtfFx4C8qDwSBDdP8Ek6+NTwxVv6vjO2HcCXXVJSg/yAI0LHLooQ
GQ6frpJgtj7t/yOVRzAnT0Tx74uXkBXBGHH0hSn/fQVlAnfGqn0EIQMH14AEUnbOXVSe2ZPM/NSF
eCk1zBzYqKIXlRKq06Pn46OIlRL08LqVBQ9apCyoGVPgjKrdQoBMhvaiRCOZheVruqY4gw8dA5Y1
F9OlfaL6MHZpVgUVBRAVoZL+BEPCIZcdiwbNjLyNh2W09PyhliLVz1Sitf5t6ANnUtl+8FexXnRj
IPPqNoUck8vZYiPIzdGI8qTqg+JI3CPqAYmdxCfcwSOen//KU6N8RD7sp/+Vn8AvGSm3Jax52TR5
fXG4hK+5vdRHZnIhZH/Vw/C54AGXeEzyOkI0vlp+QrOx8UtgNvuHQohKBWNbO4vDZLGG85UddQkf
FUiIRLg/2umk7JVsKErVZhCwwBgQncDTjRgVq5hbbqE71o2o5DT2pKudwKjGKOZLeZ2E5QfIgeMK
rqDweY9ZG5bxUMy0+bZ+dB1TWBlUIxO7qcPdtcFIpk72lstQ/lijPa2td5EcAYT4OmdlK1r/qL01
FNZ2f4WUE5IodluUWZjkFF6qUKHWtahtZrASBOSQPN6KPDVNLMbAbl6r6rkxc3xwBotVsAftldpr
5xbkLPgpK2osQbUBqjxARgIsVIeteUS7l3vY+8gTkYrekODaywTXhhryhQWMkzxW0+ondtGXalw8
9gvt3/7sQZ70Vqc3rT5aETU8lEDvC3Ydzpo5RVEyQejSuoNZ09gvfkD0RwW026jm42kpPrnBTclE
7xo3SKobL4AssP0hRMxY4UFTmq/pj9/6oO5iXcEK3IXDzwRtWB5uw7iVDSDPhokjlKy2HmRVeOYU
XBn7dxoofud5zDCEp0XaT0Y3SHvxB6bcLyEm5h4WPJrIePDOvbNeyREwo5enhA6s3tadtqAQunjM
selwIoS9H7tOpp0dZYJhXa2X/Eblu/ulyPWJldN+kU4wf1z7I6F4NWT8G7qjRv8Frp0M2RrpuzGW
Om3S/c/NFgK/uJhVmTNaRPNhncsWvxbnnhuWA4pEnLSZHlyvZxDU+C8G3AqV1XUeMb7TqYkJQdeN
TNQFkfFn/oxQyvzdmOOCpq+6hDvh6txhvbCYje5sGsi4ldD/ZenPEbd6S1Qj9k0Mt/RdNhxPy5ln
5iQ5JmUBmVvibaF9HK+kTwohmQU0DNN8fdHKJ0DFGcvGYTETIaeJnPAcA+nByq7LrIEntFhsOb32
8+2fF7a69NIyz9p4Ig2ugKnKqqpLuqjg1uYRiSFIWy6YTeX0wGeWpHuwEA38PYESazp+aKnFhBOm
7OcoOgFhx68hR9f1mkkOwSeKnn4ZxoMNtgQVf40UmRq/CR1wNr1A3JD0UZs6YC9T+U1P5ggqQRhy
GYnBYWvyYyHBB0HGiJCclBSIPqS4isZS7mkpLsnmIiu+5ufKNWNhSMCGNPl0YNPyHkghJ/KzU+TS
1hqfjnyewtScMxgSFvsNqCpGzucBr+/ApqSeNo9dRINU4QgZxk06qEfS8igMoH7s0ytWlKbnjnrj
90/nk3ui1qv9PT/DNirKqUlO8bWptdESirP1gLrpExZ74b9v61I+hAM7iON9TIL9UdjCuzoYEhqc
D/KmXfMRDeCV5jg0pL9Tj0jesgUFNmHsifZ6qP3B11uaoCUe+eWxJo1Q+UPzNZ+EdV7qFFpRpk0n
GASEjDA1ArGfYCZRyd2QIvQuFo4+boJnX0u1afd5aNtd78qnX7fkX2K1eMOanoXC8gqmnDDDpA9M
d2ZZBDAGOa/6JitFhITEs0RDXqKosdbiGGlZ8iFgK3V4TV1E9a8TtGfWskfcyr3W/gLqDyvYFRdX
mjRCyBLuANrYuxt30aZhKEfbDadcfmeXNYeMhs7+Qlw5j57UikwdU/1Z0UyR9dt7++AjRexzrmrY
4ttuzSpOT3VYVQOJvDmS0FvT3ntkdubALHQduD13+Nk0pmx+hfeIoXkpRZNPfOJBMlrt62kycWPZ
ob0QVNzHIycIw+fxXZ6/WaFNZ+LDuUSgMtN0gU4c9GqifcwswykQ7hqo18Y5xPvIbrQvZBeT/VeY
NJf8Nlt2lBeZR6tQVyGOGflBLXOKNT9FfkCYAWZxncMeuwsaf2dCEz6copZflNDx44wTLyAtfwdM
wM4CI8kvukh1TTqNazJc6XNpXVjq2GVpEhGFCrg7YYsdG2jT2ISf9ukVbT1JhMpbPfrdAD5/sS9s
VlO7NsLlSqNQ/R81IRGqRyRoUvkDRVC3VHko0IeGQvvflms23pQ+1Z+ncl1KSHrZ4iVuLb5Ma3km
ULWaW7a/m+fRllMDRAyHZ8AnXNBs25FDnJBNCa9BvL0UOlwEOwjOWvweDoEostq4QxicX9j4kCik
PcQn9HMnqAo414ySZEAabzVtBmJbQ4erWP8UGvR1C2OsF2jQYhggscL7Sb8qqzfSZPmfF9ZZ6jTa
D0zqzC65+s2hnCyiBVEGKWNRpFlTbs8Pv4Di8lLP0WLDcOYMTbPXDrWW0H7u3ODAMmK7unM6ktwB
m0MUZb4x1cVEoT8z69YpOPqCZcVhWDQGhKBFbPxjIS6z2MVJ+iDila3+PBlgPjop0oxIygOy4Mdu
IhaixZrSiUJCHW7UiQxiOfojnR2mIMeb5kizeaLacGZ1eFZFww6vkKM7A+dScRVlq6kRm29eYE9B
cEBmLINgrrxxqDzYLO5fjSqtvMKGqEgCa/YvO+hjX79ppkQyDyxP2t3kbztp9RCaPWap5mum+Vji
Gi4t4M7vUXrwjUcdBpuOHAuUrz+DkVqqyl2QTXYYNc/V4uP33NlVSBm/4LukaCVwI4voofqvMVip
frCY/anktmJL1KN8cftPYNPrg64gva7aojBDNr2UbOxH1oCoXHcgkG79rxrGi2elcTIPKctPs7wM
htSV1uiaqQbSDAcqc/+kzkldjL0u9C1PZiNb/RgMxH7DfXPWhT8JzrRT13Hwc0X/AnU7XxTRrsMR
mTOMwts3JG8nKQee6Et5uEinwtit0WKsgBhaZlQgtfLs1RLjKYWVxnP2Dq/MTbaOMyjeZ2EdZCQx
oCEkHvDRKSJYN/IEeb2InH9b9mPlhQYCTasBilg2xxMUveXZOORyAKSXU3tAe1pQ8GbB26GI40Hm
oWmRY54yEPJIDh7pHvqUvf+N9qUS3g1yKqiad95vOleGZpsmpbNA7gkqzeyWcs5yc0xcYwNqYPzI
/cs4xJqzG70kvq1IgpIQE8GAhdyh7QsBR1MMcFrjyocn+Fm/3uPLUFTOvxffqCpSaiQu33CP5r4E
vbom9jJ5ojni9pBfsplMhKjY3V0/wOnbVwbohGzpAlscJ1c+TtXXDAykHb1OPo08UoD8TGvT73Hi
Eq+zagmkUZusdXgoVq6XrQCSfpQI39yU7aOAF12rOJCZ0QMjuj39Qr/iDhj1zUlSaKNyIdKz7IHP
MbFt5+VRKm06/KStHWS3koxxiJZNoi+CTr67kOcSiPoXoSl0cGOJ+hZrsWHXaefgn9g8JfyR+lg2
w3uOKYqlQWDll8CXRIaW+PEv2tyQV1HvZuijSfO1lsm1haTGcwIZblyBUhi81jfitzesZjL5NSMM
GS0MvrsxgftjOevk7t2DuCRd6XQ4yqFYtvDn4MhcJzi9/BUketoI45fihujGDobNdPenNrYzxyFS
8xpYi5obfNzOoBJbAdC2FyIASqkUtaMt6LJoJXbpSIcEe67ttktuXIy3GHE0y5c5XdaG5PBiHvWS
Y78z+4s9dYsV4ZD0V8BgMcy36/k6KWocP4tuAKM6bc/97zfOLDon1iFRXz4PMIJJG4VfkZ9nJwE5
zdH7YQ1GQrgS587IhUGFTIyGsrz8xi2y206NZ5t2fUW9oLmDVaYgKKxqA65e0afbdfnPAOtR93Lv
hbEa+Jdayci8QhmHnR0jqix46LvNFD+bfWNicXxoXqyxT30JG/Qw54eFCLfnCBwhPlNPoi176pxL
I+EZVDAwfVlJFkAUrQ9kh49Z3A7KvoM2muZuWDwGbV5G3xu7V/6PykW33XZREabLb5F+lTVC8OTW
9UIyAf2Npq86agNswIFh7LLHuSXefh9m0XO1Uj/85agEI27Xk8anzbq/HLDMpzk0p6kFcNOk67wA
8uy4sZgeoW2A0Russ0sCn1IMQAHrATk8+Ac8rhawEV7HXMceKWswtkUzQG+PXADsQwfsE4hK+XG/
VZ7hnRdQ80+7A440/ORYkpyQ3QwWPz5SbbONBzI/CIK7g5qnUV1brCEFg3Y0kBqlH+Se2GXNeWNk
NDhQLS4Dg+62i0+5j6njAIKRQdIzc7UHJsppW+tqUV+bBOnrQIeLxWtqa7B8j59sChC34nHeUeUl
tpPYoRRlsDBJvHQhssEBdBVMfF8MYeni/h41mAnS5RSx3ksmEfjzOJlo207kIUDfnz9KQO0Q8cBy
veTPRsrCGH/0GkDAWABmeFJ5OMKlhiOz2PukuuheUJqYdgAQWUncR7ZEhWBvbwXBs0f8E7Jv1vTc
oDjg8y08tHmKQMA/FxBirDdtDAGfmLqPiYKU3VdLx0If/DTn6nt3JeN+8SAiVg74voAuHyOX173J
AI0DEe6/anpFGdIhwYXiKNd4eNhLST8EFEmFGg7qcln10zm//7TRnyoNm/zludtXmZdkIsm9NLWq
tsyobeS9YkuJZroMzKXMy7iTdcNhXRe86j2P6CYRrSBzmcLPh33GJYTsINdqjSAwrxfHGCOGPeVQ
2cokB0SkUg+dVZIeQcLZ645txOFIluXvzs39ckrTd+zBVk+IRfE8cO9FTld8Kvv1t2eeQ9abf4c8
qVeMXPvAWC0cQfEAat0BjqUbBN0jJZADaF7MK5xpxF3ZwVKGWAV0JkuHk+5O0cS2+3fLuDkFNNTF
dl+6chrgPvANsJMupfwLvpVuu/TBfa9guALvCDfj1TPgcPdymMi1yElQ3BtJkBQNq0okaqPfxIni
at6BWUGG3CEh5EKll/+5rJnQsF+TjoL7/sxYg2u4S6IJ/Ao+cNMTKaMsCB7Av8VXGwixAlV56DnJ
tP3EUatRteUC1HSneLMrlGbzFkZmo8Zi4/t9ko+x7BbnXpQDEcqpgDBHI/Cj/NCUGGZBftwvdC+A
n5gfIdd2ViWRmQW3cfhzY66TLFw3i/Scp5os6pZPOlZ7ULcpzZzvlW1Q8VVJG7xsMEn15mqHXdT/
baBtjGPl3fIW7C4J6eOZ+kQOEXrp2SBYx8COZNh/5576jk2K4+Fus8/ra3QZP7TpAaAjolx4E7/p
6oIhKCIuyxmIAxH+pjZq/IsiSg1cS3oJH9LUUWd/b7mnuFbn5ghGF1l+Lr3idE1dzkDPk8jhDfxc
tV1uC3M8hDV0JWydM5M6XWTIUBkXJKvCOGgQDu5r6QEiBcLqTFuh1nGx1sqHd9eKPLh4uPFVgV5G
sqMxJPT6Lbq0b4h6rStj1tKh13nc8kFnr3cezBkoD4SibktLGN436YpakWPTsHjXQOvj62p+j7wf
glBslhPR73hC6ilU0ZD+KVLLx3k+YaSrSFev0AEAXymAZwk8RufBvM6c7ZMok/U84odEfz1Ww4k3
7rGhwpk5PHP6yJjWdlvM13M7B9qiorXrtaDQ/7k3yJJp+IeyuQOTZ0s0ctaNYYn7QiCshNsgQ6fw
pcCefxRlsv4GZUjyrfv6YbioKI4tBTgiraxFEzCDwVvIXK2ZCUQaGAbyLvwkFr/JhdQqXSN8pCRt
jEu7Kbp5ENCaPP7oLdmA15RDPi6aJ5m9zenAo9xEQaRlKFLfUrylw5x1O3ok/rKroToy1a0bQ3Ei
enRIYiyTzFbukgpTQRABxS2djqRh9617tP64+GxLY4hPeiV0yZSLxTla+9T0JqDDfXmSLFcu5cCp
I13YxQp9hSnLATRzNjAH6RQOH1EuwAqjawRtWNrGO4jVNwukc4j0SY0Ha03lXgvCvSMsnIfKhv+X
uXYlzMkGLku4Xe3utHCvOZFlyR6eOSprWcCtj3po6fqLFpCEWA0cMlTWqfTsnXwBswsYCmVhCn+w
5ErHhU2tvo/7z+3MsjV1V6Na8AQCnQAIDDXJUNcPsd2hmdMO65zTkwevHs0rO7HgfRAZcEpI7iRf
9SYqFkrM5a+HFmieVCa8Hgy8DisLUE3BPn96ZwO3eBogbDV0wVa/MWm38sUKTJuxWVAH5zcXdEe+
TWs2mp/pGzJHYIhqLjlFrNlLX9niZhH6UTIhx/S5fVs2wsXsYivT5fzXzAWetK0KklyDt30jv8I1
0waN+TVZE4RFdT4Qp/Yf220PhfhkNRdL7f+E8pNL9yw9J63At4RYrx1sO+wLr6TnIQsQrWVZiBYU
e/mu5rmGSq79OcjP+nCf58LF+tZmIKUpI8nYSfOG9NOpFlnuyFLDSyMvZJsHAaMr3Y924t4m245c
RTMLSkO3gAhDgDc+2valBcfFwPkvKqfeifXTGI1ql+hOsjnhiGNQ7vlUwOQNBBgbBvqw86Pot5DG
MjIsaiZe+XFy3G6KVw8+y3KHKO29XqBNfw0RLOWAvenv+7NGVNjhqxrXKYH1955iT4VzTHWHOROq
epH0CIZaG7Lkp8YvJ6UXtQAEjodL/9ZCqmHAvFBTxOvJd8xcBiMImIhaR3BlBMIHJkRBtT86TOQe
JAh/OcmANYaApdkTszWmJJRpRkto7QryILWR8zgG7ZSpvWzpbJQnq+uj8IEptEDyp0eAdTxXN/it
rYMpjpws/1jU8tE6s4SDFmGZ/J18ECvHrK6jyy8n4Sz+MHNPy4g+6+jSSjJPaQ+3n7KFclV5miFz
ow9l+KirkyrMCI54+SuvlvcMw/QAopd9hzt8MpTG5dkNFWiBnGgTpQLz6q5YHlTqgRRqu80fbuws
NgUa+nOeWxR5vVIN73LB5a0BiP1lh6NqwkUbCODpt7EbnEMIti8b5Ah2ziDxjZQku+DlirBy/wkE
GvGcWQAYku20cb1zPFGALikOB2Ku/o8ltgVJDYT6hPzuYWJIf8vao0Fije6LmYFzzDx87mcMRY6/
RuEIWzWlztFVMVCOVMsemOvUmCSoq92lGibmLc7XzEl+88jfl8o8iqUb7A7xTA0s+J6m1WF5hWKr
4/4i0GqMxqt4JgNMef1leQrHqExPlfRVqIK+YM27U5lwxk0LDHEjzeuBx3aVew3WjoLQhxt4bUhz
oAnFaBiJGTQng4ZBkFbUGhONLdNSI9jLFRnOLjhhyGFq8TZzP255OZjTYsP8qKatLgTHIaL2GCHo
7nPnATFZJeWl5rzVy79xlA0ftX7npky6l5+2pt3F36rbo5yVJoBuPHccORZ2ZBRzsKZNYgQj49ok
0l3OLtFSGrRiCUiVJpR1YMmdXHBhGLdGV44fcsRVopzbdRU0ia1Yy65Ef+Qs1+Yygfe8lvnhMcnI
scOJ3Q0DegD+TwJuDtSbg6wtpXpHVe+qnnv0rDfbHLzNC31W0IVP4iJq1H2rO5+ndCdMUkFxH66q
WcVvVtxNyJJ/XB11hXS5f8qAjx6HM6tda6tb4RfBd+MRKal4g1coiTvDmw4rqt1DdE7DHq7Ms6su
ESNENLEc3kOrY5/htNN6T4tweeEosyfNOr7FWmtGLBesO+QczA1OFcDok88OAgp9LE7XV9hWS3rY
icTREbTcOiPTR4xkU/ApFx+u1AlRLaZtKIjJC+v6DVArHdHYB70arUAQUWG6T5J7ZQ2pLzKCHfTP
BGxyqRfIV+njZMKYvEmYH9xWFdJJ6LQHRzR846XLHe1+gDYzw9ttQVwfO9/VW5Z8LxMuU3n0jTCE
R8iueBdEAfEV4LmY5bPTlXp6vn/HxKBOUXrENMVG07d2IjnJspJEogmdh5/pj9rxNjPQ3zqt+jI/
JfkL/PBrGsu+bQoF0k8DoEIG5vaJaH5PvmWISVOsthegGFr7rtKrx3Sn6yoFm3ZOUrtuac/2a8Ok
4gw+c+u9Domy1g9thlUYChly9yp4TQN88NcIdL4bh9BmdRqxQieei5JcHaM/pQcZ92U3reUVLxTI
W3JJhjGyC/SJu039rxtd9OUtOIGTbwTb9htdAaSA3gbb+VZFDhHfnHyxLTXTLDkfP0r7683vhw2Z
CWvu38mmXPki8jyc6AWTPDe12ZdmneXZTZFhVmUd0ma4MXX3X9GNULgIAnQHCRgfyu4aPK4ivnaO
L4+aqJtkDzwRWpBhEL7GoMcmkbFMs0WaaTQLGqCrdMKg/vhpmT46y6Wnpi1EECm9YZccMmMhWHMs
ZcKRMgTF4gqk5esyYvwr5IXp3uYjOAG91dunnt4pat+JqB0N+aCnCyKpOtcxL9QAayAHdvM86mqq
JpF+QQg1aQam+Ai9lGz0YwUH8ryOb2zP0xSGdsfgdpcDYobAPgvw4FZG4oe8YJme6wJY1MK2wGgQ
2muTu/qmN6gb1uZ6iBMxQ65EEhvEeP8qvN7qqfy7MNYGUq/svyKMAB2nY2gC1lIPKQaWwij8/aXO
e7rLLl2DkppJ00xGjh0lv4WddXKRVRxoAcMy+nWt0yH9VSnx0Q6b+T+E67Tno3ddwGo8yiY+9p6r
cvO1Q5YO7sIMNkcSM0Jcnag5VUwwOdvTdNSMWa7KnPOOL6HM9AYacBpIAMPu6oaYhYW+L0/rf4CU
wMhucLUaTbFv4YpP6iFAHjrPho1isV+Qdf82zCvoZV9Jegx+pD3RVaH1IxrsSb5tW7zKkXMd5E8X
OJy3jol34Pzzpbv/ikYgijfcyHCi2WE3IliqK7pxUtU74JIzHguMeXruwzEdu95Ba102Hmm6yp2g
UdVl2JxXygd7HybZ5wUB/FBDeRPj93lK30xL/KWNtETdmYu6RGtdVHMGkwfTyRF6F1X5Vjn9evvm
G69f6O9EERSoMzpOEmXXbI8BXTHgdGFkYmHJnavjBNlOVENPiVupXazJD/NuABvOuPWMBgfbxyxs
30JRBwU8TlIq3bHD7loGl6ujmezsTlg1UFw7S5/7gA1lL77MzOMBtQEEl/a9S+4jehO1cqVAf/va
8rapPN+GUuTFq4zEXbsvo1HYkJaHVDkdWJi7ujEDoUU4W8GS7dSFzzgBACJCLv4UNRnY0yDPOD5j
iysxaAMMaj3MaZfsFpvunDBsVNw8XZyeRB+TNQBoMR1Ri2dahN1syP3JxgHTJaEXTxAkGCjK7EJW
qpUh4T6Cs5ScbDNt9HQnVVBpxt87SaLveAJUeCPcLwAOLbfuoM2dNqsDlhgDh0QpOP6kcBMCZqqT
2qYXGIKc6/Xqvst8Q5pDqzcHMzYfcOPV+25iCOsVL5+Gl4Nna7SW9A/+GUSL2RLXg+WiPZVAYkxn
Zn4VPg0+FlRDm9e/RDKWhyzqigT885+NXgly8E0KQfGUdKLomQ0J2gw7k9JEvNKAM1gegulIiUAu
0I1xQfqTxsjQwBB3DoRIP0fcMPRAB3MufFF60q0DIghiOPVYeuFv14Ee090MT7p6PzblIeLn40aG
KXwYosf+m1oyfb86Z7boAQXQedE4k8pnCWZjpD8AQyrrx6e2qF7imCjN1M+csujHow8aMPUHKCMr
q2HHe4hxcVsT86oQTuu6EvLWEmXcwjfIaChMHbAdBUN/txxPQ5goaCiA6s//3XXwlcN+Brb8G5+I
3ju5hIr38f5dASYHqUPW+zEmuilt1/XbOUcIXRKMAZ2yn4FFYg8xu53yX1kp8GwHZaf6shh/Hhgo
Kzydi8hjPQz0pjd4hsdvbI29TL3ocIr+vsgJbMRDYUdmbFJC3Kb5em9rFsVkPml7nX0C05oiepPU
paw/Q18SA+Ej6NSJMq9FlrgncWt+QIT5DzISCB3vHXGgOplWyw9vYP+u3kzFUYK84lBkL8/2dEo3
SP2tTnk82CwctIcLC4KPt/oQyPZo5+hJ7pjopSehnXtmihbxVH341i+gS9mMrdxFF8kH51MshnBQ
jjiRIGdmNz0yX0d4WPt2oRUq0cJMEgS2THcbHBKuZ2INozqz4B07A3g/o0YMa4tvtEtdwJ6Gqujx
kSo9vTnnLITdYd8RpxtrfKH8/FRbW+GRycTF/RPyfw3YIZTh6cznDpxXHGhpNxZiOxAidVZ3tCh7
u/SHfMv/++URLVaHEQjhEd3hNzG4LLDm2fry4lnsuGN/JfZ4CfD4HFU9uh48Z/68+vk5LlZujK3O
42WYjvIDnQqjg1o5l97agh8SCCkQ9yYf5f3O9yadyM36X0KKmkklaoIuCE6O6Z+T3Taofk64+fjQ
G3lNF13gKi/nLmqhHBtSbJR9aV3PxCrzGayYg1W0IjlQZ2cSDmo0jw8Gspwnf5J09dAYUx1mY1RK
ctY3B2HSp8+xXdB14ErVPYkCwLCrwLJjjKSEhuoNvQhEhCtWWVfZjEFhARFIpeFcKGxCsTBXqFzC
TsOiI3Vb9BzORqqlW+9kQ9RUdHZ+l+Ux830YZpmF3JzbGOwi0gP9N0WmX30AUcD0Om6EXKf9K/Ab
t4aexFxHKf7gdxg7JB2BIOFsp6TMiqjQszetHw2XIdqeDntENxQiHozikHeunHS77nu5RkGA/14G
xo2ZR790FfcgEnsWW2UxkbFdfqMrV6NGUtRW5jdShOhMeAe9ZrKKbciybyh4/H8D9sbWf9eNJ6h+
t4HZetCK1aqyT+SbHVcrG4DT9VNi5fApmt0ODYu4fXIOamWjFimnjkOi+oOadBMHoM5BkXnGM/7B
4BNZ2INkNb7Ji2MmQlASnH7Ca/OuM8S55i25Itn3QDOI24um9tCoOlfoiJfbSM/ylgp8EBRuVK0l
uecAmyjq/Sr9cSqNl80q0RXsn+XL+IMCyjG7Ysip9rI5THGbu/jXNiYly9aaraKVPernAMUgEwzK
Cbi7memY3cgi8UDISUZ+2ArWw/QCqQJrnQT+aOl8MOkWG9jd7p3v2/Kyp5qKvGFKM5AZAeiZzggP
otNST4ptgWoKBZzsW++jF1QHh9T8Ejm/LAi7fXuFm8DTVDDQXEnQVx0DENeWvmL1JTzsUbpoeBDk
AKMAEkDZIcd2eEzAWVjZrKs7ntfGBs4d6Wpf5dTZOp2616RA6Y5gPy+v+pugJpjbTqQxOnpeAhZQ
89f+OC91O+RwaIG7ILh3bY+1ybmaeweAkGdhVjPDET27d6O/oVuSei0WDfHjnReXOc13sPi4L9vS
yhs8h7K1cXDKbzL0Z+fn2t8p6M3QwMACd3elStjG6T0/AD2QPcCcYhPE180Bdj5AoUnqZuE11N5j
jUDDieCZ5RqXjeDQG1CbRbygoNZYBro8BZ6L0bV0uLIFZ/oo4l65JkOfi6wmARjqZN1zfx5CpfPH
gsKhvA6MEag7GDmBAJIGfTDWjku1HaoQ6AGucbD12HG/AnELegW144Mc6pJ132GYNMowmQ9v8GSz
NFnQHxH/p3tF5u/DPc+1Bn1lhwuzgMtGJY2gpv1QhN6Su+BxWZe+Qv3GtWkDzN7a9qj8OKmCOjl8
BBTwsyIgGY5Yu5Ce3IekpfyUPcxjX/dZnQPCBPHtcnZ25Ok6g0VPh+BbNpOOurDxKO8I3QQbRlvX
ReUDm9+AocejvPiZmDPHPp3ddL8CJSMrxwTTgudDZerXnoFoSfm7fxLPVyQiXe3Cv7PR5mhV0S4x
V0Hv5HZj3v+HQTJYlx0X1D3fmWvTUbJzbvRfsQ8W+TR26eE9EEYrE3eauMCww65QQA0CRqCBdRBN
4BdBpmCYsmBLL4gABtciOAAsmNysrHdEpTnwJ3+s07IcnullpVdoSxXna1mZTlCM/sNdmxnjdBDY
3iaxe/plWen2DqIUTkN72xojUkL/qwdK3mBBxC6GD/k6Rh8JL4V2whJifTZUGM1GC+Ti5By278bD
aYHSroutu4p1nl6g9uBb3glTYdW8AV/cJuLa1IgNAKyQHneQf8+gkrTaGOHNQg9b8wD9cWDmOYUI
abrXlYPNbsyisScz8zPKLhoT5bl3svhrIk4asZqzrzptRLBwK8aW/wZxToOFblV8F6vjx1VIBJXR
tlw+gR7VOtoGrQOIvEVUZxrM6ewl8vLyACv8hRE4BbnpMEwkhe7tQHwMEbppe/Fj8xVkHejxz/v9
aFxXqQlNZJ760zq7coOTFKC0fapQVRvHztg8nsuPmSv9Lx3yeD3yzqpsdAL+OGEVuWVez0bGQGLl
SLbpbsmEMng39Z1GfTbpN0yZO+2hlbIAsy8ugcEOQR6h6H/ICeD6dQ/497viQ+kh31oWCe8d9Dv1
rVE7TulEsXsnMQ6IbP7IGRhwsLXbaHV/I1Y7bEVKTZcG3+nF5nOsxkFAA/ieiBjMB3a0gmTglYfg
zXSluIPCDQbR/OaLNKvLLycUNLyGzmse9jh4zWoYSp51/NgYqVDJub+AWh4mQ8m/G3/yBHPxXi9I
TGKGwX9xvIBfzLIa6JpgpzV6WVVnhuqgxYmcv5i+DRcXVj0HZgAKmlLZHxzPtzLwJIEvCDYjIdoI
cmR7CmV8Gfis23WOuuKK5XZYP2MH51VGhXRdpwAwnXjeueTgfwrs6/TTaW1tyKaH5aVq8fQ6s5Vh
6h1ZGN+agkxjseIHzWG8L2J4ElMyR7VdiozyGv6uIfrO2T/yn9LUg9TXKm4NrRXxXXHne/hJjyHU
2ibao4uWPTFM1hWiaNK3qvmuSiycrJNGibCDzOwK17mr2Os/DB9WBT/MR3q6WVxvXUDwN+JwckaI
3u+9gVYdmZoRLfh9WjuDsbvfogxfcNLgm9zALhY2eqSvS7KDuPktLp3p/5YkxWq/o+z0fOSo8oni
n9rjBzP6M6y5Dx8bR4qG400I6VLvqFb8aLjOoshHHo2og29CqkzpP4V2tsJqPxCKv07jVepqJOTw
qp+l07lbAHn3YwC1IB7VPGPUjOtKoW6aIY7JUzGiMoj3cRwYNe8yAy8Hng8HeKmMKrIFHCgWOQod
TJbhP7mqvOUJVz0dagLHhO0n7vKFFhLUKIfMzoOKgw0TO5qA1MkV9jHX/hBVB0TSP1zQMyBFz+R/
4s0dNG7qvmU2N6PjJWktHgYN26f5RcPPfJDZCep2TfPTB/8R7CpI1ZqLG5DN8KeLwjj56IzriNt/
WFtt5o4EzR2i9qq6SrfX28DcPI6+HBZgkqUPmpvopiupk+Jgjr9CcdnJ2kMmXjrhLk2+OzLQXD/y
VssxWG2FLitq3M4q3xPdoir+DcQHbNgI8ZihQ6Lr9LDnF8YwGsjKUQhtQXpp/+K4jcNfMRG5r2Fu
4hqAcD7nCZCjxI2+QEWhlR0wC1OUeyNPACVO5IdN2HX0LQhRBrMFErTZ5l7kniChorv2HXJFSNOj
vkUgZvgNBhGvQbIBePX7Sloa6AvkXmBlWe6KpFz10U2BJi6RuLOt9qN6miPKq33BEuHt9h9FX4Xa
xD5QS7TnANPu0EPFF7s83u5DSuRW34XUxCnzFJvvvchumrozY4AAsMvSQNgZXzg9AE7rG3w1cwoK
PQJYMJmLUnz5tYKpCY99Qt3CVw18F0pyELt9vLUyYQ5HADXdCVr0SfpWR94tDkEC8w3CeMRz5z1O
sfHRP7+nB6efJZfaViRkWmDgEF0fZVZet85s3mQostCdz0QPlonnsdAvElKOWZ1958/re6EF1DRZ
Ql7nm4PrWoJjj6JIVOmeGPIOwuIb46RyOHs2UVEnf0wf7xsS9DCKqaleFCtxDDJXgazEvJAPO6/D
P9U42+5R6lc0fuSheID8H9gfNaEG81LYTsCF1ExoLTUGXOO27fFZ7tAnsVcDnnukEGq1djcmYtJy
QGXwI0PaXseTKO4GPsgdIETxMDd6Ik4iglK1XfNBhhQgW5nWZb4DZkcskebsIJKcwMvZf+aoYAGw
bShjN30ZgfLP3+r7e+qtjmOnLwhUcNoW8Hu6M6BpnaeRsvyhlLzmkAGkczTPF9wsmcQ1AbOFay/L
yLD61kyz4xsUntwIyp3pybbvUHR38Ykk1xlRSfBBoA/lU0OdJC0nxDNfISRFeu5MCwTzhIRounEH
Ez16rUduISpkTWYsfdHrLf2/cSR9SvHxoDT3kZtJPM2hFQEIK9p0msQleyVkiza9aSRwvTi+P+in
oxv3c/EoQ9Viise62t8A6FiSGhLru7mjs562Cs3rDjoM1PSR7ehQwOI70JGZBmHof2DtEVyvLbZn
4PDg3fgrUJR6n0lnDXWvrkInKlVguV0uOyzgaNWGGReN1xYBmg/665ieo2ee6cKEUzb0zR0pSLr6
6XAbJEUQjxneBA/n6tOjASoqMiBkTLQybIaOgHFeXHiZ0ZNHQJR8FnGfpG2HYoGbdPzegcIDLtZD
xXHTzajuZexr5fISAYST2kyIyxnomh41zokVqGRUjcSNLbNRmkq7tXgEpo+sYCpLPx/No7qC8hoV
Xy6m1h7FSyYj6KvqnZBP5fOyuzwcFjTS+lxMteJcGscvDCxC3260Y+fE2CtNhKjm0Sl6QX5VgJre
AT3fk9epdtmyoAv5x7PcpDrZ6Bo0sX2/KxIio3dSnchHOOEyd7mVEMv4SxhMLlpc+lwlEEucvmkP
P4j6xgcbDtzHjHBntz3yTdyBb6LVaesm/Czet4149Rpe2gzHl2ULlyYBpmWk+ttZUOVGq+Pl347q
DPVNy9itqy4QZ4IXby84G5kXmffekX1wjspMvkam2uEUGpDuJhJwKmmWJhRI3tytpOnIOEZT+AkP
erCQifNe1venu1ofjNCpyYylTguaFplRuDNvOWLMKjUTaKimXxPkvy4RhWyNUiP4E8V3DWC4L+z+
bSsDV8r0kiegHL4200rRYv4RMMGkGjI5j+ELgTnB+MLpFZL2D8RCocKViByPGjsuv8cqhH7mGw9X
jJznJBtnYIPYJ5bVqCL4JKuW15bX9ltPraPOE7K3DkO/jTsSjaxxKLg4g+0cA++W+W5zeL/68Ugo
sUHIenylyh+eofC/yYd0oIn7djMcPUohCntXqc9l3UYL/Z77J7v4j7I6jDrbcSkXVt6xeHRZ8b/b
QCWYYMieal2GLHDIe9Mq7hJi/bxhGBgtb+7hEQlupVmzH7pb8jQjxJOBoG3VSVx0Vwck3ndHBz5g
fl8UDvIRfUmlDrP520ZbtRJ4q3vLUWsgxI+4+xskKN6tX3Mj2EpBAGUpYkznADVPEvW6baZGcrcj
G9vHfdV2oUqpgAIqgaO4X3t+lQi7W56F95yN4R6Sv4BddzZ+2zTzeq4x3KwxXbkoVK75MfYaIMxp
tjJm/ylxQ/SxSq1Z1Vy6cBKpnXpbrHnUycjUHggc9UrLnV8GKTM3eu4KAz9Lj53vM1Hq4luzizuH
rtLLfs8JZtYoPHIaCS6jr+BaE/iSghrzg0/+BETr5wH5jyoL3RFgntRIUVtrPKrm6U+atXA+XPW1
Yn95fv0giRd7LqQr9IaDl1h8Z2aVoVfmvIqgEYo9Pueq/j/i0fz/oPbRwZ0KNvr5fE/DLBzTBDHP
tJ2J2Tcxo6i3fsRHiMUFSM0+7osqL2C3/XEr354E1RjPuRNRowwbFtqIlGf3taCnxOFif77usK52
QH3TmEqEPkrPfSwrvon7gfgFWlcs3XooGLeHAE3pWhPXGzqT00hqdKvjaBFrCwbzBhm8614FdaCR
CpHbk/J5EEuzSTrO6OHj7JMWUKVxKQ3e3bvtGMZOkmogIjFPOw+wA4d/sXnKJ2J3cubRQWt5KtUT
0QMHCjJeimEFzlNngcAlIhjHXROQS/kdksrHQg5cimykKMHcYNBNnkc3gQ/dZXGzo4KtLpbEYBOH
KDFFixwEfNU88UDEAW53bn4fZD0GzOIw5CFFRPDpO4qCT1CwXEGs5SZ8thOkiDNE3KfAtdm89xGa
rv+tfWynYwZ9kCVGcadlkLjBCZ3Nwh9uwnthi+JvQULZpPJEYL/aXz3TMIbHSI0lSmpjCSqb4yFA
AtLkCIRAUsG1Hi5WL/DD7OAGPkud+EPECpqVSSfwZddVc5+RdOdThNFGap1M/fffTiIY889uY5ne
jrpn1+dSDLWdAuLwr6sw32D0R8jLVLe3jGgcFF0zmQBEvxCvgHUrGtHoIayEbbR81s0LQFmA8xyL
byS0Tl6Xcpi/Vt1z/EICMDM9nMrq08xm5bzu76+6zdW5wzoSdj5WvQ9r7yTPCqlPIVvwRdJOL8jQ
JSL8IYNTDYocNgIhQDHTGL+0HfQ6c7iLxCSvq1T2W2uayB/CxO9GJVdzT731uv6YFDwCExyBW2j8
FL2/XO8pERosMPvE0HkUrV0RfbUdSYKXTlrdW/FPJLskc5vobitfSDA4w0vrcGn4/JOKrrXiVPKK
uw9XAco0/TTUG1PzgvrIxLle/KK1jGkQlTelfYvfXPtfkOEnDBgE7B2Ovd9D9KxgHJXmw4Mz1bu4
HQJ9jHZ2rzFGPf/H2vuD+Es8+ydLG1XySZfIi3TItg5kbAMXBruLPt7JxRKaXOsvSr+Xp+aDGcvS
wZcLAtNjCHkv0qP3fZz/+7AuUsenqBZyW6m51YO8Em1k0LxBxWMCUCP6SZEbLhEtZVvAhjQUS31B
Ed3dwSKWmJYH0H2gZDRVOXaWTaAZdRaJnmOI1suGiJitJDw8xtPf8y+02t9C/1dhJFSrdEFi1g8U
UMkIWnC28CY0ZvjMTSpYT3d7v6MNKgiMZyXT5Iq+o02sugMdv3EMX5q9//DNyw2EG+XWkHIbKjEc
3Vmm/Ic0xwSYlQ1BTu8baQYREYchHBJLUxNo8HPyHi/NYXaP4GehAlwSF+oA1ztNfkztFQusX8MB
UGAZfYEtoZy7SK9bCjorZk27AcUFQWHjorgwdcnQGMsKbWCv77478FpNindZvE4o3dYZaGTSnZA+
v+swGvzJX+BsHJFJcazLFi29JjceKQ7JH4auv6uzwqhqep0hCMs+1aJtH5RriVY72BLTj+QGfNQi
/2ZbU6zggsNfiMVTOwVl9ACaAEwClGmhMZcxS34t4lYI+q+VCiU2XWe2gzu9adm/9+p/zGnhXZGX
pfimg873VGpGhwrzmFWKnNWcEFX8L+wuDATmzUmj0hsPfQ9EuOe0+lNEXooONffHMGyO7cXuqm50
I5MnYeWEIMLik8QkrWlhODwIueWmbw5DftOIkyOfhObRADuuE0S9WWKqnu2bJz32FTt8Hk00FXDI
LYjODTVMCLCC5GhJ1l438AtMsHPM1u0qHeGpBjW4ii1fVxlLimcxNG8wDrtQ8dQegUNQ24jG89eG
0egr2wkvH0Og4xw5FryXd+uuhMXx8EJTlYeYs6JNAfEFQs37gXoYU4lphMuWhDpCXNm6S55gfv9d
5LvwtbkrHO49WUCYVUHcFXin/9+uL/2y1X/CAOdFLiCo+V7gKjvbO7LOx9nYzsFMF0WqOdnAWT5B
uyN1a/swX8F+hISY67EKGVYZufat/5SlWK8c5PJaGxyKzzeYQwTN6ykxtuZHYE8Brs2WSDHzL+v7
26zzj3S6+3OlKhMjltH8+Z8xCFv8IEa9K9YoiiiyDrCxIdrbM4SgYu5IHYjLDAn8V14dlmQttlyY
KKKiUcIelVAOoU6+8QybuI1s4SqJdKP7tWS88iQTlqKbBtMKzlU/cvQFeAzj9vWABzEBYSquH5jK
cbSgRnQG8PTIsrHodVv6W3BBbO7b/Wf/gu6ea/d4P9mYDaIv+2zUg2zfnHLP/vcOXcnNib2hvYeD
QXf48I4e5bwLk7uyMM+7oERnAo54gUrRXOLSuyffjCl8UY1LlblUrH0BSagmRdi9X9dObyILXfNu
xO3ja1c+EdqwMiAusRqxrM6lXhglWiTA0+kkFkWHtMbMyKl+Q81eq8pYeImtfiovIUFZLSOqqslh
rfyITK7KWJmyMwwbMHtSI/1hGWhlHv8P7ZyRBr8I1omviw9OXYlTGrgN13/RUF7mExKe2oXk0/0X
HFPBaPS56ArxAjIfCTzYj4i+h1Qx4oTAwBUcZjNou3iSiYZm8yLDJ/izUzg6ru1eTG52nm8UZ/OO
LI7UmICHy2u0avNh281S3L4mxm3D/Q2ZGqXOZzhRKhY5IaEHIIbsiTH0B5cbLMB+2PMvvkEj7Kou
Lsv2eOnBSGjFh0OnPN+vitLMK/AHP2ewqk+uIviLyRUN0WYCXtYNAYOF88qtB4G52fc5KjmdSKNj
dxyjAag9xhOYHgMjBpbXob+QPj3ErFEqjICpkcvob6easnLACgj6duV7tQsy5gD+wK1mKz7Fz9oW
zkAXIjhx08wXYqymwCvQQmVTexWW95nZqBGFP/HJ4lBwAsy8OYy3jgfseuuYtdhOclM7IFpkOKfy
vKrkXJqoufUkk/kxbs7j3c9GXc8ROnjjZmohlW2zvHok4OI2gGQUECDTcNEYLMkAX/2rm/Qa5p+x
cbrqkjlJcIIhUhnx/sOZgoEHNxmeuJwJQghVo5U5WLXMokJ6DkF2YLxSMpE6skq+1i2zjJKOgye0
cvGOP2Sdskvg9+j0zMay5bMDqacZc7T8FY74dq0ewwkFdquxuvzcbsfFnscFcxaa44ER7j/pqm/9
c0wRzzKaf7wfFty7NKujGmiuWnmXX4zOHwpEm32twswWPb8G9h+1QZxic6BXWmmsRt/YA+KKxyde
etbXU1f2PKG+lbzK/Zz2AD+zHz2c/SdMp+p4LrCp2A+hLDxO+aMx4WuHG0zQmgj25Kj01OPJ/IXY
BvIv/6gtHVkNj/CISlnhaxCmqrv6CLI1vnjenTfFYqMfOaUcGsw1oJsU09t1Jn9L4W9LovVlnmOo
6eQF+w6K4GRB7QzOKt42KLFE64EkjldoAl9rs+yX5t/DAoqXcdVYoRDEnKTnWGZqT76MqMrn3s2N
bgLBn/E5n78UYhLRThiMOKc1RRlgqqxpER8F7l/fOOoJ4lGFVfI/dRjuzO4Jpsnj5tlChuw4lipo
9D7w/yldH8uy0Jt32CL/ohBKcuDrHczttoHlDw4drsfwR1asJFQu9l7Wofv6bIxabytiKhu8/M5G
6EhLzcYKELI92jN+MK0cqQpFM/iEk3VaC49RURXYmN6+tZ+ujAt4YG8VALja0zsPxZfxa+/PLI7D
g9auAqJsn7xh1tRpFKnaR1dwDdk0Kf/KonEnw5TQLA1MswWN5QjICntm7ALDax4FNKLYqR7rYULJ
RyhyhJ9jFg/GwD/oDv7ld3V4lz80GOW11lJLjKiTK4MSKwf0nTcixzw2BQTKoR4iYn1NMYLQUFQw
Mg6bYSwIWcv6BAKC4/N9iIOS9urhiD6zppp40cwxv3N8T+HGG50kGvsWKEvORo88lCZ8tzmwVmZR
JGOdx35eyeLf4SkEgZgqcFWoKvbkKKRE1T/8HkNIW9ZRRS20jXpKQKhYGTLAP/Dzwe2sTkkFoj3x
tm0+96VmX0QxKFssbXDPLF4hON+oy8PRf8KcHlXFlJkYLR0wWNNU9JAdt+7h2RINpDJ1Rrpe5qL9
DRERrNVWEeRbj7167W64s+ZcMueeMrVOAMnT/pp39pe3SSU0xXTwCSyF31UzEwgZWC60fCuydRug
y5aitFmso6THEWSPFEMMMQsyV81DHtwZzXOC1h0SQwPzoXh+VZ0mTi3FHy4jL17Ng91n07NzDmw/
Ht0NHR7hTeU9+0Iq2VXeJ9cTXT8Ji/svm/sw0HG5dFWjlMDUl5s2oDAtCbd3lj/KXVAmjOz2aqV6
qcwP/nC08dNUgOHnmgTusm1LGIPnduFJ6X58yqPic5pBljJsZP5zmVMPCV2Ph3Ls2IOqZ5FBnkiN
PGe7kkplxjdMURLO/OpzN26KLMak11DAz5VilHKfDfJ9tp5h5WndE1WX+hK2SnPpQ/abqyd1jEAO
i9E3s6MPuxMxxnqw3Ljb1//1BxvDAqfXJDsISmJ9ZUIes0R0zBZD55WQzNR65tOQM8NzZim7GhHe
zfTNrR0tFQ/F0I4YH5NLlXYniuaN1iLx7kHerXGUnAN5iTQGVYrvGjG9dt1XS5A7oq/wodMc1DSO
WIEBliXz4+wEfotuR0G0PBy2Lfx6CjvmxOXxMIDP8+o2xFnMm7RoVWovZZk6Pnpbj3n11vHnFRmZ
MgFinOsi2ytGqlbtlPcWQbJoELTdrHuQCvVVQxLsTij8neAUVe11yyLoaTk+A/HT8LS3sWqvZXNm
jclziVR8H1m1gM1vmXZ8yzHFPQ8AVqcFLtk3oQ/yZDcM0Xk+9T8jqiSmAWxI4ek2LsBAcUAzkdb8
FydJpBCFD5/moRsjGoizo2yjMSeVVulJn862aBjwJIQczwwug0Vmn8773xO7k/DnOes4Z0fYxNZd
dhkvuJ3qAsN2t+FwDpm0LFV47G1mRkyVQuaQ8Va70jEfHUE8xz3osm8uOqBNK3z/gew4UNVHEc43
48JWxUZtGl2DBYQhs/kAfRqwfeBBNKqqXlAAi2Ufi6O5bqEA1jhY9z4D8I3YokIcJovk4NX9Xao1
2xjETOx+wEaIlAet2a6HWZgfqq/+NMeaep+LrKEp10MKH2vWe3QubmVAE7kJBzRB7mImAgK21Sf4
mVELoou2NtKMi3xOEWVj8VUFQnXfodOqHH/4jl+0az6TiGyGz9YVdtou/JxCO+9AbtryoKBdy9+P
+YLNrr/VHDsxM+TSduO/9CpXJRxjt7zFNgWrFCaS28HCuKO3lOIaHyFTQmxfLZ+jeng+nmUqyHTf
dkWXfL0phv8suDbV2Z/+iAoRwyr7HLZk89ERXriTZHcyXFtCsibphTNenFFZFv9350wNBN6trhfR
JWjHozlRkB8YVmzs4OLVWLg0/ctjomSiY03KK4yu0F+0XN+63JG2+EqrTGoMvlhnKZxOOUo3PKbC
9HNWVuT+DRcttviGQFC9DMH2Ad3gyfTdnAk7ZnlApg2xJtgYINY0BCzYasf/TrIypavwHqzAsSRg
T4Oo1Z5RnaGAska0rY1lQe80rCMH8BaqWR/600pq5yfjAUDETvmeDDMlLMxXH6wqAoTnhhuY7rEm
sulE1siixpPXjnQhkAGQNxaac8UgwJgV5eddGKOKC1whZj7yHfCCgU4s8yFhw3eMESVjr2a2Oyul
I9zTJxEUb3twPI8upMBeL8ahlYPZuY0k/jaqMapUIUq9IAs49cHlwKm/6VsokUvOJvEZqiVRlSlM
QOt3/8R/KKgSC13XW+veWOMB6YSwTljYM4SjhCNr3LsXZ9SIigoAo/BbUZ/hhw33/+Wi90UkRVaW
EQ7WkQYPHx4rOSCge1TAjFtMrWZnLKW3Mr6i0sw+mKD4ZJG2TspShJeaW8ejnaol1/mTSqPR5WJu
UKT/Hea6O/E0puUK6NkoAkDe2d5K45PZROpCOpVUrqAganNPEN4YRPZAJP4oeLp2habBOVeuShtC
kQZb2wSFPHxarMtzA7cqdeU30kTBDFV/+/j4+EGUxPo5sknC5ZMi7SpwA5ky/amjV6PlqLh8/Tsp
N4UYEXdazJ4zfInw82XH91DS5jkAMZXabPRg6or/+8zepPerzsKYPRyos+1N/kBZLFzEMxua82L5
86/gakY12C6eE9/uWOB0je/bolcYb4wDwDQc4kneAgpJKAw6ijMFYWvVWjnhBQ9CdaDyC8zdZSGt
Vcjvb+8tKdbIdM6IgKVuoiJKmwu/edWXuQVF5d7++rXCyg2CVEWz02/65m0NPcJtm4tsy1z6sUET
tjUIuogClc2OMM6vigkF4zk+oJGwPUwKNSRXGIwFwKB2Sl229+Lxy1jk1NmUvuq7cf2RVf1+iFlH
xZfVXUIoAeYqClxa6hwnhgS/vCoAdB2oLByXmiR7zo+QD89OhBqs3eBdjHMLuqr1Y++3XnyZIgaC
6x2j2fYRWSR7DTS4RTvMhbjfMFKieuxQJQI3whbrWwvBKn/xbtjO+snd98BRwWOL7a5ruyv/n/cL
zPsxDyY1INh7cbsx/vy2idMnOHfZUebtf5tttU07NYpz9kCNetSO/XndOiVf9Wv4d32QBXUwtla2
j6RIjQdFNYmCeHubGZS1cYe0R0V2Yw1UioIfQdAWdcTJzlibrmcTO9NR8AofadN5KBKDBDeW+UHk
fy3QlRctUg7Cnm8H855T9nz7hOt8Z/F/NemLcMCnRWz9JbtY/IunWJcKh/hSCo2WYx+H7oidy+UN
sj/BJuumkhuQcEJcBngJ+B7hjMUQdia5v0wJ0Du8iASrnPznxk1XFz4zsFhtoIewlxqcmK+NRwFm
CIIZfb53tQ8bJZpCcuUVA75JFPMAHmiTkOUYN80LCDZiBlu59Z1bxRXeOEla42MI2Jjukf5eYvZu
faJ55qEMcMaVAkTKJ90RmEG7x1nko2lDhdMTOPwBVo8/AxbWq4uQFgzGVfzlGAtoUmtw5NBuLCyb
LUrlKKrQqb0usPPTZj6SuslmieO3HrW+eOaILEPfov7oBA6+/lRZ8o9+REK+BXozH6jWQE5Mq2Iu
f5C1N0S7HNWXJe5wb7vHNeWJaQQmPWe7a+5e70HZYRI/7/7bvNbnsWshy+/aWBRAkpudTnatac+i
aBlYYxbTQkvgC6Rb3LwGKRO7K9bl1SHhcPI4Hh7yNwRdObNpmZrp4uyR9SSuReUVyFXV1hNPI996
qzgZ3X19G8Xr2GIi2pG+AjVsC42FFqCdiiJ+YGOTC67UfqUxZVEgTmWJkvx12on+uadqFLPSMnl1
UtbUkdTPFv895GMJaCQ8Axqnj1WOm5KM7ry9u70kmRc6Rf+qB+VH6333Xjc142cmqOEYKzHYyy1V
tntWqftI1G5ANsiIl7pFfUNQZhq/q8rK9TliFUwVq1SOfTNBGkoiFHp199wfmBaaBNdVRQ3iymmw
VVYLdU5Fy8ceKb8+Oo8pGm/t7WPSw/a5jdhnWc9+8K0CKsJtr1Km+tigdJ/1ilsOuelZIjs2aXk4
u2UUsqyPPUQyP4CcR4+0ITjS3U9rSuWTFnmBEYdiSW7J2hQ6RqvceNcyzTRpKirb+0vKFzaZ2Svi
i8ohhseOwjUq4Bl6e+qX+GM2cDfZ8K/zcDLZGoe01BS6X0MsZhaxryZYW+ONCgSYZkLGQpWky7Kc
nE3bAHL5T6X4C1HMrgNC2a/YO8mlGuT/OVVSCNgvZTV8AvmUbjkyplOjl953nUsM2AV/Q4bGEqgR
rne7Rr2D6PuipgjL7Fh7DpwH7CJXiK0ZudoZ4KCBLkfxVh2C9X+hsplpYrd2J2sDtzbOZ1bIXvbY
eIoWn4ih42HzWpVms1Mtm6ebRiqTLGFZjR1+5xgXFWotMJtG2wAXC2DO31Lqkz86u9ZQYeM/5R/x
+bKZYB+MLtUqPX4ta0tT2VetqLFTEvQSF9A3zk9By8PgW8sYZKcCzLSAbYJFwf3CQVbMZ1Hjqfn2
pQEAGksBUYy6+qT1hptUuJv+v2nzxIdtCS2V1+q+ZQ144I+tjU1NaWsix0/aI+zMij/gWmrNiaGU
3M3etJZRHrsKBPUr/1dv3Cr+uR7yaMMPnS7o6infcWH0Pvq3SpLOKM/uV+2carZmseYcJun46EKA
m6eDyFyYf9Bofh19VqlcsKiqCVkzn2f9MdZgTFe3gaOrNpRhju1+ouVYjPxRILJLIxEIMo7Bka8U
VQfm/Mu27y9N26Jal6ne3pnIljLz3O57bnvq9PVRqzoSjouI0DsUkE0CDLpFXY0GYyFw4PyJ1E8I
yxMENMioxhOiwsO8Nc2KR72lFsTnMbhLyHy9IU2axRw2MxzxUP1PIAw0iL/lwvByQtc4jImoCwcY
DUY0uSP5Y62uPzlgkJTLGxb88eCB7XkIO2m/EfXqfLQoz6RvDN8tRf6ZJEe3GjK60RZ74W9VXdqi
TjFUCPGRYwjblvEPbOP2Hcwfx+EuxnyuRn1pl9HW6zIbmtEP2OnYLatryyYEmRcHNI2IyGFOo4Uu
yNi6CndWO74BldSXDit9xc858/icMyHvRGWUf+W0ScV+i12hPG7LmOAGb3830XkyoEXXb07Sgt4c
CWRTQ3JMzkdt7ZBFwsQVuLyxA3R54TOtYxycq25ImxU6a0QjpbpndLwCwgNntiqkTLW0La2+gSF4
fg5O2AdgI7F7QRk1pHDp2yag3j/wvIq5+Q/JL5OQXtLZdiDKXKXEj1Iz9hr9M8PsRoZ/+8Bilesy
BbzvsVPPzg/J9nSQjCIao+FSsKdxfjYVWWLWbt9lBnwIr6qdZi5RR67lVcgZy5COXKdOuT1vXv+5
uuIKX/fnWGrXENVDTyoW+Q1D43YXClMQAjyw/KqGU4ejtpuxA5YcWCCW1qwkUwumQdUlgsQOhaNA
DR0T6ZJARmUoPD0xUDByP6gjPus4ai7Z6j6K0/fu1cfhI/iXqNgEPwk6b+OQkPZtkLqkg7c4g8I4
yXR9btrQ20FiUIqBi/hNbJtXB0xHFEt/ZOOnxsVeoe5u+2+p6g+YB4VlsH1HVeDjO3TKfLKyJFkr
KqVgKu4gFIF+G+eKahT1PefT1fwdj+hcE8v+8kNNQpB4/tWuteseaYtDsxtv+Ot2nKesGD8SQLKf
pTIvrFnPCsLU59GSnNiVSxKO9XW4cg06Lf/n12Q/1qfqtWJJOuTPQKyBV6XoWr2MfykzWt3oK+n9
K/bsfkRfGNnPE03KwyjsvkkG9VMYWq2Kd0Ni5iSsxaQXJRM76WLfJf9SMtyHYrEhhO+rKd01J8Lh
l5ozbqkmKqb6GIwD3CWGfQxiHvJWfuWPOH3gG93txJ1S8CpKjQp6op3zNUajki106K0KICbNrWSe
QrbR6IR7/Mro+wmputm0JfvMWAor4d1Ilu0MyTJrUcMMASTr4n4BqUKQnNA8oaA7CDz+Bg3fMi67
7UqOW5XTj+vtPrUzW5wgrL4TFIMmLsB6L0EpjTCcp4zGS6hDjk61/oMdFXfbx4qSOHYbfhKTYO4y
5udNatfSy42xKRyA8D+mH1t1qdnMRUgeo9TrLYPm1h4JzXjjhfPIx/H8bp001qwXdDz4NroScImb
sTGnONqhCCF5id1z4YmW0U+sCU48wgzlKDQR+jhDILBqd6O9Fc9k4ki/tdKirq8wRUjLjwP7hkXC
mknQKR9j2LkmcO6Bwa8yKB2HmNX6c9OYY3xsGxylygQp7sA/RXQ9RMDSnvghrRIQILPyZLc2VrAp
9ReNVLyb1Fn4mgYOyUdQ7E0BNypcYyD0w49gLj9okVOXEKa9nPtC1gbOB3x+t62/rVn/eqRo4qiQ
SqOiSMa/YYWvIlSDs/gLpohaFVxwFRXR2c49IQU3UgEzJpY5x/iHHC29PFcbuTuUzCpb8tQ8KdH2
LR0m/RIcHbJwdbCK9OvTnnfL3oqeGWLgykuNkRVnYV6nsAxk74pz575JiCzBvnsixAUXKsINtkRl
rOBHWEdHgnYkok2tdG/mwnFv5+naFEd1s5HVsQN0Vnx4MeY1FPEDN/9pcAahShplli+XPsFEoUmA
I4P8IX0B3TNud8mdCJlsTHXsCxfe15MPKPMPEYWKwckxCngJ32eTOhCYN6+ZyVACS3hhQKGJi5K5
OoCG0kKXUcEe1ovA5/7wwt0z230LDb4SZsRdCV50Ftj91Es6aKLbIqeqoq0ASu1O5UTNAYZ88dsg
8XPHuAmtmyhGIuaatmbAcPOjAioqveffiDWrxveUrnfJjfkqTlNLrkLcO9m1KgQyd9elWfa3Xd9Y
Raan1f9tovWqcqE8bnOKz3iIU4f4dNXpYCjcsLMpEkQoa0QAOHVmECDHm1PgCymyxBGGhnecHkss
4zu3gQrXQp8PNpb55ukuh+YmFwaKuMhE59TmNwH20hcHNeEF2IS23GP//kdf4iFXV2++duvNpSKV
xP81lBGZRCX/NVi/borvCpGmuUrX/2X0RU1X0hDKb15WIAdk7GMD+4PrSJOnewVU7GdiXsM++4Nw
68rL56SA5kOTIk1kHd9ng8KCgZgpBaLV9TqxpGUPySwbMpV/SyLNHAaYJz8NcKkD8mpD4bTN3A6o
V6rtheSyq8QzECNSvPZH5xRi95fRyd73q2iUKKURlsgb/tNo5k4Nj7YgAmcigpmrmxAC3otojhT9
9h6N4cLmpNj3ex38t+dtX7+lSv3vOBrgutCoOnOBPXTvGlMeC0tkCCti9AI5CGp9vtSEURdbia+k
1uzT2TRkvdWWecqXazjb6TPp/ogTr+lA/5lQpPM1HK5ZycsMXv2tO3hVBHhBsIin+r87bfsLJMK/
vPvbUYtup+vJ/9GRXLE2TT7/fB4A/OkYfQt871QSKAlb2yY8oJN/TsVfTmpC3A7efJncuhQ6Cmlm
ULb2SielArqHUPbHcsRzXTIKQpRnDAcE8vI7qYx/ZrSqiMAi/fEV/C44EGx45ofUbMFallLpRHqI
J3SGJPz7Y4B71W2sr9OdPmz8axftKGMpTE4Ya7/0oTfDmVps6R+G4Mibv+910tCkIxH8lVKiSGkr
oCkpOZA2hQV/TcN1Z/oOJbtjMynsPL39+3GxLG7vddcFchXjeA7+UpPRTar5crplYcr1SBOmZDsL
ngsKRbFUAzLbrcxr50Q3pN3HezcxtDu/XbXBRDKsYaVT+D8TeppjwC3odEEEVU+tMuUiwhnOhimb
ct0B+IHW9xbCKHc//Fz4cMRDssSwake8yYW1IjfD6MkfLF9BAUdd43/Gbq9tjSs3Y7VdeS6udEE9
am8xTBjetfkfEswbb58Kq/QO45xnqeBjhANSKZI1C/AJVLMB6rBMCMtENnB3G++OrwHshCu+16L7
L7tlDNHP+GHwHEfV81sKpLI1kvoS+eRn4fd8iLkBZ44+Mm+X8OZi6ncY3atQ/o+f6ql/uoWUIDLD
dYuhXXk6huSyqQYQlY/ylKxUViVZPRfL6dpPIbQ4vHd/MY7CgcixWp7zs7geTPA1HTmBaJfn4dyY
chfUqYpB59GuRIuERpwqVEyceN4nB0bApxVOVW5kVUtHJAiwElMCCwu8u0im311BOGAkc3caeBNS
DcRzHfJH9f9HLn6EmSgR5To6L3TDsYwHW2MszjewI03FM3czC/2oLWGezW1Vha9plNS9dGa45vK6
QcNsuqL1wRY4+iI4Dxi/bxJjwQCGU942IxbLX2QIrlLfUM4XNlWWGMNBme0UI8CdK2GH4pFEpwen
OVI0A7PmRxDuMuok/k+cbRwtwr5nXBadB6XK89eLNrbHtCUDWL/CdxRny/TRal3dtcEoudVOlUyN
FkZxkIvC3Cl7KyGTs3szkHT0wEy4cOMrlPlEttJ/kR4Zr7Xsiea/QqiMhytxvSnBC889Oz6/IJnw
8rt3Bt7LAXzzfo3Sn7VKeKCby7RAey+ejHhRm/szt7mVqvKmC3yM7PKU+1+4jxIuvTTjujovu7UI
Si0P/EOnYH1Ht1ZQRaFsTj3SNzMaN9PwdqUv5/SzIPEp0UToAzc+MUHj2pHOa4Rckz/h/VxDz5z8
dM4OaEoqXrdTDtYONHP11eigMQk/FTGsrx0yFaiXWbWY4DIcznaJ7HM0xMomCE0g0U4+Lb5H1khg
hJujsHr/xCL/Dyz1LRP9EB8nnHHaPxJvAtHyzQxqUsnUS0GBSH8u4AapTjrQkkkAbSvAXaJa1ufI
Yh+X/8093001jmKgmjZ67C0rQY6foMAX3jkCCP3b20AgYht5jn0fX+WwTm62dw+VQqugeVSDLXgs
Jfnqn25fTkh5KaYKKUM6hOsMilt2MWsb74DMBQJjnr7iFIt/CkHTh6TKWKbsNNZVCHjfApkJPeE/
aFR7I8hxsv4faw1D9Ttv6ANPl62Taf7wqKcFbJxESxoYmXsW3tCYKvwymSug3v2cRgeo3LV3hX4M
nfjiPzaMKzGvMNfw6TpL73th5uNnPdumbpHt6W1vdGIFs7CcJrnoxQqbnDIZWyv/3/sr1uz2a3+M
fGNgfZdTuCBpdvh15q0q7blbkCpFOK1Ixi37HKEupZsO/pcJratLrKIvKhsIzZVO5LOwqRaoxM3b
z6VdYaxSSaHRYuCTVthW0Xva5UOAqebDkVayXbix8+K64daw+f4pXeIdbuzWEYRd3zKUPxN+MXlo
3oHKy3S1xI9Rl6gb9zzEIbCqUbUJ6XzRpY3BxMCeHXOYAQbU2yu9qmK/ec15ii3ldpJW7QQeZVNq
O2VlunFvj35ZY5Qrfe2c7JhPg2wTv9ffXn1c3p5u6HSrNPYJESlufEAJJ/e2wcp1kONY3NlY/P4x
/qSV2+invBjvJNnUIyYebfsrWU2cjgtpPHQP14q4XmrRf4ys2bMmaiWprSf1mHd8zRwnBs8jJXNI
jTbifULEOXgLadAx46g37Mi3tXjF2StRwlSNEFmolARx9rmVmDpSqI7hjn7PfpIlK2w7BfO9+3os
QBvais0Gxxc9hB61I3JJ4GkU/MCgnBaqxxRtOc/LWz/zvOIh72sKjAzpCRMv+38qm1YZ68u2o2tu
3FLrBwO+q+giIdZh0BCx6M6SqvKe24Kyq+3br0d2QE8Qnh5jlMvnOyi0qNVSwFGYr/H9rx8hiT3o
Ay2Ot12jcnlOly4jCDe08R/4Rd1m6rthlAVJRZrVWSTTQV402g5rsBKyLNGJmSi/lEJMrPErG42u
Uz3ciX9aqUbd90KfucHA6KdH/3yMkR3JSlGoulRsmOFEFxHmavxijNfdPODQ1zTnvFFleQF2cgd8
iB0tQU/zUXxSjUot0+dR8WdoYwMPYGNVLHUAjAITaQX9uDv6Ck4h6uM99szLhkDN+GS6yOl5D+eg
LKn5Vwf00RW5d+WBoUtI2Xp4kDQbO/HObPgUaTap5anaqKrOFEKJdzkH8fQtdMHLKmjvcMWoMY9N
b50GFlRt5CyEzLTDcy54aE0TpuXUolcuBtbYWUXOAPJruxAEqZIHccojlC/onDzHcK/AZYlDx3iq
IRwBwZkJbVwMco3NPNMm0QyHCsgg3xLkKaP1q5M+HMJP8DVEXgc1KSWHHHF3tQVJMO9hCQiU9h9N
L3SWY0IxBNepha0eNou8xjTtousxXlMBD5NbsMkccSZvukdFZDDz8anG66xlrnzPpQL3xk0y/taf
XY2CMGFckTJ1w4z4mwY8GJ1+1rINO0MMVgFRyV1eT3MmBjC5oiwNLkkZlAudYwIyWKvgjj49GGlJ
7R9XNa9Nl14rSAO4dPAkZk5xgij5HmTQVLVttjnDSOK2eXPDN29FA6E790L6cnajic8dxhaGo7WV
syhcouF7oanIM0pGjUhnNPys/Gh+9JAdNiy9hz90tJzJ8HVaawzCN5myzP++l1M6iFDhw1vbpcp0
BHCfjiCibCQk9z0kXxXastWJbo1H6ZVny4umX9JxJrrJw3IskdNkCUkBz1LK8Z8ItyxdGNtgorRJ
cM0BdvvPxbrAZIiWzOwZxQhp4fd9hRcDsLtdmyP2u66YiraAyKvOjWZBIU1UrNNags1wNUncvuDF
CW9OIFIMMM9uqVg7yGbMOOe1BjPCWCt6/BmTzWYokkaeJpOdjGlDg+bSrz7e0wnPKO7byNFiV278
Y7olLBDBKaoIhnn9N8lYSk9w1OO0NSlFaUOqsbydvcP8t3c4NtVwecl9iK6X/vhig+NONMCTxOzc
Dg6iw0aEpFli/CrLdEHubFrQqOteZyqbRStz9yMd1fZxf0hDzADQXPb7dBPf7vTbyXQT7cvsDGG1
fQNKnGM4sW0P4alijdLMqNWLSQHbbC8sIgAyIQ9hwZO2jDXP2610ZxVSxxMuD8N4IBGppuKa4L1j
qlRECD/XGuQJRT6hGJTbTiQFSjYrlWGp6wlffX4q+8GbcERgizxna0sPyGJ6zswg5q7EzV7Wz5Xg
T9OHjMknNAEu0tliW/bB3kjGu5JtrOsqUpSZyWABsowWd4+VEArHuyAG/7iWpqoYW0ugF7Uw5GfN
lMgZEJO4FOxtXNnGv/6VuPHetzE+ekVxIDvJPF1HNOqlbKnEAVMrvXN7inrFQeBZloqgGy3C7ASH
iKxQcp9FyPRbU1cOHO3thNfaOYx+07SB375It7GAOrR3lBxKVDgTLcfHpsFRbO7Kz5ebvRNoo1K+
xu8htRrkZjRfG13mZNlTcyg+RkkBYTgeBtbtIQEgDk8v1fTcSr0U5cNoI8p3j+ZwZ/rOTX5I6Bn/
FcVwjE+ESeaSybFcqBCB5o59NG3Hydeo+7ASQqs1ZQqNF4ULpvwxLnOZ5WjjYP+aXa7wowbw9SUc
eM+NSz9fvSxm8TqVqXjz29qv0l7LlM0ynrVxZy3uwTHCQR9JtlYjWkVHWem1pLhi2Op8sk8TXO+N
KSVCgpHpax50FMjfFhboYbKZ8ZiSdBEQ7iguei8FZLCxsGazw82pe5sps98Zm4KGBJKRg5n+OvWO
fIwjK6HaXeU5sbMeUJUSEX7XdZnWwUJoFa48bJsO8D4QqfGQ09VU7KAkDvO+u6IK7Wr8MHycZMJs
QsMVuJuu9Oa6udle4r2O8TEMq8f30OGttI55KKJPHCMRBEZY48gvh2vYabzM3yR4KAm1RW71S2AR
fWcovoptcX/wU9/p0FxzvCaXNUvoFYXAstV+HVg2OxaYqRVyspe7PqEuI7a6+BtYqcCPKGoEGwYH
y84f/9vgdrLIvBPRwjo6uMwtjWN7e+nKLu+S/5AbmoCLOD0BO6YGkjjDDm1SIPtGSVAUVMV2FvkW
8vK2ti62NLwE0EjBEm/DANbiX8WK5KRtvhUWVvvNJie/Pq6o6bdHOvQBosjoH3AI76Nfq4QL91xf
DEC35HEnQugsRLV3sbJ7xhOcHnQp1DSUqthNvJSGZ8AMTNGay7zXgAvk1oy2IwjvgEHrdHas71ja
LseiN4DkUkG2wl6UP0OGzTHyJil3Af1lzTGGuCtOHW07Vh4qbaB8FPJ9cA4edpQIw8DyQ/Fm9PQO
OQa4/qMNT4CQLoCJMPaK/nOL6GtM9BP0EkfnBHVqdADn2ZPquI+4eh7qWzQQrp0jNZiD2SuYs/EF
5TSTrFzRHF7YwrpmvwT4DpgngTsrDNnZCsfQor0h3CIt1HZoEREZ3e2x1fMOujpe49QzYkN2Qld0
IZnvEci/b+9FLCY/0DPnBFcZLfzq1rC7CFi66g1jmPjJ3ZQMiCKuxNg6RTFWxg5AgNMBuSLdMN4y
s38mgxJpyGsQfNBwtnLLq2AqywR7xSsgAgK31sbGJRIQ07/pFAbYN5Xn9Y8MsY77vA8Z2XLDn1Dz
/2UYUrbTyoNxjQRWUJUioaS/xphxGJP+XiPlkSmbK19I6Woe6ufLLhExuitM+K2dWRsQvTGlQvA4
Z8f6kNUo6zSeKH5E4+cl4PWjPzt1C9X/dxra5Q6Ahc9VjS3PwfdU6rA+S2Jgi9TXrrHBaO87oreS
eK5GQ3rCg1A/l8PPfXaM6BekWoEytL2KfVxKaYNQEQ0ONY0ulc85zARdQnUy3gSvPUqgosMnpNN8
B2gMUO+FWgyEOSjoVVHkNMIKI317cXsUf5pwgQl0JGD5gIXBCMvH62XnWXCdsMshZWKFCyye+Fr2
SJmbKnVAkRN9nXjGF7ynskJOUTOKocl65qw8oFjjID7v6eGP5m2l/mNAefyZHRL32fpCPqEBi/9C
trbDFSBzRh8sFwI35cijRnm3cE7ZAne0bzKqKng6PvWgd96EYAzX6pxiXduh4kV4dofA2ItUk+Qh
m+IuUCRnumURKoMA7OuIO2s3tM1N5bXj458ykWap7byN5MhmFH5+Vp/wWum5B1cLOG9Uw0ykLQ69
25tuTD200ag16OQbsGCwrdTW4sS9QkVghNf13tL9XlL2mY666QkpEIs08tBw0EPxh1Yt0hRctr7d
t3UdL23D1PlfBgHwlmDcBOgix83TxQqusuvoEYRg626NoD7hhJ3uAVnLdn75Kl+DSMDfXmYXcGht
4IZ2P9afwcBDPQ91JjOc6CArh0RnmdXFro6GUVofVwaP+Mxou5b7s12Qa26M0CicYWAloUJUA3cy
SUH85lF6/coJmmvWyfSksS8rpax1n7YTkcawUfXQd2AdpHNxT6GDMGlbyeHy4MO/HEWPhcwo4enL
hDoBJZ7MUEGkMV/El3KhbZKtspLU9u21i0YYWsjCtgEscN04BZbP9D9CT5k1Eo4e5f+AvzZkyYqO
UV+z/SA6ZTTj+zvBfEkwD6wqJnebh6JhUl8wvDGlEVRPMwbkpXy1bLXqivFN/fxgipI4piELKzNL
+u0r8H/5vfaYDh8+93ltJeu1xY9J7ZiPD93XsR50sHgogpx7YGLcQx88pE/CeI1MgQHiUItjUfct
2j00+DAPPtmVSSc6EskPKQJGuKlblrveIFFM7IJt8ZDXfDXOtoOOpW2pTLb928kT5ehNEkN7tKwQ
KOfwKV5/jcKotlXPC+Sbi1ChRobO+pNUkiBlQXCwz4ofap3HSRfynatT0IdEu5Rq8Z9scjgD8lli
FZlCXdai/3pVB5gsrunuhddfJXLKJ0LLLPEGODTipDh3UqQHlEqo8diGjYOTN3pk5OfZImVvUFw4
Zdg5Mk+R6nurG/LsOgPsQb56lzessNQ+uWZmDU6G7kKJMCJEuS5eFDD6GFrAdiMLVHH+iF6bLTUx
b/p08AzU6TUbPo1KDjxzrUUrcGchJPqqHe0yeGLwzqRCmphQNe1w27TMlrfy/312w2yZlQ+vdAq7
TLn5oR6qTmuM9+MCFe9PxKtIt/FZOQ913mhsZ+R7bFy9OrfqeNLR2V7yW872et9995bhzupd2vgs
fpoKoOvqAO8Txj7M7Lnjy+wHA8r2A5uYWZh6c5CM6OBxDbepMdqSdLSbVkNjjUch9PMpbkSEe/IE
Ce54a9fdb/Fjoc9AHjBe92dNQT/bd69HE3z+mptoqnzyu6oqha4ASWhzudw3rAuBbKmDIkHjBGFw
HD6H1WJXuWF4mhpuPuFctFdaKlsWcc4eohAIQjCcafS8KHNWEIL4TXSSKQwU6oh/IrFO7cqnWTaU
OqRFwya9ELHdthMdcwZftv9Kk4+Fq/80Heeh6z7vGr/g6/DbO95kls7QHu0q0kP4+owCWrYGl6WG
4YNaraylW5ImDWktFIolLGeCEA6GXq506AjjmWuibqiRZUsbhU841u6ds7wscutwc+Q2e/qXT8p6
enaqTznhKzEEFUdOi/s/YAf3YM0iTk2CLY0rcRJl9oGZB6KeJBWt9hOcZucsS8xXv15IMTU4IwWf
SrZUe5rLvWxPA/h+ZByHKHI9m+3q6Sjhq32MvIvRpsBbnmHFyHCVQV5+ZXrmMhFy6+1r2r6X8I4H
y0csTCwz46wJy0vRgJPxeZBXGwjKWwEvDf+t6HvHtlU35zgpcDGSHzdZnd/8zVpf2VSLYTeHb00t
JU5A0skBjmNN9bRzctli+AwJjsV8J6AzPIi7E4BvvcjGUULxfF5EQJVw5jZ7h0eeth9RvrM8Vcbu
yLXXXSfKEpZ8qOaiucIDCVyPB8Xyok8cKtcazQjFDjD2443LVlP3B0ELgs3maVPbNBJ+sKLSGBhL
yq4paSeBDUlD8w42Zc/bI5xnHsLtKOKvy0gnIpBR59ubvdGF+WbtdsV00HpbPQJrqQDs09+7k5hv
xxcs64er6ATKw2ieLYTjggBX7orn89w5QPkXUjNx5ooXmPMRKiMeQKnR7XHIT9iI82PMIKHoCtQk
eqWtMypT1cZ9XZDdsx/czp9MxMF25eIbqwwF7c0GbqMUpHNh/QHzWCNGWTrUkd49+w9cxVQR+hKI
r4TDvkTiBwEiKIfs5zQ8Nz6jP7WiO3nJhtgEJ2MvttskbQzdVbyl5qFO6Nhyzc06MyY7q9FBLkEe
qSmNteGJMH9g6qUnADbQTKXiO6BqtYeWoUtODYlnp+PjFwzOA9IoVCZ095l2rebecPVo/q1Nq9RL
tcHh+pDJPgCPMgLQaEtqYC6UQnKbUU2h6WWVpKqCRfP082lGitpVu+iYXA25EXIe3TTPSYBBLB1O
p0IvyrcStBiKpIe7LUZ4F9NzLQNApGqYJXasrFCVDMS6FIDMRdl5Pv7sNWbdvLBTBn1+Wo8Mpbfp
PwXPBcCQQs6mRGaO4Ada58Q+90JkbqmwKtswCuHitGFT0UkPYRj4u6wM63smr89FbJhhecj7MiC3
89d95LKq2IsSyeGvpNO+kQF21lIcxCRcuBTvU087ChD/8QsiKESVAcr6QajYeeS0W3nWBG3ECrv3
TYGt2LtUPTx9cfDq7Z5q5CriL9k1PdWp+oo/DduSuxgkE/VcQ8wANkpoAIetxWj10A+xc5Fpd68c
vJ6nS4riMpIBvcRxTyh91U0c351ZxtR7BaB1rkxjWcbC4w29b+XBkm0BtiHlKxagsoINIj6Qry4h
aNVJjpuSmmcSRyArFeqMXMWum2coCQSinwa8VO+ItsPhN2QvlaTlbXWKhpMLXkrIMDw5mteX20qq
e5uo2OxdYTS6vIoQHIsDGIglDOVw8x6hvh780LCJQQpzKDSmUAnM4/AQe1W/NgyYQ4/Xnd/SWmuT
NNRctdnp+mVfb6uMWgRxPEu8HVBPHdXm5K6djla7rwvYRQQlOBOdNeLkY8XS8Bbhqcsf+Hq9CKly
0KapVw9PFHVTTqt2Vm6qj+WvBWzL0Hvjz8sLZ3WXU13zq7Tyw1AUjaXSEt1aaWsHQj4gNcawoH46
8RHArmTeHluoG2LvRoWJSUF7lBKUBYvrQCytMsVEIzXq4yNLf+RXXILBqT6k3SrTVBOi4nP1A1V5
90C3L9QSkus8as4dimxfI0HQS0qwmnVoIxhh0C0pRiv5dydgfBXQtYikLu2NCP5NkRJ+vUSzbJa+
hvIhV/gnyUp17IABzzY+UgkyzXlqwQo65B1ccJ09cSnCvv3D6D7x7ExLnRjwrKW5iM8F6N28OVsF
9Ynrl4fAw/DPTgURpqKwUj/kx5ARjjVh2t2JpEW2makOAvdORWdZmQwjYsS7ovUg8OD3EltR12GU
ftHgXyeKi+e1xQRk5ew0rr5D9HjODHy/Lb550FHZgx64rUAMCrOQWZziPrIXP/WfVTmNP69SdB8R
l3i6zlyxssDPA5ThQAQHCLI9yuyKiN6nY1SZx8YF64Bu6YglrIpQiZ/X4tbwk+5znaXP9K6Vt7qR
w1VdpxyfP/xrdHJ4RuRyceDyFZzLmlzT/M9F9/RAMm/KQqKdW81bjtbJ7tJO/k0yDeMLVU+yT7Jf
QCz+2233aZP/kqmid6QZ5Dz7rvrHNRDlemRe8C8l2Dp/lWX4Cccw/b+lficRIRY6DbrkEfukpasf
Xz9PPWvjF4Sx+D9DON5lwVpbDv/n502DaPWAPJ/7rAgHmzjvD29WkXVhbFvX6xgyYs76pdxsuQgI
RiykVHOCPkvLoTJOmtv41kvLQIL07xdyR6a8RZtRk6Y9pnKzpF9JH5bzFFB/mbH5RufCI6ViVKmJ
XhO8bjd90feS/euuGKUkcAa4h2eWwnduHYnvnsqpIN5rfnvEV8JIFwm7G1roD8pd7tPD6Z1gB8pp
xDBcjP7lX2lQ2va234eZ1Zf8IItYcqs6J/w/cJw9fCP37Cv50w/0xdRMu1IIrWRYg7K6ksREXI7V
UitFD2m9zcN1Ydm83V25Cm2bwGq1+seSiBdYsXp9M//kmtNS/UOMOXu/olTQEz6QtSdpxt1GmN1r
h/5p2nxlw8YCFnrXF8/pjatScmQR/ULhYsUFHBUIKrzhL+o098F+RAfZAbWiOun/j7rYsKRGtHj6
tA9P0Md7Qi7uiGlGlWqBUqhGSipmzuDvmAdhogRC4U+lg8uE+ArODbnSKALD01KX80pfSVnSO+p4
ztEmWvx/1XXnRKzqnUJEA43UZNLg5idth1QSWvsI6QVmtGSwFncTFbf5cS43vL3wETfKMrno8wSt
8QDm6DQxvfAzrK00ZJHwCOZi9NSaLF612UDTQ5mPSKIZtsYju8CuIS9++cy3GGmYYSHBSDrF82Q1
yc2cThM8zfXKOloeFm3DZQLNyySeHZAChsh+ujqm33bdlzLTlMrPMHkgISjNFAnQiyYRex5ApED3
hOYP1TW9zvJ8/GrDEYYR4PvVG8aboZ+pGL50sElTFoKGydFNOW6rJOQN2PkbRFIRL/fw/WKSXfFF
Nv2B+1UO5sPApalYZQQym1aPglEpGuGUwwptcGj1ZroCLTKTKUYQY/oGRgoR1aXLGH6BqgNneNns
wEJfmo8qw1GLICxEL70smDFKHeSX7WNIzoXfDXIwVBZs75fqyvdZlHHION0crzImT3fG9onxLs3S
N2wjhZGQiaZqXeeCgKiXxtJaGZMJ0VgvLOsv1UWTzBBVXmVRSqk0jhI2T5bzpuVzbOLopBX0tKfG
zEj/oWTjHCw2li9glUO9bTdslna/uUpjcKKXq0BdEdwA0tfUpdth2kRTWdK4CYEHkFYIbm/BNc95
RLVgiFM7c577uYmBISro8ZGY2h8hXXzj1iZOYofaHKTySrV1OtHYT2KW5nQsgCZQBkhklWIdHlaW
OJrnOiF6Lp8llSUe0p2efGxjYpOn/3dBs4CDPHGcTWyWCJxNyXKdcMvPgnwhImazjsz7F01musTo
CP/Dz2IUCi3FlSsybSRbKLgMEBS20ci8pjGa+liYC8nc9iZPxt5+rz4aFXsvZ1mrvrIvyVA3hkBb
H3d15cAESltBUzsg1aiNEm827YnJTLvK2QrE8mpmqkbY/1ex2vIN3o/WXuOrei9lF6sYoV9Fqdin
CQhFfvOoGC+LITBzvLAasGTHZSvpsAF/8qPUAqkoPRl0Q8pLB0TlKND7Xvju8cqKI8MSts4YDEHx
HUCVc08D8HOkw7IXEbUup4j1WwF2DW2h+b3KdQKtDxH2+SBkPIsT9jHh5PQKxrNLkg1wQQms0HtZ
AP7dmjYMWYDCIGbiDxtInBG/Ezt2U1HBTBYGiOz4dX99TKoc+NwBwp/gm2XRO2TMaTzn0OhNm77M
RURwKnCyixEYIfzN5A7kuw3l59JzegL7e58LniztmLPpvfb0ANjYEoDQhQUiQFsG4QCyJCKCLXQ+
Y8sbk2lro54zeN3feHXI4MwBZ5rVRTqDkraRfqHB2ugrFBJ0OyyltrFIJJUWaoLMas4SQSC+sa9P
gg6K94eZ7CMvWjMYX9jsHsGrG4qqqpE2CpBh8dEht0jJ+3B8dwOoDQWszIlNsTpEMoRVecu2w4Gm
86NFOUyUZC9oJyrCNo0LiGDscyh0KKKArxn/BZBdLVWVZHY8/s9b1Yl0E4DgK3Iha/2IkdDpZHKb
efbErAExbxrIgpltEpJ1V65kOlyaPBemBKYA3Jhuoo5vy3mCfjo2Cn43hJ0gk4yWRkF8zZx79jvh
QymkaDRjNyyvCuUoiiw8ZKXFoN35kCFBn2UVtdy9Xca1jMQfGArbyGhd+aVmVgrJ6b3jDxeocqrC
EAO7y3ub4AXkRUoLiZUjHy7ln+bIInO/xN8H0zCzN4kcDYZDurLapK8mlqDcOsqj7A2Oytv6Tx+x
QymDqGD6W7pb/BRd0C5hQy2Whrfwy4mBl2KWg84qkitRg7L4B49fQomA+Ld4H6EqDdho7AjNT6ZZ
Mbee3NEpDt6ui+cFHBm+qTZY9PFN9SN0fLAh7X0tz5994NesYioanX/wmvmv8LBnOVGGVBsKszjV
Dw9DDYhpnK+KNtFHFi+Nb917fkuVaL5zuCtN29OKBpIRBtkEqZJx2pYeglpanMbErd6LmYyM0Ri5
q6Gx8J7+E/fBcz0clkKnR3M0el/PxYh7Zz6HcyE01/kQC6doBiJg7RyKcRqachCieNHw8SM/qnwb
iKx8QQ/CuC2Op/YdRgzj9WPa6TArKHkYe1sdIXjN3+YaTCtF3egm+VojKzNUuGPnYAI1Ar7Pp/Ye
TFgFJn1ulqsje93SxYe6+swGQhNuA1WEZUHkFHhD0o793hn2P7GnthouqR+WGqeWluQW3G5Zfn1o
4t4NTdLuIwEGHPj9c1a4KGw9dmDOzzopuv4w/v4hCOjTvL3QYkzizse9wDRDN+eEe3rx/li6MaGo
3qMRBqztaqfKs+AOZX+NGJtA8br6Ax6EApodZGOgdb/Kdx+Kc4TTcxvVWYrpaicug3pWBgtaNCyA
nf/422HWiAMIDcb9TI4ks3RFWT/0Wjc4bUBZkwkAyW5prKoKgGBBaWntCjF+AsUEFkJ2Vl8N83H3
kRf4DgTgW1utY1mfnc2dY6KtA+L2If5TyvUK4cAGElENWeio1ce8Klujr/Cuay82dAF3IapViHLK
eSbvIoXiSxXcAb8ajfAAhbxDt7rDhMQZXXTnq8j1TvuX2ky/IMci7emKbs7vp6dOqm47zE1di0lT
CmAAWBdA52nn6KiXcLc1TeezegMS/aD56pu19f1VWzGbM092oJ2ribFEpMfoP4Oe2rlUwcFjXdxz
mifoO4CY9VqZ3HCaJJ445h2xr8Hbd/vzJlahJE2jg8bIzNmLvQF+A1Za3fOvmxAmpi2vcYF4RuWm
qq9neow0RfJiO44a7HpLfj4nvYr0ymbpngkYNQJMoouM2ZsICmv+VVSq+Ldoz0gagh5HIwbCIa5x
OaMIqqOAJeZirhhDFnCEEqI7bkUTjQeM8tk8A0/bUl+SCc+m+lXkF64YMRbLj3K9VRQoCgWzm2wj
a9vdOI5YrY0RbrhFTqOM9fA1l0SrWrwg8RSXutvzdxubwP4hUpdxAamIESzdQ0ega5IPXQ0+NGVT
4HY1yi2/F/9kkYXSh4gTy5BoTUL9aPHVEObm2IOeC+Kk9tqEynfhYypAGeNoMgmmo4Ktm9YkIisk
dCe9WiznugbQEQeGCBg7NaJh5+24LO9QjjccL67gE3BqI6damsTEG9ZvKZpkLxIor9iTTYMWtU6R
ZBHgeA+n0xNH5Y+2OKSwcfrP6hJL87XNrm/4iC5EyaEpGbHZXAksFp37LBL+mKs638TT25+07veJ
M7jbTr2TtJqswIPUmlcgGXLG3tU7MtTrD3ewj5yKtC61F8PXfrRlzaP38Wc4tx7+4Dl3fYyqg7EL
cIcoFN+vxsnmrvL+kvL13BlHoVAlEnp2mJ+tiFOXxJuxHxuF6Xx1CPoTsT0ukNAqrcxyQuKei22J
OZKi4r7ajibJkajaaCbEsABgEqKe4OAVkT1958uNWLXRXtFgXVXdynFckaaSn1nykoREJix/1WF7
6ihnfBLJjXHfoyPchO71msrDiYN4YmgzX4n3sozB2dHDSM9Up9W5hiwztHX6wzflZG9OeK5wdOQb
EerL1i6AMdeBQdKHv29Tih63KeepP/Ud+mAyNjvh+4SezIXqjO8SanSdh2CbmN8v97dJCU+hc9f0
wiu5o1x0K/gE5uU20VgM+ePhsEoTNRPuuwQ1yOWJ4rzJr1HtAG3TJUvVLerLobP7BtmkRnRpREdh
tqWoHwQADRonD2VAKpyn4hnYGidK/3a1m/cRMF6DcInZKtjxbFfLQoW7kBBQU4Plcmm62UpsiHKk
bqFcyAny/LfVzQEW0YRTeGC5vl0EWU7sRT7CUMlJM5DLQxIz74VARXp64SvQtMMmvBax39oX9hZA
T79dpR+hIrUy/1dBSrbdK01raLS93Xhty2645jWwTP7/eodRJnUHACw4M+6/os9zNFTBBpWccKRY
XY7y5gsMpvZHcQS8M6qK5bSxRE2qKDPe9AShQX/UagQVFMrXxvBbGs3mKwO8wYF6oESIrTmNLNEd
hlHjM2o8CnfFjiJPynQCRvIFRkXxUWVP6zCZfQHSBS/XPS5JhqT9fEvLlt4eyY4u+NpD/VyVeV5v
JSxhPC5Ggv0B4+ZD4YTvuUigYJxbRDszUT90FBUC4GWIOucpHuQFSVH1IsOrShazYnawtIVh8m1k
wdfd5l8+K7GV3Nl+0fekU1LRvRXO3/dqBq38z//gQViVcJF4hKX2q1ejdj7OJkNaWAdzdm1GTDkB
4fxToZ4iaTJBusmBdPVld6mCkHa7ciOiPZd47dSiwE/EBGIxu2xd75BeAGHc+nVIYLKlF65Nnped
UzfkOaj3ax2RpfyI+9inLDfBXpFt48gYMdFKdqD+tIK8a3YZ+glEZBF/mBp1r6mUrw+9AGYiCy8W
4j9by46Y27JzCCybYgha87rlI9b82MkQnxUOddLHqOtBm/yja2gK+7Qo0c7qofi2hs0HmRY2xbVP
zwSY6fUlX23rBI9D0LqGa5e9usxrEaVEbsrc17ZV0xOyrw+UTSqtfAQPeIEpeQhcizJ9guNNRdHb
gX9mvFrCp2roPjcPgbWb5njrKkdDt8IflIVs9zMlByCkUjCJz50N2pYs0ZJGhAnygtGsqnzzSnhA
dp5ZwBwbF5oShEkUscEujwhS2OhlwFXW+bexvS2XcI77c5xkv8csMImmR0mMqyygVNyjEVczlDEO
WmB7ATSmFw+BA8EFN9eaTCC6cOw1QwiAYr1khboWQOZ1FmRaUP2+Cghh85QQhAUPsI30qB0QkLob
UnGMQBh10wynnuJ73xoGGukuB9MVsqTrjdFa2Pgzwx9D0MNKSZcL442O5RsD+tmg+dbQ2QybryzY
jYbrUfEWXxMe5KEm0Cuv3vD/Gtizbj4sIZGE95FzXT3j6YBMis/5EXEzYHIT1rsEO27hhZAWeRW4
OHZM/2jk0GQFtaRa/WuMOAntXpCYcD50jL6rjZNMYnsWt8PQTpLmv97vNBqHIqzPzNnhaEeg2UHr
2kud9ykGWd8RT9gh7Kmir0BKltA8p0kajwORm9Y8aqbrZW6wpQ8MR2KH2UIcMTm61TKLenggXtin
kfuNBnFxJc7rfgz+rCi6q77c2LOv1GCTnSpNcXC79rjf1amnrsaPudqTm76q/RIuXLEY/CE1MguV
8/K4UFscbeMYGfgnctIYLIUqRBFxgE1gpxElpm2Wyatozeg+Cxl1udQwD2lRQn/6XlOUdOsDKQgQ
Rkft8F+Fo2rGALAEYECitd/Fx9l3q5X1gFnQ58Yw9w8wTI2gcvHw2vUGdysvfiRGEoaC/DsRhXy/
w5rEFYN19nLJ2gMB2a/bot0B7u47lee6kHWlS4Z0wIDUmaWehgVg1oG3YbqNPdlTkn2kB+Q1NEEI
DvPbFLPOWGt5aPkZ5q9YDKmb0NhJjP+3apeMbeqD7o03LF+dGdOyZATYe/DLue7902pMgEQB+bnD
NNOGlUNVDA0DC6fAdlKeLeOi56uuITrrhEEJWUaLUtAcHiKPjH+2Mr7+q6RK4vIvU3LbdxaX8wHB
xOAKH+oGd7AW0cxNeXKL7bcfaJLhhl1k9uGzw+KWvR2d4ac7g+utWbSae+pnyNQYkPQqnmBdtkOp
J2ZAZJFcFVuISwM7TWE3tHf8Lc0btxLhHi2n99AoiNQPoHmkQ3h62GQ0EWsgs4RubdByjuGE9kNa
q0l7HGTln+gDMCeO9KAD+aCgmjy3d4SAmIGS05qj/wapkCsYKblP5xYRppozhbl3E1Yxuu8JEoHy
fzHbbc+k6XoWyTyalBaBhyEJUTRJ+AxrbLtY1geNStKW3tLYQHURc/VbbkcI8dIBnKnkiYJI+Uyr
zm9V7AHK7tUINaxUT+WYC9sZ3GcEtzoP/RAvaWgUZ2dzPzkgTXSlmfr07PVtrM/0bFcv5S948crO
TftNc0R+gZiSpJ4en2165wzJKlJdiN75Z7RDp9sFdbSYjeRztobm4lu8wfLRXbUlBz0bgEqOsuWs
LDkoIWaOQ1+EhJSjlBIhJAaJaKSk2n8v4jpuniRYb//NU7/xmuBzQNklOjw+7olFxiJ4N5+QGNiT
Oadz54XiYwrNK3Qr+jSPJYUmrRWsdHUo8p78XqsPrszlU3Po8WZ5ApmD9NNpZvDaWFi9z+gMmTsI
lx7rHtYjRI/cNYxdndzXilMpnmamiqyKtBubbM3MZdjHnJjC/UZGt8uabZxzrm4X8OQvheoo/yZv
GJw1J5ri2mDwPqhQdVLdMmsOLYIDd0V9SNQpF4MTqagB4ebBJikU1mr08ZO8dys1mD+hNYb8x+WB
8yUmip0lkz1lbUGMAfRoMg/hDRIuokUerqtBWGWFi2aBQHdfBGrx5hI4q04eNLAqAdt9QR7SKtat
6f7pE14d3LN6p9FClyK8T4t18fH10RIxNvWSzf9VbjVFvWmOcuKycJ2j1fpwBo7M2dPd3Un2QhF1
JfLeHxRN7eAZMpq/mZr7ufxXLSIC7BtQ8t9gq+hoIaJVFEkx0n+oLb19g6ul3VP9oiHhHEDd/w8O
Q86j/7IghUICchOEE0HtGSj3XcC99n1BEb8pEydr/tklGkhcsnXJhcXwWzXCwCrnCaOYE7ZL8Rly
640AUM/+cysdm3vcSf+4JfBFci6R8S8yEE0g7szBQdr4MuIFz26gfF3VGbz5LPgc+UKR5CqWB++B
tdCpDFzeOrWkQEl8mptaGnCqilM7XAUUhuP2SFgUFXCGoIHMQVD612untR1Z+Y8wKEjcplad38kp
OWb7o7et2HZqX6t7UD+9pOCZInwtvbk13WKZ/lAJ/rwhc7+JlXTa02eEwp5cQekcw6uouHr4yjHq
sdmWXE2ezX1jugxzaqMNZj02i3O8JfwnxyItRdpQC6u9ECx9mCBiqwUihyLUmEDrEWGI/yRO5b84
9okuF1x2lnS2dxBmbX43IghFuWC7Lj00Un5Mt124Cu9qk4/dRBfWaCUFCe9An8D8FiVc1Xiubqdr
WVVlGkzxK+PyEeUvih1aPVkav4zZW9lyIXNuO+TLUpC2G66k56bFoksm6/zCiN2gFHksbgVrSY0+
EE4TTGHEGzFMOFy0eiVcaXhG1791oLC5ihq8Qv+/j8phKSTzqgMsH837Ucm1q+6RKVrsYbUMmU2I
RAr2Haf9zScjRcle4V0m5qoYY//mmm9+UDiQXySdwwRO3eJjazY4R78jteSKfSwojqYB9Nm3w29V
XFjqQJgM8if68tgHdUirMU73zIQXdf+Ft8uX2TMv1ykNDQYopMpHqZa6PfSERCBnMG63wF8RD+pE
/k8ICA8wMnOFRVwZR2xsRb4dFpiHKP1b3C94OkMfhMV1+IMxAL8+Xu1LRf167HqbkVIC2bS235oG
/9pIXRKbQCRoUl6Gx54/v9FAT7iM4AMHIATT5zGM9Sz0oyGhReHpwAoLfAgIgOApgVMXN6nTJvUl
5bKbMfSEWG7HfElMT7YztZjT3cv3eC2R7/BkJit009SUAk/7VDMySojV19GSKXRWV718qMDBWT/N
V0q+iO76GT5U+3Y2z3P2fBfnO1PRmgeZO/piPWIEHjC8Ub3LabVu5XWzCKSnRpSJYjTHqFnq3n3T
P32zGZH+vT2yoO+zXqZBS4sXLw1dOuoOYmvMPfAlWJ8WOUJUrJ5EeeJHFRxxo9+MhvP77i4fLFPF
F4edXmDeWO8bguM+HYKKbdrMRGknhgPIGyoCbRW9KYOj1XcM0sJRYlOCwV02I5GUyhzjBoC2M8xT
Higt3h7zpnr0NWuYLYzQbrNMTN8Qgjeugg9GvzVjmuHgLsIHIlGXZjN4YkVhoKxOgPWLF2Y2xbtc
SvbcXvEP4hITL5hFksOy2xz6kPDBcFmDDRU0ksERSLav1HwSbh8mFmhSi++/oiCFuI6fUfFskux2
+tFhkTjrXe5eswpv8PyC8my8WXMFfPr2DQhj80rI9VmXoQBI6+GT5XAj8ulu1kmNn0ow4sH2VzbW
nkQ+dTQU/BJTXD9H2Wnb6tPMlTiA/x5dyeDYEFWfARSsVO+xAO/LpYpJcNjhkKIICmUvhLEzTvu0
2hsbujg9l+OswbpQrvu7AwKvN3yrCbr1N0STnh9cu2pf0BpWz/NbMnKbaEuuzV6vOT2nUgi69pdk
9lp6Yruxs5pSxLyVkxsra4sG99V6FqiiIcHwEpJJAH8HnN8Kt++arRecPXhUVttAP8puB0ZOz2dR
/uOUAFpryNLaxr5gLr0w46aTfJ19JlVtTZVGRu11icAiY1iWGbTCEmTU2duSzy2F005mTZecnFDo
MzsowFuf+ccs0roc4dhJt6kzOXnk1cj9xFLrKcGg+Y7NcHhwEPVpJHGEkFpJe2SW1dYNClEgdzcO
krSaTQ82HK4iEgUjwB+C0tAfUDR+BWc/wMAiYYJ4FuRflJffqrZAnTqA7ILNA474Rs/zJDEBN+TW
P3YaDkCrg3vujvIK4XnBxNsVYptxbqoEVWV/thLz2k/u//P5w6/QqgKcc+/pTeRj9OGTE5/eAVBA
AmYfVskgqDj3mKUTybFocQ3MolbeeomQsXdkMNfjAIJ52/JEvOPXp0U2QwfiFFVgN/b7GfNWqM/f
k3dakYxDPuMthkZQPS6leL7VoPandwUmm0ZrPWa9n5fW2ewxxq6wF/cht8hVMe+PvsocGEipelE5
lZlJnAus7R+ULKZPnCi29xXV5tjPCV6+ZUUiVC1MDk9spE86EkVOu8dUXTcxpErRdP0rPiGGB8eO
c1LE4CuRYQj879JzTA3I49UPHmkXGR0aM8p0wmo9D8wDZbhIVizh6F+umDh6F2N+i7JBeCOnwNaq
jry6lOqGI1ihtYPh01SmUrDj+JB3U/qwxp7Aj5OwRcSNw1oM4wFyYwVie09x07sqzYQ+qBmdpcX1
yPeic1LElxxqbT6GHhXeMkAeJItv859wjifuwEh0vJ7UUkAHPvzyt4CFpuGMQEXbTTfP37+O80HP
4LxBoAYBBJIBltpV1aWag/nxa+n1+ssOp+LTTGsV8VN7xkVNnfQx7tpmQzScaXHTw+XPXA2851X6
yPdroM+jWHAWyu7noQMmQqWDiK64uXvKDPj5nboCwRum3VsLEWKfi7IZUcK75J4aYfIdozXvPfsF
ag9wVFFZTVZefEFulXBmus1nLWa5dOGLpxfXzYhi+GrKHTeIjAldkU2PYEPQFQJIbrxNRarVD8YD
ZFkRodYoJ6DWBfQroa3pBBXTD80n8twXcp5/M6RuI96T0o1VI+X8Ic2Z7Iajdt2QBvhj/K/ZzyVZ
C0RyBSkpOFPxoA8cv4rjOOn4a6SbOYPpe3BSgUPnl6IoZd0jCntBROU6kneXqbgUtSPmTn7Mvsp5
pXuA68pjRxSQ4VquaXv6LWv1xbr0MOcG+fUYAz2/HRsDlwCq49ec2KMjMR5MxV6JpGcYnQcM71QV
1cg7x8UYf4g0bFLcGx0KZo32rwMRH8wLgGVsDIGIZ+Ch4D4KNhOp4rHcbNOhQIw2PN+p/qM6Mk1f
tk/01c2mB5sv6EinibJrlQqdIpLMCoDRRI0S5sDftmoKRqG1e1+JX3cEVo1xC+Ahg2QU9GZwf81I
Xebgfz72EeVnmV+lPM3lvB6jz8MvmFLjdUGc9xqpJMCt3SETKD3PEEaiyLK3yD5UEEXdydKkIQxl
mNxf3OMTiOBfwPhyJ7VwXrqCGEHIh7yMtdFK1JxceC5Q4jrivXYChi5KIqLsC53Yu4kVtfvvJUf0
NeWF2cR9c3cSLo+Vrbtem/Tykbu48tMjCI+C550Ao9nf//v8lqXMN/cfndxrO+2j9V/h+YfHvs26
hxG+JYWS7d2RvGqkpuL3hBzd5hCrvzVbDdTmP9SDvU1ghGU3856dXuRtWRsxArXRenF9KWcdgHQp
tHCmlgiF1tyvuoBjsEjyCzHb7a6QPWbaGydBB04PH+yTk94KcMNT9FMiXwxrXmAf+2wOdgM631sl
mVSL39agaPd8QFeP6JblaVwZjTs6wQQEOuBkj+3B9ymXmRU1laqVNwekyheJy9uSrti3dSfpq6U3
le3z4MIuF0O28d/7y4BOQjiAxTjkmPrOVwv6npllezFuglQobhlT8jwIs0GncOROj7t+se7WKZAt
onTPMwpS7fFaCXkC1NcHfK7JSWUTyUpLh9YsZxRXoRgHKEvr4OwLIOWOqPf2JIlR5uo5x5nB3rqS
aUg2XH2CCcPobQVeHbklPUOne18oXqszjUdK2FdSAEhkc+Dn7hgw5T9ppuunOvKEw+N/c5sMjxX9
9LT3yGcjpXHmPpHAjqgmE74/ndFJlsTO6xQHJ3REn/svauApWaRGbkS9jEWK3PZhLQ9SlKQcjyb4
2Y76C90J60dYRT2aRrP8pd19H2VtwExgNDEqO80Ee7sBftC9br25JvU/bQZh8gtxzYnrHXmpwjlF
360zYpr22VQX71iYXxzvaaYwEI0zEtYWeyaoPVksmN7HdhEBy/Eti8O4g0lzIIiIXSrqmTW+JY9n
LZdt/LnGcF8rbfYoZT6M+CG0ZMRH3DvWCfZWPZPoNSUDme0nkDGEBdZBSPpoBvDtCLwjzVbPbz67
Y9oka2wDBKdQzyygW/LWm8o4hAaWCX/1725qARKP4LTz8m1N0vRIDI9GXA8gbkWwaYgbfgtHi1Rx
TguUcJZI4AJ2fO/9kdIJYcDTyNHGGhcZM7lkh156CPK8mq4LbBkknE6Qyp/qpJEN4EjCsfENZtFw
YtEKYL3iGy/ut+0pdRjfUQkWQp9GiXDOQCyj4qyS+2vo5Fy+Qs6wSEjvPzmKl+arXXNgd605uatx
mLgHZrDVdOd4BVngmttltm+MStFIX+Nir0B6vzEVOELuBYXPGHttZ2+ayW7UIKrOdOCjgN2sQsGJ
UnQ/eplTbNFyhUJmbj27uhyPqYpkOQq91+mbH5APJvPCuf4Od9dfWbyYEt5DS06cBPrxlUEN0fzU
pIIF3y1tsVK+i6k2tkc6eh5b08vv/N5Z0LaK49Rx3J9AgENga97YYQGKHS8YMr+Zmy/E7LGvchVh
ymVTaPyNjV6noXijzb7q67LYkw2wyEja2XclcQNV2wnGTTrqd+KTr49aY+VspRIwOqHLJT6MQ+5U
l+18Pr++Fw9akOX1NM3cMDcxlsYc4Aaewe6KdsFc4IU4LTuC7uGS3B2hMwdSLTc6yJhSKOgXpLyE
xfnE/k8ilD7KRl0hwgu1rePli3uY6pQKFheLGK9az2OfPE0s+617s7PIJhTThT3xRe31XJPNMDTq
dslwmoj+hponB1kE/VuKNTdepUTigfg6KdR70pnmCRDqOyS4OriR5Hdz34IrPmZDypMuYOB8H8EE
r1Fp+kJFbTydSWlCKuHpNld9XEvN3vTNgWKZR+QSBG9x32REwI4GK5+RegSPCKI9sLheao8Yf30h
TPn47Yy9bJ8V0F8gQpIDBMRPQIoFiwtWmr/K2UGgIuiYuFGUUkp8gBnyittq4G14Gicl8a03tDj4
48EFLxtcHCCDvDzbkr5NPElpX+QC0Fs35MrlKfgDNGCAHPWwnis4vWLstuS6MiPvspmaAdrBicj1
E7hnwjZucF4hlB8mKnORgVG3Ch+lSJIIDTc6osD01ZGp/NR10zDuc4EjN/fAscc9k00jQp4wjLpq
oS7nGSeqEk+LKZuBnoaklmhRGmdwYOJgU3OBLGmH/cHzNLgi9Ad8zi9KlH+rpJQ6xN9pNPZTJPeZ
zze2IiTj8afDrA2nwNAPbqdY+y6mtqk4oiYAhPBDHI0RA/lFnWfW8REVfyJ4wcata8Q4xYBGKfjd
EyQkS/QsK4HIkNQDhydo1YQ1UNkm/PlwRmax6TmzIjGKfOIafA0KxC1jtZ+Dhy8IaycRwSkqh+rZ
/jtOxvjPPDMkC3R09bIiZsNVRwcI/jxRJiRR1m2PApkwDDpHtWur8eZf6JcCJeqn/TgiiIGH01YO
ToYMpqvT0NIQPAujuZe8hz4Wnvj0iMedCV4xC8lqs+wRr/EGAYDiNkomuR2zEOdQ40ch39nvNs+L
un/bO/bftkrJWXXIq1J/3tHBP5ERat0JmnPwP8xNLzpL0wofykhU4+kok9qj5zd8EamGKRlEpRtH
/BDyZbKdUWQ3RsrgyX2J70fL6AVSibAuHre020BHngF3FaoP96epNcEu3QhDDyWyhCjApjQNoZUw
MAk4gavVYfHoe9TEQ/aoLCZ+cAQon6KQvNJrZP0q6eJTTV8bWPOFgJG5IjBuLRYw4O0W+XyUZQAS
sTlGJ9ojcb+cw+iJj17uEKSvM222Q/l8BW9oZm6Eam2a4s8ZzPHqMyl8Nk7J7khQQa5mfjezhsld
V7m6HYfwT721JSTtKaM4Tf59k/GSNqHYPss2oIxLjm4OTUIq8/U2sry94tyxW53ghZdI83k+5aiI
n6XNPrlq+QY3GVNQvUC+9UaAv7VoLKAzW7ShdKAK/XSwY6ODZtYJqfb2SXcJM/l+LxEocDZ6wjwX
1P3GA7EnDk4mPB9KhhOiOUZkbJVMCZ8jJuKYq0GrkPWV043zafDoeFvUjPVWHm9Rqq9K6sTps0yB
KTcGD0hXv/BsvDGuDX8GhwzVQKDry3QQQsUQFiN5EC3VALhdu89DJVOi2lnpKmPtF7cD1ebgTUCV
0WeTLcTNYeKGZLNT0k9T9b3iMN5YGcMsM01t0HaQFOcodC8sUCug/cGbdkDYUa/ZgXVCA1NuG3b4
uJll7f/BP6z3LgfnpsE6r+JxRanbDoyqVvs5SPXQVVBDzcLcJKSXH04JZf8x4FzTBy4NyJwD/jNC
GS8Zsg5lj9+z+z+tTA53QuLru6AuSABI1250ezkUxccZ+i6XWHGOhwkCaMD1hUtI0Xf1PnQ37rTV
0OwpHOGUatkhFPCvepVfIb16F01aZ22qgwkGDPFVg7k6J/SZr54zV0ILkLLgJNR3H81iZk47Ubhe
EaHJT2SjBXKN2qtouj+6sSKgyOIoA+EOGM23jrbuyA019mlWo4vKQdhiJLeHXWfenaCshdGJBC6l
AJgkshfr1RWJ8fpHpH+KWoSjWQ+9dfoBSK0mdklHVLUV23jYWtRauq+g16YdO7uoSXBNQerKtuFV
RAWHpzx7VE48WCPXGz5tXUjKRuUohC2lBkOj3i1vaTeES8y2a29VFjqKNnoEqinv8apgTCLBT+kw
hwGSOBBqj3l358ty6P8x7AmBIOuglX+l5pnsNgPSyZUUG3v+RYUQJ/6JKrmgzU2YMiqWSCamUXDx
RKlsnjuaUNoeIB4J8WnxBBPZkWsQQh5adl9MET3T0BGVqXt1adw6v7zvflFilJ1qMEh4Y9kvw8Zl
+0S5jlcpQUl10XNr5Uyvx1hEGnmZh4BIao04Z5KdQ1hjjvi3izGio1b/Up+GjdufBS4AHiXzgHiW
5K91jstpEr+R+wfxlPvH9Bnymg+3tqVx0b5TNPs2f22vNpRJvVDPb+uXC/dtLQPLzap07affHtb2
UJbMqvbUZ6fKJ2f69jmC7G/nVGF/EHnQFLJkA4WVdeRXyuFNih7q0bYvTm/XfWHe3UPD9ZBGdVjG
gPk+0Ws1pK4KYO7OZV9g+dDV7PkjY8nptrK1WM9uGTjj/N2JbP3p/jNnMzz0dfyevG98XFH7Uxby
O4k4DrriMzad19VVWO0J1L8jZP1lADitbTxEKTXo08jitYJJgFs2/vxwAGVdH4BD1tnHlCoS8S1f
hM0cj7TD7xoXqeRA6IglSrNaLm2JHgXSGt51Dn/h8qK2YY6QX7R4jyasxMJWGmaK08LHj+gXUxR0
JT5ZsE9DpgKA0OlaSnV0sPCGtB1z+zN7K/nw6BUFjjF89ZEjMK/g6MBb3hVUJCAP7JKtrO6GP0x9
bPfJ3Jp3kH7AmHhNDHA0TTcrBKUQuGtJTbxLCgeyU0dByt6dF/8YhgJa7HPiwiUk8kDGxcni2R+U
rIy8YUGqFADjAJNFHlYnyT8h4Y/r5+4NnVj171Vt351TwoO5503IBW6JR8rxz0Lbc2sEqCMU0loX
tomVphPTywOIViloS+I40DaLE5sDwB3OXs4mWO6mDyTNLg1/UCYcaba5g7RHaKobrzF5FVTYPVe1
aCYjkVgY3GqIT0WrFByoObRHgrLNAaYHBT76Du9CX1RNRyU9FmP9bJU87vWHeeANxU0KrIOYRTjs
Ee8eG5+eEdVIOHvAl6GtoqUigIfyfJ6aINzNbDiG3OnHQCWmO+VPRcSmJl/osnskbUeVZBBpJHGa
H1sY5QAw7R+pNfsOAWduCZmTw68NY+fyNj8dcJq3ST2A6K9KA18B5C/z+c9IwY55/Ws+lsceT/NK
l+5xnu0pMEieBSS9E2bUKAf/wHbz+LBovnoKRSHZ/ObTHtkVbfGvFpJxGvGuw1ohj1HrE4sKw7MD
4EOOI02Ft5Wy40wEd2OGccbq6HmoqH0JDHWpYflVCa7ZjxvXarZNqk85DOufa4Lwm+pozsWbwTM/
AO0Z59luLP3qodE/Xm0J5/BzxebKLEBypY6PVQZvTfP/EMhIAyE8lCOIqh5t+gJNO6/M16s07BXU
aNjA/KaJhePeeEgPM6ly32g5DtnHiUVFpwNst7uG5hxl4jqTwfFrRTfy+WeiAoERkEtmjTjq2GCh
sX+aZJFnarC3URJ44vnpAzSOAQYd8QvNYgMMqrUoiUIIyC5WcSu/Waic0Ie5Z6bMrYhUaE/4Vv+O
/Dkiix16ryxpv3hdVwzTlaKEnT8Zq9zXrVKLtPgvnIhwwLa7UaTRLaaALlnTXMflQoMxV6Vu+FrB
UxAJpdbA/a/6DPjzJNG0oTHWIIQCNPQG1YUBByd8E1O5exECf2z5bh5k1lDRrSvP3pF03sFt6FfV
y4SpTJVMr4+yal2UEDkPpPeCtlJXJrPHRPA8IORPxHmVMNF6NCy8oYM8lWMXiOY4Fbn2fq2wMsjq
iv+VnrfaM31ZQnjb4THiQVwmp8OXiy1SyMh6c4T2kbozeurjB+h2DrPPZaC9JAuoXbwJINKicnaX
vauLg+i2d+ycoBZnLTE1KKprWO6akaIjDvPtG50gUMfWRx39yXCPHZPNqsngpLAJVqNlPrLC1ah2
StO77UAuTm5Vi6PlD4UeaOxXAJZhEoOHdLjizHShzX3ObPhC09KhFZhZ1rfpkMOFD86HBzHRIN5A
ZdKYEZvI4bf+I/FUIu5PWQtqlkp1bGv2/ui/I7RJekwVzBSp7XbprFSmMbeTm3FZIORlg2J72tyy
6y5na+R4LC9ApD5fEFXW+ReShqrJuIgteYBx0ARMxJCjApZh6uDjMi7j7gsAY6jJO6qYGkWfQP/z
cJjoqwulZdrSVTn/Y480Xe1P1PnCoWOk5fjfZu4ZkjC+72lgnTkIM/Co1Ow1NMUle5oyD7cJQUcV
P1yqZEFhUwblvcCcHSzdbUnyWPtRR0mt6IKhU7Ncx6jgu+DmV5d/6lvWC1tAFD9uIf5xqGVpGidn
Qu2wYlR+2UwDhDhVHGiVpq5sPzcbiWrx1Hcp924TXqeiCFG8FJX3Lj06PO1jWvsgaRDbuQJ84Q8g
3SJZAUOahft3+GMnadiI1dRwIuVR2X+Q2E/b/4sRQsycJLPTbSrlxwaEt8rooyFNiWZYPcqVbdRL
aNPYP+ZI2bARX7GYr4Z0HdTt54Ay7uQVDtzW4ALbXTFzu7SRcPBJbyZrndj7YV1LZPC+nBwcT6E2
4PulAn3lchDjf0Z9iT/BAidTfV3CZor6jz8s0n8ExEy+hprg++wqw96tZsCf7NZo98P7eEl+kI18
FlRQLfdp+jV8sHfUm0IdXO+jsgGR3vxQXKrBJPGWzWD7e/eAgVgFoeM1zdXx/aVgs2bL8DTw43or
AhdhbUESlHe6vavlsw4Kfqdct9SOVFXbd1M93upG71JX9l4ABRTZOcI8s38wIi4FPLkpexeppE6A
5JmcxeLX7lZpgBULGLxiRFWqfeJqxRCHifHG3xUA9QXLTDeyrRdoJQsWaJvi0+B4Aoc8XM4cQvky
+n5cZLB3fT7Aop2FmmhLF5Q34X8n6cFOIaQbn2Pwit5TTTTGon6S357AQqPYZSqyjOGGHwSWGwJ8
kwIl2JIY+Y4UHxqjbQ+o6LkqWg9ahYzqdqoEKYZCEoZRVuFDSCpjYiRMHjpbnw9edRD11LjJ1MPn
WX6N27xea/T+PtjXivoKFjLA+Bs5feM8p4uKMkPNJXM+SC/SZnT7REkq1Lr4bQeilBTApLlXkRka
YxpMwopAcRhr7BYeCtAK1mr4W0oJRMnlXUlEPAH1ouX5oaoqHGvDF79Q6Bn59x/x2wClDRZAQORz
2DOyDiaA6ku9kW13rCrDmS9dtTkbfoLzYsKCJyIFlDheh/tJYPo54p5WudXeAqOc8WV0poONjPg3
uTQGFBAsj68si58Z9shFnKpZTMTpAObIgs/Wb8dovb1DONRZMImZLtrjywEsnXEyQKEi+lMwVaXr
/cDRYHM7CR24IzBm+j+GaYhROzHKoJZxQebhB5gsl/ZJU4DIrZcLR7YB2mzx+5fkiIo3uS2VHBHO
UZ19p6O0hN/6y9wmgmwhh1grRygPM0ZZkfBvlEnH2VRyCePS9Ohkr6Ulhh4fEVTW2dozzNMRIe7p
PgMn/36aTrcUEgTElkg8+OsCwBbnjRR8xhdSzzouXJ5SefYRDdHs7ULpWb5SmLyhGiZv7VzUyluE
YsGJ/MzB+wmNjnLrEX3YaT6N+ahsiM2jAtcxTda9jg81Pg0gX+zOezjKS2My118ATOn4xzcpTK4Z
jsultvRdvwxTIVTZXSl/ZPnp9+icSzkikzahIqAu7AjvdmcQk8g9EGuowFisJnATWDRUzpuavEAp
tNE20z8KVYMawRNtMifcaZFoUAUgpVCQv1esiApzbKS1yA1IcdDQz+RxK36R8VFGbtKqtJUMbeeR
fxPd2lPX7PfAE/CcrpAzua/em1qPF9EGdP946h4A2F+zuamT8NUm/6HAarvv/9DKCf/66UKg5sa0
K0t+l7VKZG4/V0PDR1lNhh9VOEF4Q1yiJ2dJ3V2L+IdiW9jRTz0VLZ5U5DWecWeZ5RIN3V5GlyjA
BWVYB82YBU+WbD0zQLy32iifWfR8pzZnNrhJaGwTp/1OAL5FU348vwnFTiWII0WbX5o5I3XsNUKu
tVeTRmXwxwsjZoN/1/mFWVfc38mDAQ2+PJW/XZrOjamNPO1HKS9WcpDiZlWLGX0ma75E/J1jQ6NX
uTeWmif02jYJuUjlCF4qvMA7+Wel7/95JuiR9/rXmwI38/5sD7f/M4jQCFJE/UDqKx+4iOcb1mfe
6Mc70Lg6sU250Qsd0221ZDSjrxZqmHI65/hKtZybpS23brO1AezX87cIuTjQ+FVH8vdYeC0EHakw
N00igzS5XHbJ5wwmHjJVuzhTpexx5odjWfxwqJ+hUB2POs4Gmyj71AT4aQhxWBCCGDoohb0GpytV
OvJvJ8XDzppx7ews442l5mYsRUqYw1uj0zIK3rzuigHHSGe1u93spF9zjhve7nAVraB9qn5A+O9p
nhg09z1InLpbeFLuGqOv4AhSgUVJ6kok72IzMyiwYLJJxGeGAsqjG/PVpigb8ABJ19mDK1U/E1ho
kqJUh0l0z6neiafxqDq6ewihmlahhyehap3I+T8XAMo4kKmdhQnRQaqIIT0D9gGVUsf0WtacQv6S
dB2s4JSEDAIPm9wxoDIhUxdG9A3yIcmZBcw7+gTv/0ltmt5PqNcbD9URB06XmgcrdDXCcecFiKF6
y7gQH133keUCe1ABtSmOXAyu13K7Qyzkf0FjXZqYwAn1+Cprqd6z5+5q9756BbVgxUw8R51zWsTl
/58GmDxJ+/omqMgVruQ/yXThh8q2AydaNFrbLIHbkmqswgDTw1U8GBMZfl0x8JHFGo6HTLiHL9zw
bcomsf/6l0cwRHhL1oZhXiySz4H8hD+2WnGqFwEadH0XdSQA+z+BlNPB522uCvqg0mgKcgMSMHGS
iNSTqqnnec6yoN/b1GH8zUXHI0V2paglMdC9w90iAIxKE9eEKazHpL1mcdMmAlA0BpqltahSx1ge
UpJyTHcrN8hdBcyIwH+wY0wHxarqLBw1Dxkb67Gd7t5k5/fLjnc8kOZVrchnen3b4mdbQKEFmlwy
kEBUDqq1ETLYz8D5pqqK7HBFiFbWbCuV3ffLBJ2GmJpTwvxlM9k423iVJWKUovSN/1jq/rk99gla
++8kji25Np0tcp6CZC5Q3MUSb8Yq/WjFUKVOZ6p/R0GlfzdehAnujKPcfIW5cZopH9ylDtQK5GUZ
2xfEFRSwxfxnnXhUZL6y3f42QmHyAbJLJ7hPJzaHWP3XYBYreiAV2P0w1Yqi5EaRAp1ETr2JmeV3
sDkD/6XcrcMph0ZtCsGRdy2vIrOThUeu0EdSeMBM5RXXqcscOIF9+p3VmhyjL4dipfXbr5ZM/9Fx
fUM+38gHWmbN7Q3e3yM2L7oAN7guwWl24s7yYZE1fGQWDgvWk8dYl2abRJMwdNHsP5vcyo49QfBu
Vxqgo+v2eQHujgKYnhbswkohErorPzbYLqBqTymCBiQ9j47GC/zi46A4y8baZsfjlnnTvTRgRMTr
uOcYWNSM6Zx/s3AxzbwoSJQtKm4pRgAI7OS3KRx6lkHJkdLeV3l/mxgMypanQclmFJ59IEFUQkI/
520fyAToE+iZFCDxJNgYpvSgpG5E+7+V0RTLMpG4AdbXyWaoTnrjmtbRqgxDvG1EisbwU5z9dt5O
5GviZLgNKfaatGWyVIuPMGDwpG9ul2VCPC6tDZGJRhP2NAZ9z9m/9qclWo7W/U1Lbz20SaUIOSaz
qrSoSy/Sn6+AUkUnBROwDOUA88htcHqrAqeomoj1RvkjBdzqm9RZp7h1YW/eqy3I+Jc3+ywFWisN
XusfXpTu6hqaHVPr2A27HAV+gZMmpI4hpoYA1xCL+D1qkWlW1v9U5d24Y9/s43hXTiiGX5NRfbBt
i+YiVJt5ffWUobgvQ+z4jbxypF4YYi1HgijnD6IC2GYpv2LMkyy0lNOg1iSkVbAhaWcuck2vqpLf
c+8eZWSywnrP+FFWIB9Bu+i+MQuQBs68+lrUHa2fLEZEmStH/wYSvh7GKlaLVgXrpoyhOdrEyhIX
6SHekh1gNfVjlhlYCn0Qg0obIeU7Z0wA5uE4fNua0EJAOsuUj+WEkoUAWHRl/Jm80elTL7c5jNZC
a7QuLSEKdn9QEl2v7tbDh6xDj5lHNgoYlHBHwS60HKgypPl5qZH2D0Uu3JVcUC8Z8o1QTHWJp9NY
nao3vuFaJeOfYMjGwOmUh/MpdlJ4h/XXogVimMEfCKkz15jlumZGHWqQ0SvMBciQ2HucvSA4Njx2
IxVoTKeTWN9wwSs+nnq4OElhzbFgXTDZdTYGkpbLhV2rgaCThmyCGG7w0D0RTm92FcYhgnym2AsZ
G6MHr14HwKsC27ciwcncgqRut/PbnfXxPfxlevWOczn/kcZuY7kbcL0g+355xclZmZyQ6B8/7Thf
eUrz+e6qHblh4MHzQrwApiSk+ic1yhAhW2gu2tpCiBGbGDheyEpbrMsMJ9WYv5darM4jMZH3cEaL
N3B20Do3M63tjQQi9IJ2C3gN119rb5BabIQ88P80Jy9nr119uaze+te0yEAm/MGznT4vBRKOCfdw
Rli5HD8jKfVvmHLIQxT9nOXK+hncSUiHcnKrNoSONrgWpkn//t/av98shwK6O+enxvh91owMDlwD
g33JKGmgwgIWJzkVdQjeGxCUGwPvwwfbr4W3a5I+cp/A7guFOrD7D1+zChS3kvck4a5wPBd36OC9
qSp+y5GgvdmxS9yggjOV633ScLIyoV6Z5U9ibODDu6m1WlryIJoyoPf3uoA/kgWu9fXuxxqiNpMH
BKalUneB53Un11ykKGYPE0znwCeMdZz2m4Xz6SFmrvEWOCrNK+u8gKcsvLOHtznvk7+Uwoid1SSq
SCotjXXGpth61pHlN/L9ATwSaqyIYIltbpzNSlVQC5Lq2KFS0uaqNCPIbKOAgO0Hae/IqcOKyvhc
om7PbtQiqXc4I90EA9SO14QioepxU/UBdrLUeB6pvXn9b0b8O0b/IXxFy1mKeoNjvD47qBMlV921
doO2RhH2LR3PE4l2sQ0UMqRP/BK7/BBa5rAhjtyU9I+t7a+T5e6cR9jB8u1RvfvK26/DDHIHVk7v
SIYTpWPRJxnr2JUg2vdqiGF2fvtpKWG3Ko+Uux3c1PJ0+ikgwVNy7SwOZ47kuKcWu0otqP17pyLL
6b0Qnd6vAQKaTErXRTLKU/RXIjBAktVxGF8niKueloDg0uDex7Lqeud//NVi382x6ywSgIdWtANd
NC0sxKSn5QqWJ4VV2IKz9QY/euvUDMcIq7ow4pg3BzJC/DX+hWj7SIX07pFxcDcVi1ELc26F7v+Z
wTrrHvatvFn9EOcDNSh7qZTQ48nkXRbHX+ORAxkJxIczMfgdU8bHEvWtqOVxaVZwdFtKClHDgnve
h0VtrY8bMwz4fnM97vMkp7hKwclRl3YWFf+ovJciny8FbZT6osZQSRL+qbDSVa2UqAgCI4jQgH2p
cSUhyMaWBcC/Wd/ymmO7tXTW3yEphUs78Wp0Mz3UXqAU72dnjfajdzTcQxD1DTuQ8XZjnTVD6UQy
bl5t4FIHrHkLPBMJCyq+FhjCcyh4j6TO/wlEHVGITa8LvZcoMK540++psPQMhY2wn9aIkmJ4KCFH
08PX3Aez+E1Hj+be8ihi/AZ7DlCaRMPf73Z1AHmYE2HN2CZwKfuibWDiAAnMxD0oGcZqbQN/YRbR
sZYMRYYIEdhVVabrXNjr86D4UXbcZcSuUVnNkgimN5EwTZBK1hVx6/cbgKyqFUVAvWemPk0Ma+LT
tJGOoeLgYnaEVw5z+CJ53uPJoBBkY+8LQfiHmBs+iM5XXwXG8BPatxILZqHt23yetRAXRrvP/xnj
bnKifyn035tqmFPjFgxJkSCgeGC2p/CwMr6KtHilmNJ6vT0o0uIo2oCZ39IEP8x+OWbrjst9l2x9
qKlSeDcxp1gnKaUTURsQ7MUfHxwgAqrPKtg5SY3+8Afu4CFwPc+C92oJQCNfSKYrOWajrQWY6aD4
MeyfZO4tnEyydBgqRDCAENsC+gZ+Zp6O6ZA8kVphobrmqX0isJs8Emw/Q3wsmFxM3QpCYFLmrHLX
P14SOmLbEGoHnpSM/Y4gj8gcA1qvs2Av+35UtEMrryrqKZYuwj7H2yLTIbXR4zS+thxLQH0uQskY
ZUl6LJssMVvca4ukI4SfMW2AJkng0dYkPc2Ev72+dhc9df3X0cdQKs1aCxFGZSa6kDYk3sqWXavu
DUo5ZT9v1p0WuGM/VnGPhJjVZqIaT4jKXVbFakYxU0AMMX7NUk1/hV0DOb0P2V/0CbflQHXENdkP
JkJ2NFL7u1wec45Zj5D+o7/gPjMYmS5F7zhcSWeItk82Z09Htg/5m7N3GcYeuhgAo8gBCJEvWkpn
ULv/lbw5cgX3qlZ4T1Z5vvfvWNAkhX8q+0LQn2domP/D+CfpT0SMD0tpWd2qCOznA7Di0P3D4SQT
0/UdvgZPmnDWhLu8Ne7prto176/fz8KxcyKVQqqvOr4E3cvQEOJ0DXt6RQBUDl3zUAXjryBDkEEz
PTDYLIQQiC7FZo2wO3tHGdd1SzrsIr2CvgjzGBA78WZ98kwsYbpMFcrl2psg0/zT3yciL4QKOY0d
lNcRqyQgB2WB3squYk5nfCDWXrB5fxJvD90EPnG3w1weL/KMwMV4Xe+1w/na11gluouZB+8nKQDf
Y+WJD89rXhXrZITHIthAMuwO2H1rxqwCK4wuUtbcU3ZG/Y9eAbg5fofbx2bEauosW1RiuuY27U5m
RtklKD2qaTGyklrBCxnrF42kQNR8hwB2e3bpQouOj4yi0HQIHy5a+FshRXWtx7k9RJ2/OXorvSf0
lv2pmGYt2AT49iJYCjLXzFeqMRzJR0QbccyMI5rQgucMaHlfA3l8Cx12Zqwm4c0zz+ErzzmrjICe
At1DMeMKQJj70k9GSGF8aRyuiT7N+jEvn5nbsFyxibV8gh9pwCE0n2onONFQSTX53oAGayXw+Az3
G++qfHjfv2W6UtAhEZQ9ZJgFTfuzCc/7mQYLbyGo7WX1RYyxD2tATDTIT7amEZOmUbRMDMT7bLyf
wp3iZJ8Jr5uc/dx4DP2zoufQIWTfp6gQvQl/nYonjeUBtX9xv4nKrah67XE65/120r/3nz+YFRtX
VNF6Jldmhirvn6ZonUI4qtiBnWNdIQemN+C2GR7uBIdFHeFbh9+3dXTmeZAL3zdtBipq9clad0S9
AzRBHP8eSDzXfmBuaho8COxsM9J33o4j8XVmOtzjPoifck/hRNV/ZJI/EyesvXxJ3OVQSIGaXMXH
LZUpiKN6nuNV6JYOBbCMChQs80AhgnWJ+h9tzCsrw6cEoS0WUrtnOXIN9wOH3PKDCaJJBaAwB0Ij
Vjxy4DnCi5tUf/PMpREDWxwkouS6IeiGiLjTmI81owFb8vFLbIlcSMJtViNF1BmhcQMei4kopiSf
cNjv3X3JNAJbeyspjDRq7Fjlb9rW3B/objZvDSQAdVru2ITemWeS6AGux7g5ejxFKLF5Jt4xOGyG
CiLDA7K+V50VG7csHnEcMfC0ddCFn3nClARXDFPmmCmIx9GwZA/rLg7DtCm0y8AeuEh88NDY2IBp
yXydoPgxBUKsZKWBzVzx+oxk3fSdqcjuddR7iEyhl1BTrvqd6Dspe1wMuSGGjSpfyNQ/dWsb44F4
bN8OBwMD4NM/g1MuKL8UQp8ehj0PGzT0W/LQgDtIiqeG6EpQTfN04AIHtHMy7OaaQ/T58XsCt27O
7fcWbcIUjgqX39Pn+pcVXVlFaky5KYNXVtU27W085OLnnSFIZykCklZbEiaqIrRX5QTWr1WzkzTC
KG7JN00t/bjAjdYY0PmGE7Ncik1HIAfAtIs3IV1XaUN3nPHzf+tgF4sjNQM56OnzzDcKPaYmREdI
7l1FFooc5Vshx4YmFEkDHoDnhNpPXUrx//W0ta7KzUTr+WFk1je9R7h9oiOkErojn5oqm9ksDLcO
h16ezbgCF258AIs1ePa0P8fTnlppV3bIya0WGRa1tnc6InaOqVuCPwpX2nLrYG+AIemvMSWYHMyn
HHvuzS5e6XwHbXzKNMmcfjw8jNGh0kHqenIByJLr8ZbcwdXRUJ0mDn9RBRa0jq3VZkPpTVPVAlas
B3g/sStBOxiTBb6iNkO5JuSMMyQWyq/plKPlglnZ3RmcTUEOyVbXE2AI5tDSmH6skWWCQkPKFikG
pIVAQHWeK2CYNkTeMQhdvhcfYzttW7BrBM5Y7oEYEF6o7mbT9IabS7RBH+0+oN7jfxObbBC+ZFYh
CVVslgLvlgL4J9l7/Svf6VxJEAz0qm/grz783yl6T3lcj89yH0WRbWbZkjMUX/wUnQgde4WwLdJI
LCrLs0ufbM61j1yxoxOqMOyFemY5csVwLG2W3K+DwIdR1Xh4uFfXRBQAqOZdgKcWPzuTjzqsfRb5
KDwfEnSfvttUHs5VTmZtuAmlCB1N+Krf6ZF0gx4Aa+3ugZQnlC1A/6warQ5ZhPqC81A6n8/GqDy3
9M0KZ9OqnklWX0kN+efXdSI9sDNXbRIdumd9Gs56QY7V1KcX9/fvFZVufSuN46MCd56W2/4x29zy
Dsz24ApIts6aHbN+JSUZztSlBJqWL1oQyyKYfRPFDgspXeThgAgJ0JQ4VLCvhSaUeerT373dXBCk
KTSVmBbE3F88VlZPJSyTOjAx8IBK3hvXGwfOV47CAH5TyP7hGuxTn0fCPP9AdjjPcBOz+qu8oOrC
nD0iFVz/B0GHsqOyiVZ36mOq6hmOt+zHbjxaDSnV740os2k8ppq8EF09lwZHY92VoMlWE0wnt16P
r37DjCn7vPhxI5CNoCBBfTnUMVtJ10Qzx2rP8oAPi2+DMOyBWUb1uGOEE5/GjI3OIGnGDpbV6prG
JRnC0l0EedZqnscW/++FGngJGsO3n3DH8gNlTwmmg2HPChngpXf2LaSkru3Qk0H6HCiICtclfXID
cyXHWyTEdnGkVhdzG96O0G1FyPFgQLOTaawMFsZhdWTtE/Tvw5JddVt/FrgvGTb6FJN/qZhh4f6z
HWlxaZPJjyvsDxKt41e/+7DfGeVeEATO4GSesnAflhhWtlZwqw327t2Yf7JoT5wjHZ1SHaQPT7v6
e1UG5DAYV2Jc4wwPRQcfr7uryAD4Z39iCi5WoY2c9HyRC/CJ1dqqXu1d6vJILF4iLeUdau7qJCvD
bYY1zBghe//bYrgFG+Jfl/NN8aDwbA8wJeHugAczExaJe54/Jrvf9bfK+d8I5dfVcyPgM9OmX9Na
s6F0yFioW5v6setAYq6y4FB112TggjNZwj8mMP+D8pF4bKgWOvRtPLfGhzOVFGoytoqV/iR2IuSZ
sLJSYM6W3WyugLB+lDnuByNDUV9mcqBMmYef735TXpbZPvhtJjd5U5MEmTzYG/SQLzS95OHPeit/
Ofm+JTCB+LcL/Uz16qNVZ+YYc4SBkU9ly1X5dt2FdDGWcKa30gcrLwrt9V+VDUa/Xfx7UaUWdyL8
OcsVX4ZCzCoLcxxAgjRBerfrO9houqJBhXRj1YADdi/QGUlNzqlgyQdi4R8yDSNJmPJbRhvLWtII
V+VOz8VrMOArVI6rbYCIkrCaMNKmMbM2zcwJbYKNXKBKolVCz1mLkqnWgYtA4TRzxDTJXqnFvudj
atcN+zhFXJdBqigYe2MMy9APHOWKQwFEK+6nbzC7eklqXJSajRAIyqurCFBfHLIZ+ya5USMQRB5F
lmy+I08Gm1z8FTs2BgL6fO3XtKBtlqxG8SPFeUDSSWmgY8WTSrhMYhLs81YsfAjFPu9aS2XJnok/
LFPeovCB42xBvEcjhDB/tnC2Pkmfy5j4p+ZM1epHqXfNF+naAQSL/nlqAIbTP2oljb/zkseJBB/A
MIM5FW9wq6czvc48mt5XCt0+pKXLd/+fyo1IS/l3hWR1Klo9cpHH5jcSw7Up5ck5odHeHhBL+jqw
wmB4+trlp8ClfGk7Rb1ia8lsiYGs+LXvqB7350kxjHpIcvr2iI9aGQbuqEQxihH3n+Z42JUAUc3N
ZMP+FN6aAQi96MWlnMKeGzcVgYbMNNW92NjAU2B3cZYniClGvkaLPpqTNfhzY4UYUKX/QigQ29Ga
iYNQzQiDw1TFQxC1frDZDJSpe79NHTGoaroGi188M3VFzw/c6tkswDHgEah1I/99UUUI6ecCjwCB
mZMgOp9NvL8kRo1OdgL55bYN/9dN3Rf8QsQXkO0ymKJq8oRKbd5r4+9WjsaeRWItcj8IPOTU57sI
aa9T27Ay3EZJjbVB2+v/mw06eRjbmX4C5d5t6fEDVo70de2flJHbgfjkofGB6Ukend72NJ3F8Bmx
YHZcUWoGfoPhVbHDb6kGB0/8gQn4GZvOYJFbSzKqdA/8V7LmhO250Qi7LJIjmvblvtc40iA3Wl/4
lU5VqqFWAS/eFbEbjscavThS76VtFwWhzlyqEZYqxX60Z6whlQkotqpbtmsB+9BwDuLHuxZPGTGj
6GEf8YSghcl07QMCryCjMHRDYbIJ1+UNeyM2mNvggoZ9KCFOfGrRy8lOIUl7+IRmY1ALXVZvXJqR
zXq7SCwVtU2ewiQ3E5dN88DxVQ6GDbEaFkqGAt3fh4dPkfmrrNMWikkxj/nwl+AItbQMBE6tnGtO
W+m5kwBpRKBiLiL2tYnz4ltfqeNJpEnrBob/HJdeyFbPqTlxPIdVbzHWQ9c7nhmtjQ95v/+TFomT
F7XIiwjiV68RaXm136m1r6GZ7ajE8Cq/+PJOZAJE7uspcBkY8sPT1EoQKSAR+5v9nTogSm9tYY9/
7rVVtk4DN2VspHghLEFfGRTpGhP+uuL3M/zGzRs8ox3LtMxmNBjYerwxX9zBxY92TqwSehN7yiDy
qzvDjaU0m9WjWmEfD8aHvfjuq9vKrdvjWMnww0wbYMEcN8TuT4HOhqDkpZ5San1Q0TQWFty8nxjF
6acBNpJpfPBmM4PCd/9qdoAnYJF1rcaL3e59XiuXGzNQCYiwMnjIiX/G2WUUiJljKhxbNZG9VFRs
pGA5Z+ykoHSY0tCI5j9yC0bf/7JjSDfuPFf8aAuNZs+DCOGkSQR6k4/HVWWM4SuGgQvpgj8WjQUl
Kv5yBZP6Wcvjx71Br2NVKyVJBN/WQPj7UX+XluSQ7n0w+bLPhCLouFG4DawggHC7o3BDU9aaS2NA
OuHAXsXNgPToV3dESsCwE00+5dfj0v1lCYaHPSOW2lajW1Y+uYF7VGzzSg8QgiO2hPbfK1jYlhDH
m+MQEro0e8uF449H2YwQS7h96oGhkC4ha3VvQ+gCnjMbWu+FN9O5n+b5yNAnwe/9u8ybdoiEHNin
3JsX7XZu0SUoz69U/hFGbmGainBwzppB9CTYjVw3E4z9OFyXIBhep45b6prEINdF44O6hlygiJB5
nKHPkTtUIjJtZL1y/mUDbA1LKiGfwFpjMFEyxBOW2O9nqDMVefD+nOsFMvUsdCLyF4RFyoLkenwo
aZ7zcnXH78W+olf5+xlQYynZLVyxscmS+j+7HLP/ytkfFaLaxJX1xCDLnFGprRA0Kli8dfsvEaO6
HHXYovxwr81oKuQjb1THRRD3VeoR7/5DKAF1MuX0KhjdhRTH6WwMl8iXkoE1w7SyCurvlG/bG/tn
h3zupEP2LwIx2gihV8JfLI9UZZm7aU2l5xxmakKsRhgcJK41H1cdGAb4QJFTLu8LlwIPveyldjrO
FVKgAuMdEJhKsz9t+a1JdCwsW6Jo57K6r/fb/mhV0tUkynmigU5s7gNKZUVUN4ZtvLcVfmVS8i8a
gLgjyrHSzbRTFAMj/ENwlpLD0my9DUQT8JSmNTgbyVu7D2vNvOSXWjVeuRISmCncmQBswI33lUhs
cmwzrPl39kQuT9fcwq+jG9w+OtWqi0lFqoDj5zAF4zKddu22qlbVmFkT/EiVok/itVxK3CL69bix
TPSImHyyWxe17OIj+DpqjQz61tVKJXgYMKUP+Miy1CcGb/J6YRN13QWLtZmhXGb05FwioW5JUDfu
HKntQBeDvX4LYdH/0T8FstgC3/rU2nPfVEEVYec0ZTLznIvZh2gFlPDttEWDUiARthe/rGrWjNDf
zDd/c/MT3tNBlm4g/B2Vr7Ju3uk1l3g5p+xD69pBmHc/InEaHQi+JZWMRXevejhew4cNnIePhA90
kjJjkytkM0m6wrPFkX6UFJstBAwK/0S7BQjJS3vMBMn3/0ffDKFzCorCGNUP5YckbrQQ0B4QEa27
C7qJPfJVtoNlEmPzqQ/IcN9P9megoKuM1BwwT4l1I9uqHsilezCfl1bqwonTJUAlpgtneXkDebxz
yosm+tymjlIAjCehVUblQlf+re6hUwL32ha3sUwWCCJr800YwLG6c2YgakcTNa2cb5RDNxIcGE9/
hAFUlBbgVPK84MGU456lPixDaTraBmpQ9sEy61c6Mip3Qew2VbxgoXho+eU9XKxGCtAfO4De52ru
0uRS+YqX2NZXdN8kqSA6mrAQo2mddBvIoARcMS4rGfoR5rC32aXsNlu9zFJFb00JzM2Y0Npc9ssH
6vLeR2+oGGOpH71BJ2NglfuoQU5GpOPOEhAq1epgQ7KqEYO0jO+JFKn3eGTpQ9ebhhRc+9B0DENe
+gu07ibwZ/gfeKy8EU9QgVAHnEyMFuOkODsrmCdnub+cf9IdzwmXnEBoo+HIqn6qPwS+cKFOUuEL
QqInwTgNoKgwpfNahb7+qXUeTViq0thmswpXbAsiC49qKzRgdws0v9X5WSe4VB57msBZKKeS+9qn
3CzmIeOw07ITuE/eaGO4qTgctKrIs+vUpfVGyzcERtqMxtjNq/LSGj9Ptsl2gc+XF9HMaLdS2yOq
HuVEgrGiQm2GWIK0hSCbBqQLo4axvsFfcCeohtBUIfy9A44f9+PkMTGDAjHepZY32VtwUzAO26L2
Dh+dZ6JQNmoAJ3J+/Emzz2+TzX3EDD5gaU1L3DZ7ySYXzgE5SYPdfO11E8VEHJqpHz+jwxitBLkZ
dJLQilE8MSKH4IRn15KvvaB/OkFRJrcO0A1Z45Ot4oTRO1yy7NFGzCFCI1ULth05iqjYnxvkyLsn
sFiQoAY5Hap5nRUKn2Jr7+b1ZwUiNJGkc2HzNwoBgHqdpYvbSgfOIf8VfMIHoq4KSIcX0WCX+h6f
OZxHSHxcPhFuQNMqkptYHdRtmBb8Bn1ySxkvc07KR1uIy4/RDhC81gmLycFqEO9t1z8ka7qa7Rck
1YJVsQ5T7O3b7m9jNu3TL+sKamXdE/S3Wn2EsUZaB6mBrpvuWYfB+UI0Y1YJqocSOi8Jk/9Mc6Jn
Ro40cbX+r6HvkvtN7oTf4nHEKl/3lUlDCaMEsyZU+fDTyQ5/elotXtLIwaZy4imP9uaSRkuzlNMo
n7Yu5NJVQcuxZcnOemSQrtUyISe5ugHt8wVfZu0i/HzKdqVX1ng+IK3FaPRFZbVRn+UmIHTDSG+h
5sZNCmoE6oD5vRnKsHr9/BWUN4qzcZONJ6is66UJRKu3JpjZBw9yRhBlnNuEVeoRdY4eIHm/3Cf0
Bu0WWt3Zz/UYrZ8F99oDk/YLmy0Dk/oG+kRsfay8/oe3Aii6jIJdLqkow4hXwOiyScDLpjhaCK7p
ctcuEb5hs0wpwTw9LRWJao89AoeqgcYTW9amAAUMr9Os+VXxOV+s8LL0jVTsB7Ancium/5x/u4cZ
irH0614RSuo/W6phaXszc0mHs6VRltYow21pcgboAG1rt/XfgcGscQYfJag0IHBt5lcOVMrcRbta
YeofJOIgo80SBnI9Gqwl95fOUVmxGNDgsXNp19Ku1bsrFR9/gwXVMMF/LSAywMXRggX9xu5F72BG
yEHeSdxQB5UBTocx4uGUnl47/+MymmKg/whQH4jN8sk8KFNVPYC5vMCeiz4gJzAcw8jP8wDI1+uB
9O3OW9AUnFQpNcoItcldrcTRyQQTbTDu00uujYBFdgxNqF4fYxAs/wO2FKe9/nw0wnZTErdmsG9S
j5oXifjyWIneBPvQQ1GusGBw3+eJq5jmMst70NZHY6cie2V5s1opIEsnhL9OWdMnD6YF5xnSuhoE
dLYvFZxtfsORLYwIjdt57qxEy70IVIaTz94DBtJfGimqaCnraQgAfDWVlUMBtcqN3oa3KcjkCFPx
NWhQY3ngj/PnhLoC8rD6OjbLY+NtcMIM/W7y4ma3LMMwO840Fq5HPWoTY91EvAJiLxszT0NygnBG
sgoWMMlB0h1tEKkHqwmjAFjZLpqG7ZMA+EVpcAg0Kk2feLHfVxPCzezawukU6klYhMYUfmaSjiRV
KftvtID0I1CP3VZVgciyL93OHXvW57bXMjttBGt+YDj714n64w/xhMenD9ABq+G8rP6ZspQvtXha
CwH/cr4lk1/AyGnBGZxc01wL22v3sQ6DAgFcKDAemsuDBIV/kisHN6L0VySZZWftbvdIrnyFcCWU
eoUOLQdOgbz0ZAN7xmBUBJlyc3gL4XlwmFr54mcdlgkZ1QbxoLaa67Tj0bOavebRrMDGVK2kRsfS
HaUFML38fGd5agZgSBv9eu5IryIhhRko67oChgYQkXUOhG50ThzSNfp+1rBFVJnwPDUndYk3QbET
oh+fR0NQ4w/UHNZyDee7oHSXOv1NPhOUTqTZeKFKH45vowee/snc+69qsGczbC1LrKymlIj8prZa
nj2YvvR80b30K0pYnuuG7V7zLbld65tC04kHNbYXggIaHU1Zz8L/a5EotnzqOemOjXFDSGCZpBBH
JCUGB47GiiB97wvFo048ulByjST2x2TmW/vvB9v8wlZskYF8qrfjMNwP0u/YsDi9CN1lMLDGYAOq
9YNc9bI6TEvXeCbr1QOeH5Bj1M+FaK1NCjThc21D1mHLp0Oy2z6K4q65GbkjxOTq2+l8uM/BeBdm
3zLT/++/A2ciuyrjk6rmhoGzWHIk1Gw+JxQSLve/w8HjN78RniYtcY06cQTxJz4KYx+N765m6owB
d++CL10DPIUmxHnDqOgKPn03nahejIKUd8wfreHFn1UPYq3FyvixSRGdhbc5Q80FjxhiXfyFFMrd
GxqiDdEqVF9WH2UTPKlg+QutAct1MAb5AX92T5b4KaaWNJrvmV9tTr0tfO1ykjPczAoQfXpjFlj/
rWHblleORD66XiOzDOwVxrZdLgAuru5nYJ3UJkRUJN+MMTsQip00+DdvUaCJ1saPdIJPDk6VQzn/
J/aEO/43YZncX3Zkonf8cWF+gzMH/nzs6XI3PAswbYZtnbETpEowYgW8+wXRrtctekAgkvs81eJ0
pj43DcLdIFroDebfATCIYGvc3uBOV1Md0tMy/0H/0v7I05tcQw9PyldiIDRz+sJafrc2qtmEe8Q/
9Gb/oMfYJiGDPR2m4oAwk01BXtMk0pTV0i9zdRb+N+H2UwdNRX+k20u15FuKVY8l22Tv1bHCR5gQ
JS/mlpBhLDpktKg5NiNlS0B0PMFtFQkgQnqZVBrt2UdzYvt9141+gKPd/WVEDReGch+vUeb8F/JK
DSTSTKa7JZS/+zr9qWxepCxN7voPBS3PWN4w0SSPtysn0iasAk3Qh4oWK/Xxviut/LwhHzIqdfi0
AjkJeUyer6qXbeZFh7oiufaRDI7IRR9oDllN3RbPm/HUH/2O+shBkc8/gx8gien7IGDbGRSnPvLz
g3o/KQaGfFGuTPlvvHtL1jBtp2sNdWhTZREEds2j7Xa3ROpQYddkml7PU61aMJp4pulwaFmCybDg
1yCsFCg9tc7gvEph3rKRiFVvONvsT+o/RGVz/fvoUzoBAiAXzEy1eHvJoFyfIUJZKWoMH3n0qb2f
HdQZHiJQVPt+pklxris1s/noyprgSQ0JW0OUY2w67wqAE5REX0wX7WWiGxExHE4I6ZzlQXQjwxav
A4pcO8e8DvLGWVsYj0T/XfQl5HhJFkn/ScqV6fqW9l6+I2gaUo8bmLJXtEBt7C/qTpOdyOhuwzq+
HwzlIuFMg8JSIz30ju9hrLB7yX2T4lDuutCW7rYINVIG+XMl5JTlnyYA1XVDttLC7OUWhqMvViMU
OL2fWFzYEc23fQhkOLpCKk/6QZSgnZQlbLfWAROu012LzUnJgDqo6sqez4El2ymzHJ0EK0nq0dbW
FVzPDhcrsTnxuiMGgi8E0xbegOcKrDSzEie185j4oXy8ykJ6KgMjow4lfi50bHReWtMmFaDWg0Dn
nHY2n0knh8hNgxDbiZ1h2xxUnrY/I4agbYVgK00Za2N8qBSgUmovhCORPLyRIgrx8qVYPaHAlGKg
gotpsa+sMVkjULttAJ9a9fM1xyEMEo7aN2I8BAnpZo5KfKriy9SOkgkKomlpzxLP80zg8wQcEjsr
q1FNR9crJHR7ezjqI3tAQFe7UCXFro27PFLlht1RLJ/oLcdj6P41/5aXU+3WFtvz8eqlUc9UmiFZ
0f0jgVqZfTlOEc3l0Lls4bZKGMA7l4j0v9Ot5kEFnBY6tFskQ2uP6m1i+I32NWloz5P27w/gR4HV
yPLm4usKQT99wlWzUxFSLGSnaQmCE4TQirM/M0jwXAbuEIZeTj+n28bmbSGBeSV6d5u6ISFlubmQ
IhcrWNQ3lHiuVi7AzjScbWYisa83VptuFZ0j6FfXeggNYsF2ePfemQx38RrrJCDCMpPVV4vMbYHv
ULwEDFqB32RimA//BhfbWcaNpJPhYDIQrtHofv990OC4kjTxyLuS+vUojoZJG7z54wZ5z0qRDZ6E
QUfhU+EPAcgjzNnZg0cmfPlCawvYSuLKqtYBSs4BlOn8vAXFQgzutrAp5ejPY+yu6GWVrlTePM1x
z7Nwyp3LTbsaZLQb4/f1bN5/fiNtf2DVNN7Y6JvYerNoBeya8S5W3ieWCrr9AnfFHeqbcQE6Fw97
YNlW+4vzRnh4fjpnygDMoJRXt68XXY8i4YNnVCxjiJIqZWilMWH0w7X6BXbeEO09zDJ+4QbT0ieY
fKqgtgkVTHSpbiz1DhDr3Gn9ex0xY8HBdjA9Ac9mqDRgPkzKcz0UImMaHK6YIWU/zTExz8yugXNF
CsyxR3oZVcXGsNT/dDF0ExWMTsV1TifiUN1T3EFBlJTWvTU4M0vF4Op99BP3oaK9MNEzw2OdAG/Y
JnfhIj9w0eYGYR1Dx6RTeL+riik+BpOFMZ8rr7aZnzjx2l9v4ZwnhWeg/fKaNOqK2OxSTYOcYlzS
/jAJmsb++t3ydwweWsDtyqxi25aey7YkCbBtRD7ebvlfxJg7WhhoadlWCgxbiely2pap9nze97uT
jaPBv2ywxHTjOuRSDdHrk6lEtsCGr1gwHGCoMUbBrtYT3dJRzH8yDksKPt9MrPkONNn0w99enFzC
Dygtk+UQGTNzrenE2V52Yf3RuloohuMdxSfZvpVVKv4zqXrDokjUbnSY526Lh91tz6FPve0e0tqi
vfbU1EkLn+lkUjqg4EXwycf5+RhgVik02iGdKFBdqBEZqu1kOQMmC5Hn/VvPMcex5g2FVQtsWebg
wgPeQZyX/AI+Gur8l3SUow4I+pPHewMTfkqzBqC97rHQqQVYnXAf2lwMgjMjWhryA7kR6PlBLLJN
S7fFpzhQ/NsRDDyzws7vNajPIwJH+cQ18egSTkPT/aNsxJIHBN+NJBME0FdFO6I3Ytu4X1g8sh/w
4wOpE6qTJ9gX40b6DCB2cdCsnvyBt0T94VvCFaKIIL5dZ6JPsJeuFQhXfStXc6k1O49jpwmDKtEQ
HOpFvFTZxbzSeOQekk9afBmIwb8TKT6El+osMp6ZhOIpjm5WqaSlxgwuN5IfQZOwSKzn7E0Alxgh
VPFAakUqjuA23S4jL2DVoHQt8XYG3M9TCTUFsWVkDaxs4iEj+7tjv6+au3MQAg9sSRyon7fWLfF8
qnGthRoVui00bGBoi5Oc8KkhaftL8/kMrqziX/Ein6/0H9+G9gotWWcJF9j2HYz6xsLrbAC0VCGF
eaoKcE3PzC41bhM+PwQqU61wCVJEIFZoQ3kEcBGAh5axMSYN5+UfA9cAQns7LC4L59Vs4uY3XBvf
hK6GBLrHCM1pxjflnc92wXIePrO7MMjTZzUvaQfWdj0VXhtrwDDSTzSGn6kFXPlGwsqOOOjvbeCt
gkvaaWXeb0cz5WWLVRFUKRZlteJOqNOGdJuim9Dk5rghfakMmVb6++A7r8f5siYbIiQ1dLGoHVeq
3G5POtwi3pe2osUBAhaEOkXf09yjO9YwDIzDrtLyXicaFMxSqAeFVKam/Y6oY73LJkvNg3fpDQT4
7K2hori2S54zWUqA3lDI6rU1isghVM4iUplI3FY1ka7TUl/ombLfQWxW6WemZHgGQb94FFE+diDf
lCa2edMJNw9wvBwUgLp8wuyR27mxRsBsjkSXPe+w/xLaDOuZ0Sk2Z9Vuy7HDpKlYW/sdYvqoI1fa
A68dRzRNwPQz1JXyLPBtlfYzCM1VsT/H3PxLAWKPYzl+ipBzkn4zjrxFYqP/S8oWC8uXiQOURVnb
osWPMS5o8fh3Yq4XNrfyYc7x+dErytfAcvhCjB52s6A4A1wkJTr7zhHGfZDHr+ouPEXNy9QW1Izu
wBhsMmngIOUWhCzsz5og4XcCyDdAGjUR6eDX7tolTzpkb+V6D4HWz5C6U811mW5ICcTaeqEM6XfU
j71EPYaQwcu9qIYrC+xlRJr0yq7kzhzMj9tZqWVOcb7gBqp/mF0W4G+VDf9/Eo4quKIakW4dHqLf
9bR6ZM3A6fJ1hoIfhdcmAlsSSauVUmkxOEQAci2DVyB36jZK81FDNFccSRdVgjThnIzzX94kFnnD
gq/YJKhQuqUu+yR9fxS/0yoRCf1Fo5gFUqUoPomLK+o4XIj85goKmLXpAUdoofOkTw9fDvO5/kAN
AjZ4K7cQA+CdXhCN6BlvJFoqGiiqUOdtVB7o5/pVsY6mWgnFBHLFEuN1dG3wEyq6zhL/8HFnTFBA
csggBSL18AIcKqdKEvWE6l4dALJS2uugtpNeOCg1csYjQ12q9LNT+T3DHCJFyUkQFKhBkH7VFqNJ
Y7T0xC0lTi1M7DVbZxgOqmLq62hzL3Xpgw4zlxByxIfuDx4X4P7+OSiunY9SjT1uxz0PGSyjl9L3
2WQALLmYuTASoBFVK1tJ460ln2NCemOR1Mr+mBhHJ7K3shIPKPPVolZrFNSpKYkj2i2yOqflmmOD
CeA7ejViPZu8j/tWjDsWD5DJCtTFL77FWs2R6DF53qyI6Btt/ptUdwe4IaVZ6FTe7vFjyw62G2JJ
pR4TVmP51C70iOE8s/ntQe2QyliFFNASQv/r3Wh3lzqVwOfXVWq8quOLB+3WnPI+Mz+ZD8MFAMey
ZCIf+T2FNNJr+bqgzrb6Xv2CcXPXKh9/loSuFIwdoYdjx4f5MCGTDgQ3tnIXbzVZQwrU0ankUcsJ
zMz1xgVUtyI1v48SbQAq4Po9BFY5PfrG33yc0fGCS9Dfyf+B8R4J7Biku5eVo2C7e5s7sNGyhfw+
8JUEsp3zLjQrmUPhMZD/yw2gNwurrjivfjWyoHJLQ25a1CU7PzBlAu7YSX2CXiQaO7WidODlmsX3
3ryyFWQVh+faK8mdvfmGIaP5E03AZ96rVBJ8KW0ckpSOHqellns1d4KZ5KV4LCKThbJga0BM8fbf
b5fngGD2nwXZIX1CD0fFkK47Me4SpIritHrzHatt6vRROmlW08SNzz8AIlNArwwfNLznNOD4PbbO
3r+ojQkh0q7Av5QXo8jJlrvrYc7kY4tyUw5phRKrH+s9IdIrGv/Do6TVwGelw77dAb81pxuLlkKd
d0GM9UhWCrCS9EnyXNWOKcKYcy/xOun2Saz2c/Cp2HMuSwL1NhIk+CIu5jJYx1yFKEcdX0n6Sb7+
bi9VLZiDT+44zbs+vxyRiO9RglbGrTNZ0WmOwvUy0exMmE9JaW4vuUHBlZa4NIn6WDGUpmNWQ6+j
DMeM60Fj1i4E2cU1NZxAFzulcmFpKzZJjxIDp7djrB5A3UF0W+ZQAq0xohwnRtQgdJi2QPJOjfUo
sN46MsNJdx+Cc8JRePgjS6BOJCkNUMvbN46RHZzx4065L/0aMoAZo2s35rWxQMnKm/iwSkEAQjQP
XEMNu9C28lnzdnxhyZ0H9A1uwaNRSSUWlMwG7Tyi1jBCCCXHi5Jb5+Pl4tpPb18X7RgLoUO85bS1
0VhRVpfnUpWdWFwAI594zp6ax3eak9tbcJHmoebyElm+6l/fphvnToaUrGUwdVYGJ9YQ/1vgoDLW
SM5mCQdmcMS4jB3VwGeaUUhM4D3QEf7oSg+zZCcmEPM/Yjmcyz3ndOEQc+jj5m+GyNAhoa94YaDY
01sCLusIPKXvg9KdrYDZFE6EIhP5eBhbUmXu5PwelihQ2w2T54crwaTHSaOdJoWT/HiI2JdEeiay
KpE4JzDSmmD2HYux18RH/42xqyZxBMVsgcAtJjBPqKxdmdv50Na6Wnc7HErknzoZRvM9MFyrSOov
3ne9MuuzTZUDtTJ6sPDZZPYVtwykkPDDHIhyCAjk0BAPTZH/ZJU8Dspyl2irPnBfeXj4WhIGDFE2
hpMyjaUkFxYOHS5lObytgcimJSpb55ZiTOIDrgUOpULhGFsOt32KaDsiOqLd5I8kc8XxyINk+uRB
J3rOPLvHpxKMBWtn/P7YI2aLxFzvjT46wF9XayBH/ZCqHyQIdedGhIFy2SyU9Qmy5gxCxXyji2X4
ydcAIpN6MDQhhC45ulVHLzZ7sPMfUcE3qXnxXqBebN+l+3D31pb2c2PKjCgndu8gwbG0KSAcLjzg
170ij1kZiib/aCIHSQAvwjFkuBBX9ZUvQ89F5bVoeq9JJcmUuaOMmfR4T/O2ZCVWlz2U819Owc8J
OFM7lHcZFtXWXr9nYFudbhBFaS9i1DdfoOqTddsNu4DQ/njZdpmVolGiXU/g0rJYkLCMM3PCKZF6
4tGOXsH4kKYk6qGqAGbt0hOFfFHc9oUKJTWE4g+wqy2q6jZF52QRB5ZJJvBw2e7wBKLnTJN3C76T
ruHCU4GpztJ3OUdfet6/uZTiXm9JQE8YXnHC++PCIG00A6Oz6/tA0cWXZF6rl3HdAD6JIrOKSc/O
kxQ4M9IGGmKlIhBrTZYZXKB5hHpSuxXNHlEzVixv1Z3CW2T3fHWKeFe1FF4yx7oLq54XPwfqk4kd
D2Ky/XC68GX+utw3duWB8Y0/X1Z/rJlyJKm/BcL2spsEMZ4NSDOx46NQo/eG/WWqFWg54o7zez46
z2skCo2z9aT6M4lnNxBNkmY+Z/FF4KfTX6J9DfHOuigPUo0Lu3v82fOM6/OwraHYFw5+5KIDpfzx
jumiz/SxSiOi2/0aEcegbBfPWOEH8uzDsA57AfetmkhJAY42iPIuaee5IGP2JfUKcbbrybZbzSyp
a21+e/aYM2EV1oxFhmhcGn0Je9QX6KHrjZ+sdwy5/VRN9Dixqi/5qpdvcj1mYU9v/vzdUSv3fV9z
8GNEKgj0NdomouZv5KJHkbMwGul3tsa1AtbXW1qjVeQtd5fKezhDxWLXdNQ+HHkbA5BaqkLZ3kk1
AjrA9uLEDEcERbImk0Qx8XaLxgNEzG7FgMopatMdvP4kIW6RBY+AQoXbpvG5V11FE3a+6rzg9i9N
9MjUCLOXcQRlwvEavXEPKq0dvab8DDe3R4jjnYVoMdlLNg/ViJA51HxcJ9G5teLAdYcczLmTSN1s
uv5mGRYwWrNhXMTuaE/lpNWnKombXio9lCNPfZ6dlKU7XosNqERBJ+sBwsVBzOP0BjexRoE3wsrE
UksBrWxvfcdSDULtwNmSRYFjbTXgHv/dAn1Ea3iUb4yx8tI/3dsLYbOwWSUvwLCLNfq9fZsN3C7I
k9TF5OHmW8k1pczqWV2tdKqLbqouzgcRzm5m6wQpzzK0xY9SkA4NrnEmqvp1EPeUAuDXiMh0YPPL
SB19GkOMp6Hq5kPkfD6mW3nAr7rHilBMuaN7Jb7KCaOi/zB4PD4DDKMS+CC91et4NVNtenSEYZj4
q4f0D2HrLOb3s1NL0XMt5U2HF6lK1bmUgPGold1CJajKzCR3Kk80wBcOntUjQYxd6NMBA719VzMy
OdurKDnqBwe1ShMwNna7xnKbZMcLcB7CUnvANzP6Vnhg//2vVSQCA4OIzgoneWtPVQPPGjkBWLbC
YtfjE0nB8t6xIGpq63l8aZmTq/YH4MtB3TsvQIHt4Qz82N2WdmsCgaUjrO0kbOiVevXKevUQZsSO
l6LB07Dtbmd95p74Lx+pOnvQYt7UXX1C9iVVQ+sOaJOKC3dzrH2mce2QuacU3V5ZWE/eLtSGWDtw
Rr1HRGjYwHp//INaAw53L7PjceLwHR63wqq/zx67lLNNQxHmJNa1kqdYkmGx8HFH2i3SgpG+rrzn
TF7GADi3//UzIwaP7lQJeJyZyq0rSxumXsy3K4PqKWfJG/6Bmyz34SDNCF87qYr9EzjZguIgU1ih
WehGmyQU3Q1rojTEhaofRfOPtSNoVoVEvu3bjBSzpEpQBp77CZUZUV9a2x/ILhiVVaUsv0WNixz7
YoVcgp3HLiNPv8Qs9yZJZgA0aq9AjRlezI5wBzeF78OZnQ6TTwxDFP5tYQi2FTWYmzsdle1EPDyR
mE8YLY/IybUxW0a/8Sm/mIbOouCLZ3p9U63SKdU/tveic6YOGUiTx/uLADhedLfxLPObskfASv8V
39Pe3fJ7jjTXOIvHOIlinUpz5iEqI1pyv7RT69UgmBbLp0AjFiRnULdrBY+UNwYUJZfRLIvhKnG+
lXSJnOZCZHranKIdRROagkzpCpzv3XJF0hCKxKjnSj1wn3yII7lyw6QwzVhkrfFY7MdSDCvFxvX4
54Vm1hUbcdL/Fz0ZlFbp5WJlxfznFXuTy5D02wXcGNBEyhCcvgGQyiphQX8zBkI6hx3nJjfjlUkR
cZIlKteG2yQSU5GZ9VyxbCkkYwQ48o8uezNRFwwssO/vxfsCOy+4Ngg1JUUljXc4X/PMrIcM+v1O
buIw41x/DKbrX9OHunIAaSXBT8iI+bK5qo493Gt+b3z7hhM/DyUSuoD3fA8MBK1lFcBCmivMIm8E
xrymyzfsNBUQT/xneZRv/8Q/IEPTVRx9C4Qmfrlr/OknyR/bbSOProGB9JMp7aoAL+C1S45uFJkL
PdIJDJuoH+5NNd35XL1G3JF2lTlOOuo8x3yVRwDGf+hAzUpecGbB7Zd7NgfuDC2sr8kszZX2aLTo
4V1C2/mO63BjLjYqXzK5E3wdWwyyyiu+Q5npHJzvwH1o+8b+0gwXjKfte+uCCgkJ5RWVVbuUcERf
XQCmnhDGz8YQ8BkTpkrXSMC7KHyJl/rpJnO+qd0HQSJKSlPI3Xtm3vTimWXntixc9qEdXSbHVJLX
F2XjtPrXW3fxgpBMkV+nHGf1PK6s9WTjtzBGs7ZlbzeIdxmoQ6R8i4jQK8Fe/0D98arRKnGG0SOm
GjeUp4nbbRnPCpONU24TArwxk9H5x7vE6y7a44oVViaE9M74cU+lmsUkWcElk2j9uxVls5YN0IWp
5b5hVILCVe2LN679CQbpj8n4WLD+zcgCiv/Xc9yvNCiwhxUg26IARS77oBwFrgRy9pbGVxAoGKmx
sA4nr4c07DQaD7dF3JhomNkuFD5zZecLgMq5aIVH3gB0qR1OOfOQMDd5S8PSN1xEcdMPTLer7Nmw
kkHI1RE7dkjdsaKixrc0XSQ7F4r9APzPt/MSA/6k0t3HxGvzwYV4FtDDWY9ZqSdixcJpOjf2WB33
A+0LVKa/Hhph/1yEQ63GAIoEpSV2vWxf5hUNV71hrh69Ruk8eRF1Dml0uuJwlJQaKhHa0Td7Hk06
lMueBlGreSly4EnmgRiTrvUf0xkf3+tshBpTwwsvOE70SmyyFLwkHqpifzk2bXmJMC0HjTNvsyR3
x1kVUCIWbh35ZKQdkyHwfcSTDwJp1XAJBCBUG/HtjXw2ACqguXz5F6mkkIuAbcCtsm6z75p/2Xea
7cymxPO/aPt9Dy7hNn2gIPi4IAjvahxCFtfDjPIDZXU9n3Xdy/t2YNVqGMKXQfCjIvat24sZ6YIL
uyma136XdDmqt6Li6fKe8bCK7YNsKwU3uPw1iPAlc2ZeDbQsgbFTcEscA34/CZnq1iQ+K6zj/Hpl
hV8YfSB6mCAuZitRv+x6AaQvbyB22Ntxm9Z9XTv4FJZ0DUeCCtUZZ4sDGrKPYkOpvBot7BHmLADt
dniNVE8eMxQnHPzOM39UTmQNs7z1Ag/jMa6D0ze31XHhDg/HVCWfYxLyiXKurzG2kXaDsftaLg6U
EuvFTxybLT/bFRfxxJBpSRYw1j7nDdkQdwXNPDKMOV2H9IdPa/mCvmoDkzg2FZS2HK5hQUMlQmdh
0k4f2iQfmIHrg5+pZzkEN7m3R+bhWoP5YdAgaEYIXz5qlkezY0T5EQIwJvkUvjXsl4F8Z1USxH6+
D+Q8nOyiXZMcXXaRLUNWzThitaUAG2ZLP1h6xlfKiwaiyCHIygYJTh+t2fzF8DXAPbKRRQLTxtoT
UTLH+naogc/XaLmXcl7/eynWrvJeWYbTVliyIN0qaOww+g1BxcFGU+yP6DIIBgP1KGN7cSWk8dlL
PyodbzkE7gPYSM9hWLrUoS+QIO9RCbvo8qKuWoNIPBoMNT7V1K2BksGTECgSCrH0jxH0dRiclArO
wNEH6ATM58jwW48Kvk7pHjCr7NXibQ0zVngCVlkHJWenaMvZYifGPjphJDO42Aq//3bJzXvt6W2f
60KGZXv9ywjeQf9dQU7j/r5aJdDBfpp0ntHuPsBmGklJBk6XgkzelCPinuIlQDbAwYQuAP7Zr34L
dEk2XY85I9b5XHuosFWuU8dkJ1q8vF8qkQLXpcbp8sKq7mcia0DNudp3sKS0IQY7GV0lBXga4t/Q
vhcKoEVe7PiDR8swHIicaTd+dcZzmMNKdzaQwxdbD/Y5UPMG9d55nsE8v8L9zQvgRICYFwgqkxQq
H16f2jM9yzXa3S3ileBa45XPjMNCKE//pgUXLbF6ELGRyWC5nxOZK/iuqwLzpsgT+X0vmYM/EyKT
rsGYCu0rTdqQTJakpH/7lWee3VovdgxH/+7k/hv3zSsvlEUdjeAxW/7ZppsAHqIEdLm0VE9+cMGX
sujU1Cw2ww09qFvGBZIMRoxPACQugI8jy9YK0A+03WyvuUOHmPAH0OodZf+6A50uVRvMjERRbhlJ
sup5w/ORjBZO+caARHtdxuJ1CV9GLcw8YVWk6Tc37OhL2T42Z8XxPaUU0FRu20vBgs0UD61sXICH
CBNrMLX67/TvRKnUYYZzVvdAwg/qDZLJGCDoh7fWW6V8xBtkJ592p6ZGwEkJ0swav8O3z6joDVu2
06Abz3OZ1nVFUwdZQnXt4gyV7KVXumQE4zxWoLsZ4FFZu0doCOkPp4ubzqWg5qpRDpl53KQ9zJ47
PuHkh4rPviYf63/mYaMRPK/Vbjehfaf5zoSRbIv6d65b/1gA6YVo1cnetUpS2SmkvxA4GyArj7T4
HRbyTquapm/YQRV6XQcJGcIkYxvYCkHkkwo6bhSLbXbH8omoutGNm9VoqX7hamMXJEDC4vMtr++W
I4UGniHWYRH5x7R13cBjG9T8VTJRBEqqcpRewxvIVddGfoZr/GV2NiNuCKXx65UwF/9cbwrcIy6i
Lm/HGOueP951RvMiqSMi/A4+SKgU6WxMquWZ/vpkQkBS6MTs+ESdU/daCp5WNjJZUK17h+4OyqpZ
PF9+fQ/xtNoVd1BAexXz65NwqBhMo6U2IdSSUcTJayNYSnLBR9mcUdUvY8u5cAJlnjzKdbAjztMK
xLlvejTUCGU6JW+CGJYVjdAj0sypoSD9XwP/SeSkEKCu9k2dKzxzQr0wTBF6R+y5ZJ9cxsFrsZpa
Str6cBkxhhclqWOhYlAE2X4BnN6ySPTQdN46gH9BgcuxBQnLUyHn0Hve6yfr7+/pVo3Hm1N8nXap
XcKFEsvRjR+oXCrsW/WrnZmKysP1fvhrCpwko6fEA2qfRaEz9HCqH0oXc3eBByJjrlCVQPXWw5Y2
zl2yUJNqRM+ky815MZcDXBl34wc+5hxdDuFO0azjn7t5+/DMf9Etc+mTwUQBbNsJL9cPrZocSON+
Kd7hCq8ZA2YbRLvKjSr4KmuQsPLZUuoxsamZcMax1pKt5GCGOhsrcX9ZFj59aN8si2l74ucFNqo1
eSTLpJP4H7zjiTso95vu04Krxukskz3MuRqC8O2AYvRQbrairMuqc0p104YVkstmUKGNwg5+FBvL
kDsUNyPsqmJlvuzIjB/ScjyN6i6EByx+q+WdWVVlLcOQK+oVU0qrvWjGz+IT/GTQyZswDqXKEQB0
OP4d+Al4JfhPyhoWiSRDGuc0lHXFtraencHEQZXGgs9nNG8NwkRsrPaJ2jR7RS/eAYP4iJe9OKOB
9sTbLapzEUBgDw1lQOOhClfgzul+D5xAo1sG9uh4KDPRmFqdJ6kDbZ8oGwX7A8hL6j1TZI33iS0/
8YiMHDlKYv0AQM0UObGeID8CaNox+QxHgrZgJx+zWpqtFBz5SpG5uSZ613Ruu+QwBis4Da38dqdW
XTLNKb7QTzLJmLdREaO/ieLVrBTfkWT+3KNlNuegpXixXoy4VaTFJgC0N2+hMxSNmbOyTj8m28p9
/gP+926Sp6yAXthhb3y9c3K5oczXhDb7dhqCu+z62JmPRkRgi48TqEkyH04tM6DD2QR49HbZiBce
HxJlwtUYVfzx82sfCPSK6JX0Wxc7NVC4AzjPxZ5xVVB5OC2Zc8iL+7tKb6meWSCi5wkkHso9Dz0C
SVFiNbG1DPr8Lv0s27kTKSxtet//RZ1gYknP5vmjsXi7E3x2HPCsHcTwyfuIzt++KmFGrWBbYe2Y
y889MpVGYPDbvzQk9p0Afq+obXk/lS0p/jG9M10NjEfTxUAGtbP/FwLDmQ1MtwZ79Ukb3UFNE+z/
53G3teN3tecMiSWKlhmJKStt+RoECSL4ytfNna/nRFYM4T9TDruZynFNQWMNTRd46SiHU9XiInfH
EsWeSKDURLrcvK4z5Y88yWxo/YwhOajB8eE1INCmiQGEVX8JrBn84uGxzPphmNo8/RQf8aQBuGnV
lZ5GLP/yCJPCe4UGiIWpScXRUpkrp4lZ78lnUJY/wrFzVSASHFznWDwsTMRkEiI7dWk/Ap/BBDOB
Y+MySrfdcy7eWf/RgW9yWWzmmnufJXc/2YyowXNOTqlHRzB5ARaTZ5yOZZCskMnuA1Fu82PWThgm
kYfHL0qr2Jh5wRX/3IHIEE0wxAtwrdrdDOWl56Z+SDqiE667jJIB3gzRS/TaKQEb8bBwwWDTRAIP
MOo9AYKYN0kfn7t7AZfj+g+eL+X3hQzoVzmyF1YhVRTGr5eczb7A2RvJAECG3/5EgPPk1iEMxuEl
EsYPSkmyqK54M9NBb/8cJDx6XRv1IfiGwD53PfGbffx7HQYtm6i8LEEdRBLmzUGbQl8aVhOdIHJF
EpBi1U9db/7dnt7OQQym3lq9DgqXQUfYSaKDqfTFgNMav3ovCVI5ZVeTLpsM5wKxbpR+XSGtm+ty
J7qDunPOUIzlnE7kokD5g54m4KaoKRMZQcm+vfE6HbFaJRmUy0PSLjRwBbxw5esuOgdJusFfoAKZ
hFSzgc2XlZ2N2OMOm3OJk2pdlOw4u46RurARsTAzY8/gyZFrb+xOzVXKUE2WVenOd7R9iwT4bUhW
96vIqxss5737vRHD90EhyNSFtk980FnuLO6BGLT1Os9i08wOtmYpVzlgFDhK/m4YN0LxD1dFNu28
eDpgTYg2GDlRx7EFyVQ8WAmVAOWRTvKyTGxpDcJAEn/dGN81Yj0kw0zDAIgFnMIRXTpZ5rJZFsdW
0KqVr7UDZbXg8/UGDPEdnpjbVmO+hnU07TxpO9vj/y1dcQmnDQS5ir3ZwOpU6RildcleARKS9krS
gznPIVs/w4PvAUutU17FMfwHsUyW5UM+EoPrtdxnuLZQz3jT78j5PcFTx5kScbDzY2d25Ztems5r
FKVFCaH3+N/BZtM116xU7p4oQ/DrMtxhdC+LJ+X6XwBabE3QMHWqdqtBCFwWoTaI6t3/Dm6//7ZA
H5sPhNrLD/W34UY1JPNQPaCqSDgTukRCJffv6Kb6mk2ooG/uShWFsCquGRVTyljZ8GhngCMczhj1
GD1/ElZ7E5sJEYeo3590JLcVHIbN+PNSO++so/jBtzmfD17GxlkrEGLr+H6f5RIPTNUvzbwioKgz
eUcG7UDzHa9GZYZH/wTNVY/Ws/M5pvHmfwh3iz2l0rpZVUsubky0q1ExTGkY0tF/rhJA2nsKBy6e
wI+v7JmCR1ZV985JYMx1CfbgaAYWaz9wsgYGhxbi87Kvvr+6DaRwXYQmKroWySNxOaHdZ0VFOQ+E
5+5hqaEt6iJX9BjQKgYHojrlFKkbSryScasNCa97EcZa7RQfKUZacUwZS8NbRr1LZN+fxbYMNVIE
TN+1361mjREYumqhLSzgohIylBitrhNz6BjP+FGAV8CR75DF+9c+dpIF7aLtrdyMcQBZiUkR6u0F
JZkm1KK1tffRO3oVKHKwE7NAc1vzc9LZ8OtOl0JHCwd6dGRynWtK2HMPLFZTMZ+LNIRz1tHnb42Z
3dyCK1Khl/HZVs9ewRKVcBeDbrFZYHXa1KpYPD4MdMCrJNewi1k366JAGhjlrAnep93bxXUMtHBb
1bQruBEYdLbiBdhti9ESKlq5P5cpQJLXudj7Pq9qhJAVpdYvCPOfFPJOHnnQP5dn+p9Fihphzts3
jgh0xUEwf/EUY/ptHBB8EiRsTCUgiP+oo68Qa8z8YbAGJSDpib38Rqirb5CS5VygBZEh1FoG4tWg
skGGHY6f1oDXfFZW0fK95Vxzr0X592qTu6Kr4I9vnbkGbdmvRSiRvXxeRqolk8qKZj0WVVSHPTGY
j+Gy9yHjqpAnmWmgD5MudERHg4ebb8tjIuyb8NUyoQFkJICl6k0wIhNONlqNVRyCMfxBYDfkHp4Z
7tAJfpgHS08xpWYgms7li1lY5jYpc5sIxtPmwhrc1RmE5TRgihspXr0+H2IPj0TtpPj9KYpV2e71
KknYHHNmJ2f3eieVGQiq/e7YMIJ+ULWIxvE2omFQxqJf/IojdM5lwSFoXKBwBhY1wqOKLL3w/ZjF
HT2wWlrZMAm71e7OWJ4clrYDy3VkNFgSr8K5i+kezZVal9C7ULszYzEGpB/MY/FVhufyVVjmBHGw
SC4fkCREevQvlyJ0BgCwwkjZVryqakmWw0+luQzdcgdJwZGIoANVmoIfhBL7lWUbF0QV7nBNYaMe
BHurXSj7n4RfL3EnTSRspRk0gEUzNrQ2+H4xW+fQUx8MfnSA2LH3ZxM4t960jVQZuW7bIQOwDWCW
xe8IZHHxTINxdhfasHsJDJF1QzyNUX0vk58C+gtAdDiSlgNbITl4HzoLEvSPyyFvHfkyinIAvEc5
l9vekotojEx49hi0Sy4aaZ7bb1AltPp20Nd/fXWxHw121D/3nRQwebFiveF2cH8GS3+T+XBDvHAa
vCxYidmoHt1J3GzxEPL2+lpIwXSLUTfSEnuxITYNd0v28Imd3+KZwnhbPB5Ghwq3Nkg9ZZ2tbb56
FqMQxCJDx7KAhORNpdhEsTzbIvPdYztiqoeitxbDHskf/kVE5jAdst88z14aECFrlpvdAPLr+uAG
Ldq3AmpXkuYPqOdza8Tb2Qk0s7/HQHeX1xc2JBN4leIQ7FLyn7e79Gz76e/aJHp999trKs0Al7vk
9kbNTuksJ2Qhakr4ix4bURleoPTFLFYn7LzyWitEd98z86ZrMauX9QMfu/O/IYre8AecZBWki+xi
M+yXC8NWPUly8UFUeHw/ESjolj5nFNR5jBIs1/hu+mjm2f2WGqheCtNw/KGQ8z3pfBFRXCWrrKxg
NUfWSM71OycrvPf8jRGjWpMApEiE8MYffeI31V1Pb9wk05joCTaBEhsq6ElnZF3x6f/nGZWgl4sl
DqSj/CEewXiXo1KnK9x/DOPhu7isQUJXegPTlUeyWsiWOJ12WGIDg7T4DKGvZaIsNLU4q1vw+Wr3
WKSEdt30zWnBeqKdUvEwZZWYWN2SKTDGRcgSX2UM+befVlncBR0LP8ix75H5yaaW85EaOrNbChVP
7kDjN1rwqfmrQ3gEKMWvUyKBp2YmbKOot/ucME9XNhUNm6CQmhOkNkAXakKq3tTDVfi/y1dB91Q6
gvYTMO122OQ+dpNwqnNU1KSvTQAuEjgwGLuHP8j7bpQujDVZCg2sC4aGGlz4hxLG20K7N5+d4YsR
qEd6feA+KRtZtkQSf2aHVd0LDznBjxWhizgnBH1dVUNhMISYQmX6tUmWVJiwjNBjSf9NQE2nvZEq
Ws1Sa+WeME+at9gE3TeQtxz04GvRgULeZ7VnGcnNlUYxOKMbQAoavx+D2+ku9GjLwkFr+1Gtx5jh
UVLPjcUyTq3+RfOQslLP/bsBt2k4LAv7XUC1sfhmsf2cX7PW/MKnLnppY4MVc3o9yAOYU1678oyz
B9XU+g0qX6oQR07egsf7jdJbmRvQML7pQwi9ftyFDgu+0P1CHgr9fSyVUq7fSqo5DXCdxJvsap3X
ozx6Px2jSPYk7kT9tf9WjsR+RzJhzUEOFLsAMpsEf6k0dRYOGoiBSgPjuYAKmBMhoOgCI3lzdgkG
UgNdkW2eBB4zEqCgpNwzI2KlDwQ7G4BTpkioen8q+M/npUsed3/R+0t0KNzQ6e+cKelDdnXqywQ9
AsDHqLasjg7QAnUtTJ7RiSS9lGnKLDstoYOtZUmNnvUHWa4WYD3kVJROVS19lPzqTsWsFWtCngQi
94pmolHuQTPQxaL2X39kbWQJfjYVfJFX7VQ42VNApkIZFW29AW9bkN9S5r/I5dKga26VZinn0c+E
cL6BmxQtCsJIi+6NBPavlKP2xR3G80eCNmY9M6DrIm1QE8XXps5R+bXbop031zJk488A9sPXjRMN
8ks0QbuEOg9CMVAttWCIsZZllLLdkZ6J8En6n2KgTx9BK5+8YLIm1CkTTH2EtvKGyBDQb6an5+Cg
tvBX79xk7+X2/6LXl0+5BH0TC5e4qjxdOJZKSQ/SctVRmNwsx8XtORP3nUPBOp37c1XIzGAxHWuO
llvYMsYVyWkPIzsgXtww9en/O4OtuMAKkrBQUMa08JupKm60ZLDKuH6twWnhbQRPzq22T5V2b4hP
THZ4j4lamHRwwE4Y/VkaKpWUqNJgQg8c2yFfOHcbbHbGgrRP96zGXnVyaFcD/m9LCaQSKd1pBJ7u
wJkIdre6heYTopeyzODE2K3QEzWRuSm3RRhAO2LzCsT/4qgmtel/ImQJW/mxZXq+Hdi4TVxYPe5f
jQz5zQkUzlB++kDgcgJYSyqX6ZLy77u+S3iIRFn55ELjL7F+E56tLsXgmjy7XlunK+IqNKSRc9Hn
Rkfs09gFQ2v4veHj5JyVFw+eQbucVXU+t4K/ILRoGmJ6TkSsJDUYjFm5FxsQEtxH24kQioU+dDPl
Deqv4PgbiwEmo7Z0dZKx9pAXQKE9atoLyd/MUq/1ScOxPEYuYs1dOvEGF+scuBunQFDuw7DjCCn6
6ZSHiF3wT+ig8d7O/p3UbRlncAOg//WVXir7vP9mA8BNKBRWfrgDA5hwm9e8kLqfCX2OtPnLUf++
87PAqm3A2y1BsxoCiR+QrDMU1lz93fF6jM1SYq9RbpehI72l+0qHzfdtbrlnw25rsdKGzY5vOf/C
gqX5OgZkRkYEsqFNqre+0+HkXbvIAW758Jr/JyUhExndA2FuDOTqAPjG4YNqcYmxpXJZrR8Kzkrm
/B4LIectyCVe2RQ3KYF1J++yeHkk2/ar3XUkUByXLGbi5r8DJpJ3+aYN73Pu+CVtkpaPxXUb93IQ
vJveI0xHCN+m00FBvQ0R04EhaMoDlN1tWD4DctebAV8DdogvkOyxpMbVJ1wc7ridPqOCaWff1zpV
fVpRP3got+LQVQbvZFX4hXYf03A8QAnT/PB4z97hVb9HApIMoXCTk8j0nGk24kPUR5w+WeWu2zLB
6YL+7ygb30fxXdMpp1JjTlOyrPv6BRMzWSPY5xNwhIOamcrJXXeUYk9TG9w0NHByUlBxVK/HGCsk
nTs6hSI8jt0RfWYmIooR2nSE3T+yc27J8/d20YXuCw3OBy8nap2flAoHXTeiJ6BQ53kYlFr4MO2o
H0H0URoyePWRSSCGE0ytUHdg7pnWVK1eLeUatl7bIZS95sviIZNZs5xCbBBvODkwFYl0Y+886IZB
z35uHI9MkY+LIe0wVRPegZvwW6HPrf2U/BaJIf/oMpSRFJZo5/lapmEzK2RlypAdzdxAbPMEwWEw
RpJISDVpiR9z8w6RXbUEwA1HbUhW5yHsdbNdfptTEq7iEx+JOCjmvMI7L1uBLDpSwHWpIbdvN36R
d7TDkTftsypcpxHwnhLO0kiWD1ZdKv6w/Q6oEXGEhyMOxRLB5xY2rchHkJK3jkhyBsH2ktK9yHjX
ba2fDK0e45+XOR6OQWHwqyfqx+3nX2EDa+v9wy1qIZqBfm+nEulWdvZBkaQAiy8SE8fuF0S/Mzf8
hfx5GeAGuuy8hmYai5oF6G9HvcYFRPRN749hYJX+DMhFFX1gdX2WpVfxTwwYTZL2X9ihC1+nG1Uu
PAshMFR5llMMK00bsEU1QRwOXu4ItRubIEsVojoKWKerKKG+aYFIVfSYcCaumPOURubK9f40umxM
2wcEC8N4QGpEBq7028tMakgRVNGaUJ2Qg5G2Pm5CzhaOCLhkct5aMWB+PpjCMRyCt7aDPucs2Bhf
LBEwZ7cAAJdEkFwrg5N6/TBJ15OOTUCNIFJtMayLULqYJcZ3WLgcpgtQQ6Fn3YF/77pBAqIbI6mF
ZM/u4iKvpcsRKnC4RKiG8zsbpwMlxiXQvqViSRe69scCBMMzxYlfZuB07R+zY/Fv2fY2thx/7XHv
FwbkjxYzBmb8kZJviyissgcBEqP8PuRLc77N2vjLUJKeGWdKwVUtcHfrfejibDyGUKQL/GL/T9eq
79CVbdqtVVblnkN/qLn/OMR3OGyg5HuQLFSpyTJpOMDUbNLzhKTehQZlkre/JWoLI2/HRhF6EDOg
AL2eVPeTfn5TJ32CNAJyrXucLfmmnp9FEQ9xohIqCgXAMOpI6OmHFwjwPXDCHn7CwcWMjOFvKw9e
M06PHg7vRzJlx/YjLhse2cbS+d6mVUwIE+TlhTvux1jsTyDxogUevue3r/84X2eK12Muuq6z/aYC
AqMdQm6VG6Egc9H94ItW0oDdP+DOba/EkyBsERDuSgcU935r++OPpY9qW6AWiI+5S3pstpL00STe
3gJqsVKEWM/0DYo/OL3D7iVaUjcfDGZDMgvwtRZTUKz7MFCOtYbOhZb5IL1IaRYM1KiDTz4SU/3M
JSCGCcEgOY0N0sjeO4SZvBe8bTOb/kt4VGbisZc/flK4ojbPMmz3+uwtlWhpTDzUy1i/800puTSV
0os4KfxRutYX67A+NXIqlPPA1dvoDiwcY5U6tRumVOHvcPBTYMOHtq/zhTnRbXeG5saS5G1xtc8e
OrPkyBZM6eLoBid0AwoM6YZT4fuvM9UTXAG7vs8JpV4PrA8rqUZOPu5jTHnZoL+zTv9Cp3mBwIaO
MLnz+E/sN2/rX/Ch8aRwTHqOMv9CqoWt3vkp86fjPrRfIyMk7RY+HtR8hTNudo+DHQyP1J8MIX6W
s3sfMmnREcTzFYFEk9cV7sekHBki7AnqxhLYoADonA6Y+XKITMF+TaI/1ZP+VuS0VQTo4uFF+PPj
J2Xzf5FhXhQxpX/NxuNL4xxW/wrHO0nAULKrSPUQ82hXCDHKHqCUjsrNpM/6xUB0MAB473tKTJ6O
uKt0nAHAriERhxDB1pXtl1LRIlAwXny6kYzZufY00+OdFBuDC+4vLei4qgwsVOP/6tSoYnqLzyQO
AhWMBfXUyaN9pS6Zyt5xkfZmyc65DWfCoNT6yQYcYyJrN1+Gu5cZt+b9O2KGnapUJwRnLOlr/FAD
oHWOoFgek+HKdded5JtoPVyd3hMX7Wk+Big0KXsrK+M5bGcDq5z0m1Vh+dH5Ctc2v6RfB5HEktmf
gmpJZ8ftDAq7te92T55sf5egcXQ3W/20y/Gh6nyOfRrHH3cbeaiSfpfhv+ZGf7GWqzfCR0o9P+L9
BePfNILL7vBZvBJIRTHL7GXHlI4O7DUSRHiTBCrPV5G+mfKjLN3Sp7ikXwncr6G/5DYRTKyMIuMV
0EZCTyrstzrD8TjlFR/BE/nyVLH6gO7dRUfTTiRKNqrkDZeHXe/qWXvtZiHBwMVVGA0swSaLRN8h
bNtHGL4t/dqcPz0VcL1q0XuVM8M0psig8R4oevf4/VZcpnO7AQuRjnO2H2+9gpNbrxoDUInOqxY+
DdYvLi3GIIiteShdp5Q3Dn6HcfoDBVwGWSoYNVI66NpQY684MkoVVzNOjJKdvzD8/30zuxFJqfeg
XlDT1NxKkn7BLqKLUwmjYnNkczCQ7tHz2h6lA52Npk5Mw0aDlLQdbTVKLmAhVmHL8sksvHP1/RLh
adB0CFc7gfBRbZ+1fLUJX7Nx/3Kzgo0ECYDkGxc3GSAOAWuyt0MeJwRUjzgP83Np2b6XQozx3R2U
SNdRGwulj7Imldk7hYjd4vFrmak60RGdze1Ko7qeswYNKaKKSNuBoo+UQLcwW4ZGn6ZZLHQ7eM4n
s2vBEgKmoaESuYNH3UMLjwkGhT80G14MOd1T6qSW5JCjqTgC0CDwQOcLye4tHmBiHzSyfG7jtO3h
RFtAKN5kAKQ0Hrhg+WbL24iJqMdBtzL0+JyX2ndD2YVDLl/YvHjyKIvRoFZSCVVQiGiSLmp0d/1g
JdAh9bPg6n7+3YwqAg0wWvp8S6HRXd+e+yXC0VTTRmmhfS5pbCihzGfZlYdMDeXQZz1hFdQ292Ue
ylICYvAIyog3KnWguhxjnIXzrxIIRHW1U9+4Iw8nsKe2d18co309lGGaQ1zppR8/k0hf+YjNLVFB
o17N0ilPttxmD21cH2MRa7JU7G7vV2876t4fUM4JO3nt33VmORQ2HAcYNui9kiRmud7PHsibwIYh
7Vn9oLlK5TyO+sSypTn0vz57d/EoBZYdpM8QqQH9Vq/lhcSADAt02rOkw+jj1b3nlHMoCTmwYlK0
hA4Ckc5TJPrw67ONc7FHqHXO8xlGXu+Ft38F58KrF+4rEOcUMOecMHmAKs7yzExjUM6vORabwp/D
gKhKx+3p03AMjqN7xuDj64QDr14zTpd3gtg4yMdUFf5H09HqPJn8o6C6QeMm/1tGM7tHtlqZ7aiz
r36qyvWZz+R7fZ0m+qdYGQPCjXllO3oLPzCtCDOe1FdJihvQFtvBaK/lQ6jEZ4+rP7JfnNoUnO37
W2pkvbLTeXIYM2MxggHrtfYF5ltHFpDSaYE1iMFqrk+gQE3V3isWhBcgkJAszps/MTcxvbFW+gdM
CpsScZxLCRzNdOJZOR2rTS84T3Z/PC8qK6hBF/9F7U/IQmyRYjdWLRBedod+6Lb3vG14LMDHxDo6
9uLxh0mzmpYaZ36M0J0ZrNwbuNkESiN86CUmxJErx3RysiwfbgXF+7GYR2CMCnEyXpN8ykLQ/hzL
6xMVVWuUsZnwz2l4JafCos2Gb1jY/Jd4SisfgVse35wCmols/N4djKJxJZXO9CUK8p0ZLSfjgrZs
uh26vB/2aUE7MAKolotrBj4NegbRHllVSdW8A6oPQDHKLZXoSBkim3dbrtMEw3CDRbEQMdSDdyvn
JxhxDZL4r7Yli9mqVK7GWt591H4LxTO3B9SJ8QVGVHYDxLodPikcihOInUZXOZom8q3j5SHt6gAG
OvL3U5t+/tz1J0zOn+7RghtwfZr6/ne55afgBPEcRacmS0jr1JS5us6+vQNBATIwEvZ58QVASZxH
ZL70vHH4xZjrXVCzBmhP6QxFhOtOQeddcYbsXGHBhSgzASNVcvFqwa2lJOTqTLlckuZWi2wwNwgE
yW9qOz32lEBHde6OKRakgBU/rbywUPTFq0w5ZthcN1FqLaYytDduzOI0b+iW+wixJFXc2CGGATlo
Sqmt3J7mVLvSyyGeUIZQh+PRVaOcxQcYHNm7aBpXmdSNdthJBtGrgg+BSJuHLnf2v1IX2ANARuuu
3XIncKPKIL1WGluu7/sLapapeyM7VxxyayyEjS0BdkSeInU2z4Kcym0UwAvbdB/hchPD6CwJHttz
LigUYw+LXf8iI+66wnXgnlf2gFfoxhoLO3tR4a2YPt5qk1qBdaaDwnTeI/CY/5OwpBVJvSAGOO0J
XTXtvS2GjvFAERkvcE5kUIh11pifzW8Nt9W3PW1WHgMgFphXoJHxtZzbeVDWKm8GxyMP80u0kLAx
8sl0bFZBZdHxwZ/3qZv2LMxK4LoAXUSKfh2MtoGIbS5KMqWE3MPS+tkfuOUhmLmBK0HkTjfP786i
tOLfquWGGO/gHBvy2To8HgDWWlT2LblKFQogTXIAQ8EMFJc0yVsO1P5s8FGmUUVRZGODe6BTphxV
3JrhyF8MaPfuHT7XKvopgiQ4jkzmJ4XJI9NWZPdLqSI2Xdd/JX47pcBIOjoHLiFtmbq1TFzc9nqU
75R4QWfNJtAtGrcl8a5J2D99JFpJ1UhwgvdmdqVTna1mCUpRLYYfE4UhjBwUnCoUQZ63xiP3wXqT
D3pUWzDLnR79xB6G4qMEvcBoQQeSalBse2xKyWyntOJX2ZG6l6sMeDuQ7oD0eJoJ/4xwsS8t5Xig
nVej4GOwy+S8j7aJgq+vl/VjOPWcA5/HBDwbvvKIFLwm5YGVAKO2xGC2Wc6KlroUtEwKi//SAkJm
6qQ9IS17pHEam4LieaJ8B00Yp0bbiGb05EJqdeAYl5IF+gvTbm/iXEnu/5qo2uSjlMOb+6K3NiaR
dD9rzwa49fDB9ozGN9oeUOUwzXVf89B1Ji4SgXPIlabVR6DImCcUdkuj5rG5D6QKE9nbaXzYoev5
UPSs5ztqjaT9Eo/ISvHYcw+D/GTvcx5jvoceERaStB+DGjRiGjeHIGH4gOHkKph2O00vGwen9Ej5
0e/o9kEZcSBOSW3mHONJyTdNA4+VOccCafBm/J4xcwPBdI2G31WGs7+C1orvBSD8H0hBAjidQZXC
wfRV/MsMdlH4ChM7m1J1eZTeeCK1o3dxPh7mBB+SAf028lFEceU6NKSQTykeEy3FH6dLdlDAf2+N
tyxWHbUHSgs47FcbfDzewT2yPPkyiIkYyCl1k60e6DbDZnPYZRFr2bGPBWd0XQkBpExqCnC2dfru
QW35fze6s2JfgpN/K8sPA+WMAeGA9LqDIkW8c1IYqC9zcxq2YsuCp1dWFquVf3cqhreK0HIHQlTV
6bcQQFPN2qMHKAlkbdVx/HpY8GXVF41y5ja5QOLI1TYipy9CfcxiXiOq2w+3ORXtkk5BYUyFb/iK
cjcq8SPbATq8UMXIhyJxm+ViAWrjN42cbpsYDpdC25puSLsQ9uEEnws9C0WobrzR9CtjDZctm8zk
jVzZANeM8JhxDxTlRu202Ws+4Fl/7j+38iLzcT4/xzuiBO5P8dB/sVSb3pk3Nye2hxu6rYEIQrCz
V5gqdXr0zvG48KO0tU1R3g6+m/a/ZADj2mjdaadd2QbQaB0VQObxmrdGBHO1dZGDLEH/vANG0AFd
ceTnjNXzhPMIi+9KPlwLOrehp4om6PbI/XP8sX/WYtIIf9WVqUJnj+9AST+yuLMOOZ05kFfD9gCX
xbNuAezon5WUBdoo89DMHZykGVUnMi7Y3X/7U6wsb7j/qHe1xSt7RDx00X0e1t7G8SEXU4PYs4Fj
TNX6gJ6jqJWL+LsPZqtT+yq3cDqRUsJhYIFy+soLlrJvy6Rq0d5DH0I0vkxagbs9VuwBWxEBV8cg
NsCohUYFJSYPbOigXhZcssaKiqlkSmqBgLCFJbdLRdkedmt+fgCosNdhK3DdRfKYfjDq6sBbhPZ3
muuuT7Vcn1snOrMB08ICmIggc9cdnPQJGN5AhY8b7Swrjtozln2DRyvYU3Zx/XvpxrWIIwHQL3dn
Qv+yV6UgZWHub8ST7bfeUpFy3i8bNQvGjBgMddmPITR3LW2uKR1yqaWLBSXTzfP9NRYBORv+oKR0
jZX0bX6PLHY9VYha+aEK0VGGGdA7w9KM0U3Cpbn1f6pBOaxOr+1/YLtQd6FWJhHK2VTQbpDHcWDL
5pQeRvaReeWA/tc6WWcKNRXHuST7mX+9dm+1DxfSXblbKRtD+GsvuB47Q+en4cwdzS7yeUzbagwB
fmt7T58xaCpc2I7BOnlokBL+RqURV0mWcGmX9ZsiR2UHG6VIAHt96AbLH9UWOtTN5NTHkv3BPR1Q
Ub5ZtAK++sfua+pNdNXCs86orJWyUP+tHxsODrfmsUSB3zt0qJwANu9vThEI/rv2bgeilf7us5K6
aEiJYhMQx8n1BwYJpCfaMs89Hx9YxM+NWN9gjftcNJof8Hp9A8RiQDT6NG2RBRXoldcWz1JMCMZ4
hABcCLwvBMWaumT0PjMmR8cmp7hYYE5mtGV9BN/6Df+Qo3Y/SFhYkfiDfQQqrpJK4J74L4+8vR9y
mgbnX8X2AzW3IX4/ajd043gPK1JtismxmoxtAs2W1w2YDoqh1CFdzmh7Ne9sro4orPD9QeMKUc7i
rINW19uX/2RfTvuGeII4M2AHG41eyWN9EHVm8cpjfTBrrqT3ryN+Q4TNBokdCIp1Da6WoEBB7fBD
jGJO927D9GwIHq/gA1xdbCckWH8/iD+8NAq0CHoe5p4kISsrUuXhRJEthii9RxRO6FBNnRbN82hz
YJ7vN1M0G1kR9Vr8eu6FAWgDaybQhyh58rzENQiBxvK+D3ZmMRMbCf6aNmK7YVV1v9aKmizi4lPi
0AVlLWHYVl4TFn2O/A2WN83KJYfVhLeKwake8daEI72B2NUYt45ZUh5DA6QCRIJ8tbqCBHUKP7Sf
v0i+Rrww3Rwhc9IIOYjFkUF76dOQN/Y9ddJkulEjSj+QS1N9Bw7V2lreUmBcj+jH2bTx3B+zG/Uh
20csA1anxplMetqvFuYlwMqYaz+e3RGmyJbJ0K76TidIrH9HWaPsqhNLxFYaTjDj9boclAelFlIy
zSpR7rrpCvGEWhWQ+RZrnr+Br03VwVn2WVF9EgCQ1fsDcUf817Bjdvh+FvWuR3vuquVOZOLbuGtV
+J32+jhyP9RQ6WSaZ6PgY2pazBFUM5PEBTnHSi1iWWq/N08XXV3HQiPR5ljhse74sKG8wXcZJoxO
MiQAHEaUb70F4vVQ8el8KslyTt1A3nFHtooPgk+F3J/neMFAQDOfAuS9EfTSULxJM/jC/RveNLrG
Nyc2DEB5f7M83BO3AbN7MOaY5A86tm6sHmW2j99l+X/i/zcq8sIdSKQ1zN3sJCiM6BRWQivfjKXm
Zk1mktrO7neQS8M7CMTboEqk/F6ivSAUDr0wzaLC+Y7dUJ8DJix3cSbtxuFYfXdh39CCM09zyIm3
Co4VcltQrH8JmOeHqfzjoXyHvExgj1uTqYoFwAPRxdANENNZ5hPAD7bh7OpldyqLyck0VYAh3E6e
vX8v6vjlz+izr56D/ADlBoRD8p1NdVyS6/0QNB1eFFJKCVUzBWx/yzMQ7daeU4TnmnF/NH2Gfqk8
z4vbjnRrg9EZo8CPjK7luANbHU+EuAmUHQICMmiE2KHQUYb6EapBUS48c+Y+0mevh0MH/tBIQrWx
CM7BdcbhjqRLdmB1BXYuEHey6IXkdRdNJP0XVzlr3oIzzUOFNVjIL8RI2w5OOzjhhxPtzhUAtFW7
i3cRk6IBKO8o6sI7QjwcqyS4sm3RjFYj2oJLqbWZOxqHxI7T82+vfe0vmIRugRCHy1KHl5xNQIgw
gDJhxDTDq6or3cj2c2bqscIULs/nqaK5MxoJq6tyYtOFs9uFciH4+Hu1um0aSOYzqO15vHAyGicG
sn53m3J7LfWvoqtyzO8xkPqGnE1Cq9FbMQvXGgydleMOoroYjKKc0Vi3C43y1J76RC0E0gcT7Gza
nj22unD4716vmcquQ/fXWagDx6R4OzFRq3GDHdjexwrgi0BqMBRHtIa/zZxfaTGKbuIxBjkmg/d3
OpLchE3gRGznaEVTARUvuYMWD5rgYDrJWvetddIrMnq6IVTIidTKr700ic7VdGRKIa7dYPwHFoGM
KfMpnkx0gy0vIxUNkfM5cTJ7PCOgEJWPH/pIrYczLNYqTjVV4Vgk2ZrBPTjx5QaFaGWxxBqkqlKE
x//q1t+0Zk40Xz/dGXvn9GCLq39WFX7IZ8HCsLlqoJhc8+bX06EMLV0srJhIxRwGJgBu7bPBZ3yM
9Z0ljv17r9wARIaE+6m+BdDlsMXiNDBAHXe9t3sHClb66EVl6rSP9ZJBahpsscNJ95+N5vQ+5/Tx
291g4h8UcVWs78UJs7ENtxyRRU6TSpIZqmpW67TQf+ascjM4DZlIFUa489oDlHDGviq9Bt9wy0DZ
/vx4fT94C86YpwC4uaeSj5mmF1qXNFpdAr73u6u8AbihDcB0lHkUzSIDZyvZxN5oDBdEbGJFIibH
6ofzxXUH07sFe+EOHMsMgkWTDNcX5C06q63daQPvtFVwfeJxnNYueVVKmQrw4VqimUqOPovAulGD
elqTnSEHEKSUYur8L9/mR5TMoQELyD76/3uO+Hhk079ghaBPLorRUbN/3Iq730z1MZtLbEtzV7Y9
Tnte5SJFD67KZ2PuqBD0TDnBM30nqJYBFC2TAP93ubUt9ZZFT6PSU/vDfwOr5d+AjqiGnSb44Yru
mj4wavRig9fCwZLGOjjieh1leFwYk2+DERKM8NOGuG3A053dP+5Lm0o4KTbWyG4xMS3Wkf/LVyNJ
la8W630myZqARnCcjangg+TNlq5III2UWrQARnyj8uX96UxRU+OV8DeTGC96C6Nsjw+t4VlLrIbj
CRo44qQiWkJ1OnbgNQ0vSE+AROkDxHt5zg8YN1jfWr/YJtXRpBcVN18XTVIa9KZKn1ug/64lcJAJ
n4hHVxLKwGBrRDm/y7N0eH1Ny4pB0o54tEHUDjIc8NqSeKm+O/ABdARD7UzNr3mT87YdxiES7vg8
4eR5Pusm54cv+9LXAyf627FWuY0WCBOGB48ZrCpxrO/UVZnFMsH9oBWqyqKTSZ87jTxkY3QWro7T
Xa6cY4lSY+VsNUZHtG8nV333K+H2qSX+102dHOEzIAoMcI9mOOOnB9UnRZRYbU0LjJCrKeLh4RuZ
zPpIQw3fDTyKwYULTV+yrfe4Dcjv/dRjD3umXYL+eAoFJkhJzEJ7mKEzFlMbNhq6wHbsfUjPMO4P
sE8x4nQU4t+RERAxbFoHA4MPyxjYU/6FglmXFfpKYTFhC4NmOw5XltKIH0yeVGompAsf/5sCQ8mw
NJ2/YYiEHB98PSnrRDzVuRJmIfz7Vo4joAKRQJJTUkOHeryIimoNhq8TozYmlv2NDElZhs8X016g
P7cpBXl+grplsLFhIP2rfE/Jj5oNwxhcSgRfuA2Es0NENximzkU3IWTvanPyrTDO9a1cOhzmrsCY
9796Y0POhsMB7xYPSKrURl/a9g4skgKIGz8tqQhafEikmd76nrHr8tI9wQGI5auJnX9QEqdI5f8o
mamUN2FugvRMH+IlLfTTQT2c8AtUdel8rZZIerh5DNOq/T6bPeOdg+zLG3UEm0fgkuePmbnt+CuV
zsN0vOD6jAktMra2K8nFVM7rGSiWFFg1zD+CL3jjRHwo9yaAYWVUFN4h3asgTphRZSYwxiVFrLam
4sCUPdFIKUkJaVlgbi4xQDhMtF+iOgD7EJEKqN/P4qWDCa3qnoizCnSpFnm0dOtwkSuhhdCJPjw5
xjn4gfMTMy8FRoMyQ5cTwc81MqzarZ6x4178DuNpyOiaSjbjLm1Gnz/5vJmJI/ZZJWimOccyqeOg
Leq4MSN+44MSsmCMEtvAebJc/1Lxqk7vpU2Jq1fgHKJt3kOYdLTGPOqv+7PbfknzC4k1PCMzZa6+
W6UsxcRPYfY7unHyYam0WommxK5Yoi1m1obZPfM0puhZaDMsYQSpHB59rh47p3EDnjbQD5TLRTDp
Uz65XPGbLusW1XAHNYlFcOU6Ev5dVNisx5FTli2oiVo5mKd4awohFMsyDRQxrbInO+gecPKlD22y
hs3bxBAkLhpnq27DXDJnNUH+T+ZUKwOVR6BWSfTcc+SPdx3dIGvJqQmL3UEhRRGdHkl6RO2jCR71
jF+nHFG21DV8wXcnSxLG+Iyct3pPUuDBMHgoq1fYbguCuETT1Eb0auJikGGbTKcybi+bckptrzCB
cw2gPD8QCreTmQsR/9e+0kFJjWlk6jrTy+waie0Kv/gCH24PHJYs98oMg4b7MbyFqEDyyFrC3ggJ
ouDiXleOmrPFzp3W3BubOWcIbbhpA7LgaeCRIne8jY3h0MFg0LxCZAQ1At3b+ctPz6JhzzLHPQ2z
Q8HnNDIXqSu+ItbacJnrT4z+ki8frqBfjjkQUlXVjFEG+3kKMTXQQHTQkUTkI+Z5NqvnbU+hbE4Z
PFZnYiIBPezo00ZRjGvuzRYKnUAuv2Y2lwIod75WqdyqJ+xp1fKPFHQSlfgREksWack+2LTYu+Dc
9UZ8/RH6OwnPb76GbdYSw6EbEK6nJso68jsKPgw0zNlRxnPMdjvCZSK1MrbOCnGm+hLMCPJIBDGb
2hX9AMYGwgnAygNjlHvmyYdGNULF5JVZtMbN/BGzfCKbd2A+e940sMrlHsS9TVravR3gHVMPxF3k
yDqpxi1JbRJi0O7vcKc+fTlQYAhASFL2Pqivx4NgFWsijZ0eGS6Hha2FMq/gVVmConv9AUhj/t84
68bBKeyEfkowcLtMxutqpMRojWLnMItCgTYEvmN5fprjLhpcQro8IsDZraJHg3KPQ+gaIMKsVk+t
lbiZe75jTaqXy+yPQBho0y3Ulmo1Fx3iLd9oEpMXuuQjJvcOkb5VN2hiiDBKhvqbXv6wyBvx10jC
rvLDNQ1rkgBnyVuPtQIJGCIZnlgCfz2U/Zs3t/Sn8Qtfj5YKPb++chM1fSNrn1OTj3IzvuzBBJrE
aqvBWRKC569e3t7CGgkCw7Dl7M8h+YUEjeax5VRhzPI4jRe3wX1bTfKpPXUcuZSvXOgZwtDlZdBs
AZfj6yxoDFZFegjwiXCbX+uD9jm44bEBpNEf46SS7oiEG4IDIMocD+JBxQcsfR5SiM7CTfvZXgOV
Xa9thxfLLaPeRvJnfhu2KMTw4ouR8AY/DO8Sd1yyKZJyAe5vZ+CKRoFrVtNwMiHTEwqCxKxoNQtA
HTbiAWXrrrEffRyID9wAXShpoInZCmfyyqoGoIq50kukqTpz30qRXRt4TLVEyY6lu/Mdupo1rtaE
fp6MyWkQ/7bthwCxIiSOnkhtWQsxxpJNFED9gV++/UvCtUmqHNYdcPQT67CU8iPUPQgcD0S/c84f
2kRzLU3+IABOhN2GHhdDT9qwZP2cHjcwhz/lqmTPSXjBjuJ9qF2yYGIcUoG8rGyOKfGKV9fA7pd/
IosRYpQI9vH+/B2cbKUIv5Apa0b69jUbiJJyvaJSc1nEkzbxGMy6ds/1wSdaLva7vvbbRvxTHENq
PtE+TniYXERr1js4DqvVhomVb9/bqrFJZtheNyS9zcPevVqN9eXh9BL63cfahD76KYqqKHakwRBe
1PLNLrpdueQbZhih1KvNUpRjEkyWi8A81XCvYxD/3/5vm6aa56iKv9B6n8HhlhUzfkCRJhceWEix
RU1Mwr0NgPSd7gZ1U1QeZ7DapaqhXKBDWK7+aLWRuGcUcwWn8p1qI9AW3h1GEHj96dXhz/G6cr7G
rOq7OVzVunJT+zaWjPr+n4l4oxCV8YMuWhBPPghqFaAuSIthMxk6HPx4zVA2BUdzOJuZsRcTgiyv
FCh8NLWNy+kCoL0qd1alG5R1vKKEFJhJ7qcrVTuKtpGA1Npqn/HB1k83jrdAzhi4Kec/YkKiZjvc
J850Ydoy3mmMNwaTRZomV6HkVqID1jjp+iT8aUkS88MnlE2joI5EGKSlfvjzP+HsPXZG79ZkYOaN
+bStnjkNsXhkxmFV04R7DheUB/zeSrr5C6iNhXOEEeJhyW7BP98s98apONyde8YZNk/ja48EtqyG
snSISAqbDWKRi6GkPytRZpoljWxAxlBFhNvdQWass7ti+Iy/FrZem3ZrBmIlKri83OLwI8JZzBAA
C13PHVwXGs58YWPfO6dO8PLW62t7sJc0fjaJabjCbe8gsIWbfT5cGV9rV7aqx6VIGZZYyDV6N1pN
/SwoSf5gtIpw2YxFyGUTTWLr1MZJvg7ZpUpYeIyKGAWA/+sDHujb7S3OgjWSGFec4Yx9PZk7SyqJ
y2BhaL1pPlT763bklHmGJQ6OMpfapYu2sW2X/G1aB19U4/MhMuZZc5OAOuD3GlstOZ7HPLozmnTJ
7jPwN+g8ZTOZOm9LC9kxugRygfTM5HGly36nacS4ArUVioMrNdZ210QKXsHVFsSM1XNOpw2Ll1MF
BXpJ4+PxoMbJcU8QMpbEpl1LqNrh2vDCTlN6gAAkp6eb5tsGQi46H8prMY25HW+wh0I7oQkx+p2d
m6mBINmv5TShKW918tZNfCxGBQ/g8/yDt1XSQcvcs9itJPhHqs66TXoy2wNaam02QEya1b2MMTAv
OfJV4AoRnR//g3vU1bD/Tj6NtKbp3SdPidKya5+1s2x4hM5/D1cjZ0HnrhHdO0VkTXDNcbPXztfs
dAcVJQeOlZDvrkwxWj6X4HyT30BqvB7m7qGIvjNJ4vc2zqJPs7SnEAKyLNVrFSUG9vHjDOphCRWO
qLQhrIiqgs3uzH9UzTVRiLNghAM8LXXaZjV/Yfz/ISv4ZNnYPtu1YlBWfrYvimgFOfZHzsrioepG
aJ6gM5CYp5/bdUHwUWTpmcnZcJ0P20Af8rRJTf5YnebYweN3/Jr1BE9oKK9vbVdjDCVNBPcuJ8ky
NjOexIGsGG19n3GVGixCt9JO8CoKjNtJX/HyZUjPBIm/H6XDkqVw6iMm1JW8EyMVmVBuhK1hNJwB
91HI0jpFAGPC5llWBirbCck1JBw1ksLXqnMj96Sx1tvMUnJIocq3+9cs31KA9TIsm9akUB1OzMEQ
IK2bHcU0dQW46R4BKG7ilN/goP6liJBZs8Yxp+bRDtqer1T4UCgZgMU7+iTCHwTmSUyutX2EqWaE
J1LzZaag/m+26QJAzz8u5eHxCUG/ji5t1QFatE75WUXpQSdZ7hAZnppBaDl2I97x9hGaNbL715X/
eIXJ+uy1nyOJQ3G56016usLDopszqFPJIaHEaIuRuxFvyADgIy1oQsPl9EL9sw98jaNju9u/Js/2
hjW4hXWIooGKT4BYWBtxxfpt9Q6nbvWwjzP+ZOpJ0y3+4agssLPTd5cOfrfP9gLp4+N3QDgQ0otd
+wd04sAMu6zJIu4SBXHQqx6TEOwX3AkQzVKG/K74YeV4A9Fbjr69J67mXbeLyNZD2FEvs37M1sc4
Z+zW0kbzulZUgdDF5t6U4O457NqtOc7V5SEWAwSPjFFuSwubRjCU35E85zH+ZW28CNYAsDjWi7Ya
7GllrS6C1LB78sMzyt4zUumU36jcn8jox3eb2VBi5QziRgq8v9vMuzYTu6h9tS9946gaxMHh7tu0
NdCcEsUicuvjbB5SuT2NAe1yKOewnccdxVgqiBDVzZnhEiUzWUPNyeF1L3FYDgcO1a0M6KoNJ2Tt
EC6fvESCB8ZlKEiRnCcwgGkJPPqIz3vfGM7YOoeQtkG3Pk6+Be1/LWmUKgmS0ve4UMCW7M5hFZJD
WVdf+0nC67WGu/RKyGBWabv6N+Z77agg0atp035LpyZT78DpwjqxGXAOInjnHylnPVO0BWsaQeoP
womjwAtz4MR9XGMDCOqeRHV3KxIr6TDHYvMON9VAUFoIVD3ooCiaBChe2NxBCEcIQmd7+y4d5Dks
Nmuu66cO+mXWrccb84JsOdq4fI/FIiwQWaxzHt1DYy5PedXQW1bTD/Eu2Jd5bMMvluXP7EGbPaOF
XNQ1ngEIbW6sRN6SwI32oQgbsaUKY+0HLhH7ilNrOrcbnn9BTPRqFa4qUynKQSVAr4uEgXTnr26P
k7A12rsEYi7Cdn/Jg/PvlVI0+L5WiMESKbrxNwAtVLjHbzC6+3A8wir6Gjei21qJkq2VlxHyH7Es
u8ihYZWDrVE7UreLbuE9w9wzwAO5laWXwyARdZ2hz/Lyok9glKCKLgodA76mPhw1kJyvYjZu5Kxe
thCqLAwZSs2OS60VHRok45F7PIsB4ICT9HuhsL2vCj6Y4CkCC7NNPQshLIk+WM8MwiNX6iNfHfcF
LsNLcECX5fOCAS6dkAgxQnQ/CSkOXMYgV5GQxkRmfbr/3H+y19Z19raXBwoO41OsS13nXZ70maEV
KO4fFtyTVliCy9bOWPXVVHsFuC+ilIXZ8p1nz5wVEwiTwYE/2yi1ClEfc7P4eKvZNJxQo7x7rHAN
S5rtz26/8+yoScZIUiZTNTrdmLLqnRpM/cqMSn3a5quf73/oRNCAgfUn+/KN9O41RqN6a/6ogYGD
4yzOmPKBb90+RYig9LhWzBa5kd7QADJCzdwLAsCJcIOUMSK4gZdsf11+loVP2SzBOj43hszluq5p
rXohBXRWfGcBSQzJ3fERjuAcbfJPYo20RAJoLDi2BMuzxC7yL8T4YiQwfl7Rtcsj/SdZuwrzVTqD
OSU9q43ClIf79zw6vGA5d8ec2MEYSvsxzEvVzHwRUMxesun7Grol8S+5xFL94uvZwxa/lyOhZCF5
/hDq26RJ+FMyo3HszKybZwiI8i+9+uE/U5TgiVwSGrGkRSz6gPn971uKocwK+4SLm1fAjyoFjMsm
Fv24r1cJtLSdYAJX5tQD4hegCmYP1yx7FwOq59LjXWKywldSGzgioUz77yNqTJHaHE52iwMaO+hc
fqPubwmSPwYiTzI5cLvvR1kykvADkPZaPIfx48K7r4nnnIPkdhMZXRNVlK9xxCzOY0gdPXcApe/n
LCNBOrcP5Fu7lGBkVsaLLJexVDKb4Q9ngQMtd4WJE7skSMc/3Szvjg9e51y1vvtV4f4cW/Zbfn2+
4LAk6nJFXU+ecXbJGiuXY64WkiHHlpNNXwh3hmdIYYpNANmO7odM7zjjBBk4bRLkMG6SDCn0yRdg
NPbPmtSmS8Rc4rFLHWdECqtW7jiceIGTHWXQcAqwAUZaYn0AqT54M2BJZG0peviqcc9j5rwn9Qbm
0XvhKN1D6TiKNPjoM/h6JHJXKs4tsO/Q5uw7Ohj4GSCCtstk174dysjBqq2kDm0CSMWGGpDH+Mh1
7DKiljIliGlRQP3CWqadDjYLXybotmFK9/iNOI4t9uw/VrZ3InM5l7uUSef06YmnaygDJhcICzNm
DduR9+BrCoYfIue0sOvnq2yRxrjbR+l6jOW2zpqaNVmpqy/YV0rfrdWdHc19ZaMLO5PjkTxxCjrm
pm1uB+dpsjS+F1t7ECdfdH/Tpw4Z3O47s3fjDuUtqHd+SLCT8BiHkfUX8SDYkLk/MIXrFZwlL69S
cZ0ubTiIZquFUvoa/1KK2tzCTt62eT3wFmWDX2XQQksDRzLClMtcdKMs5OqOlWs6pFsNYSq8TyoX
+vtDnfVA+assELvHVnvVtFSEeYQAdbeW06nOV46GobXzOFo6xaL2nTfEnJvPh9lqj/9pxL3uTxIw
oiZy1lyEtZWI9XHEGPGnIlJNLaYGr6Ms0U9NUFOuhBoYRIIE047LBJA5S2XKZOYTk/reXUnKN3xI
IWnTwT4MeWdbweidFZ7Taope7f+ro/Ugj3TvJAB9CwoIlhDBy+k69GHPaKrb+hxqKVwPvooCMYq3
JMaIOaBbynbaLkbkf87/Vg2X3S2CuEYWLKujDVEvX3E/jUzgtugL91YVWr+HHshk0eQsLo+7+kc4
G1WWwzSHeknNlec0D9tEOBaU19BwftaXWVhKM0mvDorgQ7wExmmEi5/A11qW7ux2s7sXj02zDeou
Mv+FMHGfSwmh3PLjN3tuBUdzWxlvgF7UainCP+vyABdre+Te9iIRjSmdJXV5c4lu6dJzI2Q9gsS7
ZSQ4iftwFdbyNeW6E0vlUdiedsoE2mqr9DY20aDtrgWzSOmVPOxVo3DWHaM1TvHRNwZoT0FIYBYf
YRLWapSDNqdzHfeTKseeT+tNFBaaKepxfT/YYIm16dqi2cW7QHRpYZTw8w81LX6BFjarMvlmbPXe
25X+gjm4UFbxCqKkKMEb+L5tdPm7JsFlO42c5R2MAzQEOYrsJk8Tj0O5RxjaExzV0yymYJLQEeC7
wT5S8TctcQPH9G3pOZ42a7PQdqttt1s+fiIT0beI24q1Bg8KkekL3hC5+q/ZVTGcJ0Psv7pbKCEU
4W3buy+0FefafjPFBCWSEkFhK58hFJOoh+PhHqXjgxCbZ5HrWHfXez3pnOzKzUfwLIQpFEo+nnPI
U2lw0dVzXCuJBoB8v5RKfCs+a2wtLmT6rdyQk6ULU4mJRgDthACuu15iz8cEltsGTF/VgGW7t5fB
GujpMAcYxh/fpkyfxy+f7OuBB/hPq51rJyNGXryWgnOhUNWbCSQSczpUVYsTas1ye5+eAO0o2opW
PnwI7be4DD3aJYxxkC+YQDCcp0Dsn74WTPmDtJ9RYQM/IlSop0I91X+xT1xLNPKLu6hxFkVRjZqG
dBps+DB4qIW7J41SJkbKYru2BgEZgF8Z0LKaPt2646qLoeSdwt69spZILxp/uwsXmwM/K8Hznc/x
SRbcr72rQRxLz/fngB3yNagUGExnYZ/BhOHlgbKxHGL6pt4I1kLnQ2g560xzI3Hw3rBJ3DVyqg9/
pu30PmbBZYyqzXnC4X0YZjEcaO+/7faizLCfoRLbbZ3NOTIJumo7g9A+VFPT2hkBiVU3RMQUMmAW
DGh7EcfbDHauN3E+mAjdEKxr/FsODwW2yzaRLSYbI2hhxpSLYP9CL8vsnJQOmOvhVIuq9XEvB+wA
2URhJERQ0vLHn92UyZHcdUxpJs19B/hgyhLfYlOkHh6Iiub5D0KeZlQpdYEdmS3vTIsfQFTkw9YS
D+sBQc5JfuIMz/JkJdlRDENpWPt6a2ujWesolsRj8XYDtZJ//E9/NqjGfGb0/3HMQjbJOmvMxXu7
ZIWoIlhp0I+G7Iw+heGzBEdBWzbhZWaeDHw3oznMWMseE0mLLzLsgI1NZLXrebzLrh2jVyAyXQlu
r0KZOJkdaooCCyTrCV6P67zBTkwJIHJGLf1xAAWIskkJAIHGYf+xg5oH5/TJZgXifVJ/3FQlgOvp
yGFhyY8f4RAoK6/7bOlFWGReidqEvBW7Lu5h2TmaHlvGaxJaF5A5eXsG9jZaBB3GAb3HAxocRpMC
oVqzM+pMHbc7xA9grQP7g+j8uLWGW5fO5VdN9QZqcAQw+mLFzHCEjnvk3U5sTyq0W45VMKWSEMku
b7PZ4WXLB6TnXJ0ObYcZ07DjXpggPq+T0X4y8FqBgDq9/nHB7GGicbHClWmSJlFVBzjj0LVqH3WF
ChMr7Eh4OF/z3fhmBZqWxpkkUi6MLFpJjJPE8B6Nt2tFlnK/Painx+gxATdaOAdIv6mKyrLzKi7t
NK5dXzDWs3JSh+XxvjXFoRXKo5UnjCBr7VxcP9UogSXoUi5c1rNEh/z5un/oMybws7yiLPXI6b17
cL8tElvxMa0MkuxhYyY0XZTEdouyb0vKDwfzZazQWiRbsjYw8xzSqH2CB/66f0wWPtLkBYih5SCb
MRlEjfbz95XioavjgUCgrSPtF0z9DjZnX89eMCiEm9lLbXmWVv9LkKP370CUxV5L6rzokWABe29b
eQYa3BAz0AUUmNuerOIep29laDOFWPuwB7IgLfY+2dJaHTBeOUS+/IUTWOe9OjsjrTYPwM9VGbmd
/9k1IEMr8e0dDf7pzVuk8COPkSbpIp1ikkRifzjnC53talVgkG1uwvKuadZjkpdo2Y76xhniiysL
uOsQ2o4do/Lz8YrgioYgdHO+kgOlX884JzN7sEqt8HO6jCwqEVnwBD/6QB4Jnf/WBFiWp9aKuNfv
wxT5ssEvupyZLjVnbh3TnT6FrU80NN1InVUjncsnt5SIfc/zdNu1RUTeeP6aje7s8oaNPL3JCf0d
bFpC5U83BlNteS+FsfuwczU1dkRBtzgTROaS2ZZaOQi3TpHtZhiwWlL/iHoFR34F4ts37NV/okRJ
wcxf85k8ItI6oidY3o4J9ift8CPU6evPecKhk+xxntgCLhpMGFM9hhVSjWoOMGK13h0GhUSooLdd
kvhHPOehyIJ7/oz168dLSIQRXhpwtW4bkMHcLqY6I7BpSsNsYxjE4zRUKzr9B3DjVXNDmNVqoNCC
xYsTYmhplQxK9FdRsrTwg4XBg1sYZKvITsW+TK3sNZuVnuDmjwy+6z1OTpLDDCxyATMEfwIGMilP
IecIm0NH4q5nsjs6sl9B1YuEBFE/ohyD6yBIsh5dw4hgtaod3P6fqRR7hTFHcS2kZe2atDGUYZHg
aRSHVvAqG+hXMRWD1WhVET+Jj17fyi6Cl7gqNI3HF+Xgr+D/zbVrkNXv7oxCdlnTEp3thZ4HtqGA
wH/4rDZagRuUq0Wx+Hd9edHb5+DGn027H4d5Yo7tOCtiPU81yYWe9Il/Fic2Jy6rSHXhZQfbu2h8
NCZjltDdqMhmeVhgD8EV7mO0WfW3QZCtLB9PZXR6iO132/2u5VUnZ5IQqJG8CECez8RPV1AjZChZ
5bjHhxzMu03XuRL34U2xiIYrwDGVnOjwpkXhoGrzbCrRaHY7CbdeQyRIrvlIxNIFsPzVlDKK3O2e
xmoTEO9X00VItRl/DGyCIOXgaoVTGrChTGXNJ7xXUGm+l+z/N+SdC60UDMsW/HfRNxAqNtiGkq9J
T05fr6IaaNbLjV9GXvxpiPeEqv0QnIa4QBJvJ0Ph3BUP2shk07R1iFIcnr72SDLC/cOoqtlvqexh
NTcflSXx1Vu6D9AVAoBrKSqYGjzcoS5DK1bt7Pl5lg+YMEI4rIUxSxQiqk/OSvUmftKTK0ycI7J1
8dd/lEPbBELdz9bOmGTNc0yKCsMD3JH6YhZY0DuEk6e+7qIHV7ZJhp2sI/xRaU5h9leOVOZC9Pon
nsyS/Q/PWPy9ps2KjJTde3bbZbRwgoSME7DLJoTHar+JwCnyKTv+TreVQOmYJ56SI4n5wmWbDZ/i
oUJNx9pBbRODW/6ffRAK3VdxYNx/Fbr0FXrHOoGAF0XRmda2A9hys2CSDZd8Jk8OyeTnFnCX3W64
P/fSTfD0Ync9GRrPNunouIe+JWNKBVW1Lsf8sVC8yGS44GtkedjvfjuA41Zz56HkgF5yuoTDM/vl
Bh7TGZEJ5zrld5mGIK5VCVb0+4XbSzGHV/I7dg36WAr3erj6ehNg/qKKOJ+ltdv4t4cy40vaL2Ih
oGxdspK4j+LNroCF3POSIoZATQL5XtFmzH6SgwhYzrtO2486c3cmovmQnRoi3gULx/+jtGfvYyat
C+H8nX5N/4kvRvpYJR/hk1UfgCezoiX/ZQSzK6OHGyTPMHThoj2jBXdn34HKr33PAdVqvSY1oVpH
E+LIFabcwCNtKFDoz8E96o6YIwuX7w2NqQCP7ENhBCZmpX9O7vrgG6m6kEsmHzEGDrfKai+yZCaS
2cwllvKZvGkJSB5C2etOCMLjffYk7sUX15i4fesDdzoGvDQ0pcqdHmFOaZIk8lEY5qtYVFZv5Bvo
OVOx9S1C4O+X43g2LqJaPxa1PX3uT579DPCNiRxLqUkAkcfoVdf6SMae87kZ3otkTQT0JrTFhThN
oiP0+OdzVe/NPx7Gg6Z0P8C6Ggv+Ks9qjJZISo5dqwHsozB1P8gAZpv1BsMi13IHSvBP4hi9ydW4
llK94lsP0489xCU/aydrjXgfj1DZ27yZWpPTG37WdB2Q3bgJGP6bKMp/RWwC2S9xifoPwxiaChMB
U0aJK+X4F+me7JrMmY3Nckzqpz3dPq4/T7LZvyWbg5Gi+iWGPZeNPtPoBgAymSeuFbOlbOQJ2CH/
zMIHqiKsIWxdvFoO9w6u3BsEz7Ekd6Q9xGwk60TxpeuPjhIa33bPjB86IrWWqiZ9GtmsNeqFPcay
liAwQqYhfN5SU8pmf2PcoJFjeE38gPsCdN2XKzdF2+6yoV3TCoosuNbB1pthFhIPwcM7Cm8GcLJU
G7azr6pPBizmunKf/gSl0fpkFF2H7PnQ4EjkqhmmbYRLzqc2gSOO+jOd2hQ4QQwnc6xHXP3vk5Ui
Un+N7w58M+r59jglbBXJuyiuCRCsOyEsjRfolILkXJBxgOtYgArfuKOc5keAyLTh4Ly7uLdI7jmR
gHI9Lumko3EDlZmmpExD6zr4+H8qDmfKauWyTW3M4LD7tbOeRmKAxlKEKUjilvKdP6An4Mz2Sr4x
qggO9DmDIvemDecBxF57xe07+KX2FPGdgNRnT4zEgG9WCecgcQn+eoG7PRhjFATBPJtGTw82L78Q
MUSWX7EzQZsu5MangM9n1z3hQml+OSaqfO3Sjvw+mynn65X9UqHVi/HJ5vsQZSJTA7eVHsawpvHE
ZQu5qjMvtJO0D3EOjvm5Lj6GyCnQLiN2ycbng1PD0vB7tmqWEWByMfWVOskHLPr69aQlibTbChBB
r8RVqdlO11SF9bKNkml5rsRPXGG0X80E+RhCNPwu1fUv5tG0SAHomd1tR2i3U1Iqypr7ScKIFXKv
/A+hsK+NNHJjbyHVXgzTrd7Ma/fkPFljP9W9gGb0NEBcoAARos2imBy8+E421SivUiBxLYsVyF3y
J07yubbG+xEyRyfrag89WC138QObOMaBke0bXtJy4IkUpIwuF64gY0VmK2q80muig48cOIF7SSud
g3PNC4+xXSYfb062CrXdhXdxgtOQteHhXhjfvM05iav1CXgkMD1bDu3t9sSZlIzFrhBew4eKdoOb
EfnHFkdKLamhkARm6ghSZYcvLEVEiN9jQYCNOBT1RU1+gwWbBE5cgeToTwFoQk5E1zs8nthW150/
oN8r0z5PO2D90X9PSjV7gbUCdRhdepSR82WK6LU1ZkfOjAyi2YmhtYKCg/NDplHF+GlPxgxmLoOA
VODKRphPIVGO5+E4Fuxb6eCBkc3DkjmQjKkymwfS80N6Jbe8Pqx8t4aEZtP1vcH4sDkyx17oCeR9
ZwUwO8uWZWKd22SDRAao+E6pgYrHo6VAmXqADHQDEnvJ945l4n+ldW6W6EF8FZgE3G+jNXG1ijy0
GOZML+y9vkDyfQhOISek7Wpljg1FORAMynz1iypH3qoEVyLX2gi+Of43stBiI2jDAxU4YQFqaRYZ
bTgmlWlE+0OvWW9H0kM9GVs1kEgeXqCxVLxBvso3BL50695mPAThlMtSfIiDqz3JJVmrXab0kjwk
+2nEyfX7syTcgc+COw817hJ0UhKO4K9brbfBZdtuPSMzbaXok9o4h6Oxr/LfUJu/+iGYkQzh7u1Z
qAZRxcg9woa59GZuthspizb2JS0TnuFVfEMCBu82cIu/NhbM0ZseI2lNDMjz9xx/GpdtlggpbQoS
qu+5jwmC8OLdZm3S20wU7WHW96puli07JbGnuEsTLVgMIaWf0ZIHfTmRDRb5ivNW9GtShBdBNvLe
nQEqBQh+LnFYsBXi/BkZ8YP2H6zGQvEHYhQoz0DkWng9++CEqf3nQE/qfoeZT9qm9n9Yi5PpDkBJ
e8wYS+pHSU/Y75Ha1Zg1h6hSmjdg9HjLQOqOZ/67h1P9t3uGUjEIPPiymmhZO2oNdYNxxbwp7xx8
QXjKVKGE6nf4DhWB48kFKfvGJYlfSLgfgp9Y/SA5JnO18tRn+mKegwmZDhMFS6ZNv7MmNTaMstyI
GYtQyFI2vPQJotncDX88ojISGQ/EvJL3k8S2LVAiDNXcOCmnskbEGH6MDIxku9faFn/qzsMHBMr+
dhnjSwownxhEY/oByVuBJEDyipJus8oIKjc0X7aUyX3SWA0HTJUt4uiiSfN8Ln0RsvVFmipcPLMD
aiQVUtmooP+WvbrCf9Gld7pfdcobaer7PHNWvAnbUfWhu26dtWLGEtIA2MvBUoi48z9T4U0DglAa
NdKnuLZDxUXWlE0+FYO5Ka4mvjDWOxFnlYLnY7p1dTg1/Lwfm15lCZnEiMExehtVgpGMQs5WHAW8
Hulld1hL6zlZLRZnsxHMWlXISyci0/IXUmcrC055XLng1hC8hSJ2uKL/YIPqTv0zxUQsmHT1pOko
wrfy7xiqwocC06QKxrsUaOACyj/V+RIdnfCZXWa5OO1bYoTwfkYE3gj0FLxFsI2/Z14QaLAFkPl4
CbEbbvWIL3cOKbfUU9fKih4tEyc4bYo/NxLaoH3nUa62Rn+RYLVV+SxNitj/og5q8t0wGufSYLjS
+lhEXVuXYYhsJGQCXWPeWIWHqyu6UFs85b3fbGPEWLlHEfQuxGigzKgfx5sMGLXQ1TTfha79mwCH
FrSd9VOTMV+JX7cHrSWdjrR1s7MQEWgf7Z5shEX0w0jdJkp7RChAGFM7BPdrNR2nYgQuTeeMGq78
YPkn4V2IINk55CHU/4oqL7LBthYkvT9AblXaRZaU4/oT0Mn2ucs48brCN6JAC7c4imFmK+DATzEP
I+PaQYyBBjeAeik7gZYant49JN3AFQTrLukiBeLXL1Q7EeeWCBQSJyOck1Zhp1OXQYA098RWmzX+
eAMndtOrkrlzAc4U1Iath84wt6e44EqXb0ffrW5aKcVM3gXBSDCr7V8pYW94srjxoOvsJqKXvJ8d
tUDO6vrizGhjXaduxIgF0/74CkMPFLr3PeEJ1OXvzamvuE9JXNeLE5bEyUAfhcRKFrS39xvU9NJO
RpREbUKgSRhXgG2+ZWqQH1aTzIAxKDV+YdcSoLZxcFMacd22ec5jHsbsmhSiXuQoQVHd/91+ok5i
qNXq80VIhc9ZgHqB9onGe7wKfDxw0+MKptRquM7Kbwy5TSS9f8Tuf8bdz761Rhf9dXAnnp+MD1lN
J+dO8+2ATiQw2YUWsCrHka6xWYhPviZxVg9k/C3bDTmyLDgUL/7FBL5HIKfE7BTCe5tZHWxsGtoe
LVVrufHK3VK1FlYEB6WeOrl8l9iF6fhHITxM9CzQgYpBStP+DR+zyiEJq9oDQRLH0AnuqaPjDFUS
UTlfMgXx5QMR9iwhROUaml5mhQwJN1pJVJ0uSXZD9oOklz+SCLY9ps1KAcNiyQ+e5gmjS6ndxCbS
x683kQeQSy2cXyz0bVJucx4A4M4gjQuF8aKzLfWBEwsd03o1gY4sJF7wwmlhNXYINX8RTO5OnDH8
6DCdJ8x6mBvSCAts5adp7BHhuBZm7sM/ErvVnnPOdl8tADiDJeHRraHSFxHy+Yeu2AjkFedSdi9c
NljYgVEd7duHHkYGFQlhEhJZOhNn+F1AGWuCcjQx293kvKj6bfBiyjQK7P4/vzdm29qSmXxbTSno
+XdnnKNhH0i8gMA/rkTnibWJoAQLDZ59ye/WZufHCEMguixxAU/D66dg1vf6tdsLsI5LYOf7uWAX
iyu5aW5L1wDwyxoGRPcjhp+rTUnVpFGOVmE37O4e4+BIFkcFeTTbrsivLEyC54a5FleRzMP/t3TM
VvbHW8aGc2y1nHuVltqDyz9Cnp8Kcx4MRcNDfszoRMBz025/6/5Ls1jI6G10H0qblxCIScvJX5A4
Nnqr4yHSG0spF0tWF4S5zSduG5rhMkPaX9SkCMei6u+ojSM4qGk3dEK/EbilpQTEA4cMSmfK1kgI
ReNz2G3/ah7bqvRAON7lnB+wAnOQ2LP78nS45S+qD85alw3H1q9hF8PosamWCoJ/oDVcmHj4Cc8p
RdxIV3i/sPZrOS3k3sya4V/5KxMisMreDapnPYI4Mxdn7sqhwVMMWiqbVjvPXEqcbwV5OT0fRS4u
EN18s+6J+i+sijimV/BdQ5983bx0Psgr3ukgnDzVgnT4vSHdOp680sS3f+cnMiUgMkolMaIgiG4v
l2IUBk9AbgwSH455m6jUWyfKwCxwZL1h8Mk04lwNPuS45iazZ8tFBZ4nodEVnwYSLkMGpI8UHhYs
e8KTVAu7aKYn8ZakTa6XeV9Z0XyIJPzlhV74VWvzgg9zEx/npCP+9V3xzQvJAgQLBfFUC0neLJsu
5Sc2pUINiO7MLwUdARM7gurEFtNjXY+oal0Lv4GkK/dJLKLwDnIowtsCvE6VQ8/a13DcYMBxEqtp
qErW6FgbGzEglNYeR+4PI0sSR62EOf4TwR9rfBylV1N6tp2VjXB+q4Xw1mjkvK6AQVgoKViQe5Xs
ZUCBml6+8Roz2HIipVF4osY9s0H7A2HvoK+NhIHv7uq7noNmOhuRE575pPl6PlZWaalg53xd+om4
yEi0G1ePJFAhZzyWd6m1wkiCbrDKzdBVPuVvD3hfLhwDF/hpgcNvusZciD6Yhcxi7hhZbZka7nUF
hEO+tnuJpZWfQQAi9yBd5ZUuqHwImwFK6K9d7CIzkBJwroJ1/hrLdpPVjF3I/jQKIGL8f2GupBtx
ywskgRWHTgceoNuZTvjFzF1o9Bd6uldmF1fviKwI4ttRIdFVi1oCWEieBV+F/iRH8zJo4ljFBuVB
wzOfY+zhI6kCRp3kf51kzWWZD6WydWvT8dprbr5DNF5OdjmmF2znGyX6aBfKfk8vhn5P1F839dzW
ldQapYWAGf00DguGXE5El2MpX6VDjDYrH1YyxlK00ZYOz5E4oewGx4IvvWLKbDTGXZNZCy4DbL9W
A/CvGGgIH1Wl7Iorvkb6v0TumMNJlpT5W765cJkrPvTBLZh19k79sbAi0dID2ERD0jbaK93EfZSb
PUU2vFmwoUq4h2+zF6h+STg+SU1dTY3smxSO1vRxQlVZvE+uL8ok05Zz39ASlHN15XpIzCJHBhHL
EvmqPIYlNose4rM8tpeKPG+ZsqU8myTfqVCx743iY4So9KRSluM7GzR0sKszmp5zsljuaFvt1pIz
4un5lT1rbOYF1J0oM3W5nkzeGWwD84KkODbYPjvUakeYmo5rykAX+vUm0D2j3CnIFrC5YjxJoY/I
BU7hwQG9YpFaimzqZDDGZMkik9BWuyRuVweQ7R8Sp87FjF4U/ihilc8FZmQuJt/6wfEMdRkAHmdK
HMHzouHs/R25VzK6nSwdRvosr0E9cEJPBVSVtMaJ8rXef19sn7YC4WkAAqCPcdsYuogLONUzBfwQ
328FajVgxkiMECLzvVHUmeyM0tfRo2tdejHxAD5lQrG6v/cvWIUFGOqGeFDc8o5WJXRF4D2wcaDR
DdPZDtxfSCd9WAsN1ql/ns4s94xPpQpFYPEc8TlK2DHCxQa3hdZe46uKAbvnozMilKvMuvcrzaPs
+iKgDqjJts+Nl1jYx9zIs43o8TOy9SJ2R5u1GH43qJ9qjZYV/aiRnMo0BPjaIMLZvpCefb6UkCHI
vzF7NFq9PmogNG6ZEBXrIOvbjmeO58kPquveHfKFAAwjvPAHEox5JvC0NzscXbd/T1tByaDdiPoh
Xb2cLtroX3VvDCryzXfCAQFuFI0wR+NtsnzyGX5pb+wy3x4Zy3JBNV7/KnqzttHWTnapu2VzyhUp
qN/Swt2dkcoe3mwClIkWRnjaFB4+X1Eh0bqoRsMTjrrL1JTNc34t68CiG90nscek+AIj+nHaEs7+
/cj+oMkw4jE/ZyP9sjhUs8D2SUkn/Q5iBYIEszxH60gX1qGV6UKh+WKrY3Bt5O4cXyNknymwfeo0
U9LJueq1DmSG+82uagDSsDZxFukkBJQ72JK0bjrxrpuxNoLD6TGbghTx0wETsXuHbHz3eFBbEDUt
+amTKh7IKhMioCp/TP2Lyi0EbKHwS8PzLzNMnjGSXf1KQpR2s0pClEbq4ETYtHYcHUj37IzWCsqa
qym1gvmF1Ts9ExoazdFnE9QgkhTOjWuzmU4JEn/+XYYP7zW+h5Ccn8dO3vDCMvYcEiqe/OAd5U/l
f1gW0YZlSrl22LNWo0hvMXq1oNCA6F8DFcK2IharpO8ihyuvol03654Tt7vni/V/NaXKpH+XiKh+
/hKMp5vdbdKVBzUVKtmox88gOSwVaiyjVL8T3SBOKs+LPqid8iwH5xO37o00+1AUeexUusldImwW
kAhlArohyBiCKSsOEmGavmSNEakPyf0t1EXUG4jHwNcsj0SuBqhCTu9YmmtkPiYycUYEwyqrBdZk
VVNrSUqxEVJcbedSSq/QoBkGj6QYnSz6PmqjcR2EQlpdqBsrEMNssHHNww2ZDj8azQymXZNJTIdG
jApwsrqFiD4ov+Rw1j8CixFi9NPAJWAYrVWWvl4kG3Lc+xRXk9udXi2Qi2Jl9rMOPp5J4n1tPNW7
MqYEWUvgxbSHH4KqpaI1Obot91QYJ1RA0UyauQroJTSicbFuF0Nk8vJ6xmmSJNfHrKS162TdQ25C
veLgm0+JOlcg/9qNOTwjhiP94p2retdIQSCPWcnS6dU0zF7eda1b0wHi2NTUZzbVWUDwIjdQ2Yik
tqi9eQivbf0mx1WXxOSZPL2KcYZtW5Kepgwa+nU2mUqud/mQUa9yDqSnj7u++mDoIfoih+CPWdD0
AWg8wbGS4Nv7k5DbPIDj/XhoJzOvQglw4lWLR/ozvtXfyzGs4DNU+g/cTJFhI9YZCwus93N9wdgz
pJkS+CtkhZVQi7vb/H5R25IfSx/9c8u5KM60cRPAzlaHmqgofh0/NRFqApVYT7XProUK1mXVEC6m
HKxJxmK+1KemtwWH7iJljwCqYXztyeUIvcVTDSwfzhtfmCnca+fHzt+TRRafdzStvABhXD6DCrJA
rlSmCM4d90pAlA51daqG7NG8cHbe1BnvHwNm4csGxG4dv+1SELr4bwwah6imRza/abPburQPAuqh
q0AC0w1ofagzTuTC8gfkKcAz+Nm2UbZQovcLMT3QYlA/2o8z++l4gJcmkHy+sQfiR9Z8Lo1ONveU
BiO0OQ7dhCOh/iYCzMBVQuDkuIH5xQnritznOFh0lIfrty21RYC9hzR1emh1WrfSmmzzvFqLS8Lu
w00pcKnGfFgQWofR9/K989K8B/pLwP7pJ4L6h2D2kyxxiph2O2DJ4tWNexCHeQM+a1Ia0q1SxY/J
9M9tTw0TodEvNrYUxHs1HDty1t8WBRMdKeE69VSWw9XfNnNj7cPv6g4z2/rxdT9rx4RZa3VejEb5
5cCzX1xCZfTeEpOa7YKhjF1nmvTYRcRazAfNTctLQCVqtzsgPgLttNmJGGUyEaUHZhEdORSYLMgp
dVHd1BZ1ZBZnno/nEgBcb5L2seO1gSuQJKHuQvPx/rUQgUoH3/4X3cO/Yqk3vqHKMWA7V+QwnpT1
tbz7oXPAYovv1hoJOg1Q7BwoZKCN0+FnjE91Q9ZNf4TeSOK38NNqviSoOJmZ/mUcosMVPndNZ+u5
FxRzoN00wVfDKcgb/LK87T2PrdyZNYHW1X7chDn+MCnfF8RWWPcY5XMzavXW2/FkhhZ7Oy7xauaI
mXe89tROUY4GJK0EcOqmuPulZuETChGufLgbCITgfm8V8X/XQPVWscWRIeTZf9/dnmgTLKF5i+sd
Qkdo8luvC+4g7AmL1Gz3WRGQ32SFIDzX8s0VxNI4cOPNjEf/UNVHXm0JNzdZaYMLOCJ+wKOGf3nf
bVyuGqmAmp2h+6NOoN2AuB1vwQTSXckITVvMXMNOH3oP0/4hqH7BbZVTAJTbpSy66BIJsNjttfpJ
ahxy1x9fL4kAS9ghQ5ifXf14cxVdaOXV155gMVCMnNvgSi0lrPfV8Bs/wRciWx399Kwf4o2HCWu+
0EqmH3RncrLe9uB7Mk9z4Mw/Q5KazuEhAmvDbsFr9W/S32fVpJuzZZVzkQdPHYM78nH9uUJOx5An
w5eb2SXYswKDRDg+BwqybC7y5ylVNid90J4Gyc+zvNmaPGIbK8tL0wONfA3MyDqbbB+kFapthVHw
IaWZDDc5cV3KnT14FfI61Ae+GYld56DkJ0qVfu8vb1VyapLXhZMY6s/mOXD4UTz7bfwDOMD0WBfB
M9i+InOcH3rZxEU/BoGjS64gDrB9cjRcnGXf2kea221Fhb4jPY6U4+Vwj52QIGCrUuwfPXciXj3C
lrLbd33CBL4hHt1e3WzU9ql3CUA1BJGhW4XVk+U4YQ5uuWLTHeR1XsMX+zXQR3qr5XwNKu6RCwWe
8kxehel0ektpAfcK6Chx7nrv59e3alg6iJiITKf9cjzCrHhSwL2A8mp1HgyMVPJKlAQY3BU5o0q4
Ld2+lw348iaL9rIaeqrGqalPdCHDsoIssMLeIxSLyojIG9m3cafdf4Uyr7W2UY3IYs6EHRs+SZfg
W/NtYWI7fjolr4IMtHvv6QI8zJtkBfcID/rTiShK/aNnLXAM5jPgO7iF0htaKpduJAtcJEB6kRC+
S22GOnxzG+41Z07UfwPGuVkuWm6YLUjEUFdwRixCxuaBK6fAMmsNIW17GXBOdxVvSQnsuDhHgIOy
hKj65SpEDADSFmjFfZKVLowxol5EU3MU9i7dhHh9yVBHvhAEkzPmiM1qUPHtSecGxM6IHYx7Hp9g
HMvr3oVm6khA5HnUG7kUVMF9HCLic3QTc0EAPTWj322h6O/ByZsx+Q9Xa6z0oj6A0l+pR34YMr6W
HnjZo4njvq0YQJ+4kLm8gurNWWVhx+kU4eSs3vXivNBCzoqD6XDWLQZqHu8JN1Ar02CUtrszA0r8
RaclIsxHrxlRLpLCTXQSzse8Cv6d5i1Z6Gxt/GqI807iT3ZMwo1OZv5i0XSnit38kjMqoAN0Lo9Y
BCwfT8HHsTZOltPu738Ylw4XV38XoAQABBnFGkIzf5ZN0ZP3hP/C/EYUERwCXce6Kqhen0HyXYV+
UKEDYe+zxFfZ8Cj1CmjlhYSyR1MQzOH8jZXIMMrOeTEKxuVhY+dtKmVURt8IZBKlXVRtClspWIeV
3TYXmv1hSnzrDjxvnNSIw7TVLBPYNSrGMxe+mScz/t9imIAQLHw6e7sGYEjqsE5CQWgKVgjXi3nA
hkne+IUF0bQ9NZmXxzwJDg22l9SLG+QzEQsIE7fhwcaKF/hJHOEmkZxfQ1mskLJwNFm4WhRVXGPW
kd5BSfPLe0Bc6jv/D8c2hjPoBTs7yLq8LTn6qSEQbW7zuGSxJfIEkqxfvut3cEkhCfFGTTh0uuy3
T2BNshuWCKwJFxKu4mlbOCU/sY5lEPQGN4RUcaeyezD5L8NZ33HxYG0/0KWfZ2sNLcoVPyRh60aN
OBP5EhZGljtXC0oTW9lzoVc3ZM2iGQ2If4ADPTqjNP0NbL00g1IhPOIU83lYe4GNUTFS+cFws2Mk
W0p/lXhfBIPJNM+B62VeWuZ4HzvP7E/8ZpM0Grrnp2LNreOYqLsdesYz+K4mVVxukCzGktmLM/+s
39Yaz7sx7DBhYQlWmRRuNHJvoS01Lor5dN9DylC5yAp/wAlZbgZWWYy6qHTF7qH4VgW5EcEXzwJR
6BxiqH41CHjJLZMZy0AKTHqu7vpenWLcNt8o/mB3Z0UxiyVFkXckLxVaqUxZ2JVNdDcsiIaNilbL
ODiTYuaXycIegnzc6W29sBujDN9Iq35/ae9qOE2soP0i+nCPR2MgfcM+YzJRUMhbPzTiHf/gI/eD
IoG9EUWBuyyPlP+1xfrPaV1QyCL0SYNitkxKZR3ZEmpB8lXDqS/FTFDLqNapMiJeZDndp7bglEop
UyIkqyyYvV/ax2JebMAI79ON6FdC009yGR/oxtJFc+oJZCiZS5hhn2v5ArU7h7LHGKHGx0Ki8mvO
H7UUlg3qu4/btwvrJ617jC0IFhTyngYkvhenCh9LTrYOtii7rzHgZmonOzV0cKMi+IzILuJf5H7C
EJC7Hnn0eD5LkMcKxylRLzT8d2Of32KCTBYdw4WltYLUnQtr7QVcM9AfuF13JXA3A1j5XUTZ0Mj6
/PujTMFguzQ9Tso39jaj0osdFG3FHYSJ103Rh27mD2bSdTUO0zLrPnNbMoK8PgztbinxJH009dP5
91ghPIC+44hJeIQaffd4gzlT+/I1tMPBHiJh/ItdWYO2Caaduu7ogqKoer1CTF2CS0ZSfKcZZzjy
WTM1QW3oj2v7RZ83/7ZihEh5h1ibJoaZGNRWzzolnNoAJ0AXu7xFZHMIO0+MDuuDb44sytHSYhMy
xXitWyqJm74zaNrnSxBFib8uMeaE6dwg2ZXEq0aiFetniF3HuoTtq5A3ZnrEq/2K2JiSF2+0/Tyj
LJCRVcOgniank4eK6sctzxW51jCdVh6pjuu2ygy6uPCjiwlbsUaxxoEKhnbbO7LLF/szJy2lhAgo
YZSYYd75Z8zraw1Zsydu7D5cvV1tyefwTsdXQS0FHLWo36+MoP/gKUuYuIt31HNu2GPqO39XIuaK
+8GBJ0vGd4HM1HmL8GFZNY8G7+9RS0IPnE1FKrkv/gzsJAsEEYnFpP7Z22CWUC5XL64DyCMiOk8F
KVT+7TDRr/du3FphWcld77GBbSorMEb7ZmgM8RjYuY0N9nI7T93OA+aVomDI1pgEyt+ndPlsf5XE
5COnLljmSbbNqrI4KzeGOTYpOzAhW9GmfPBbCJCoYjdME2sSrpTs6Dl9Xto1AfxIeZ1zGrQbHfRE
XeYcMGgFQ6mnTT98LNWE9vc9Tqs7WJVyjQg9goucrZmPNEYRVnyPXjTFX7HEXLjRzGpxgLu2Eke0
ex3Spp+wUK5P4700YxJLL2Z2m4+7v5DE0MLHjT6oSCSpG/fGh+MTzNkCo9vK7DhS2Wax/JVxWyO6
oL86zZMQldyQx53X0XRUkStMiL+Ihw7OJX5K5AyFvY62GXZhNtguoZKjeHAfn7JKofv3VQGM/Ps0
zEdMgyzjVADKfVSj2K9cDX+Zug9GET7Dx5LWlsqLOjz0GrGZ6cJT8lx3F/LkrYctsGNI4wHL9LEn
Es3WLXL/ysr5KOaxOsu4ZipNtocmnmNlNq6qK6IPMnW0DxqrHT35zzHOwa+5f5eNXJM9aEk19/9h
T7eKBappaqQUQr0mMdR8GyRK7uhMZgdirt9gaWgtIofs2GrI6kxR67sdwhyiPXGvjI47S8btAzOZ
xHtuEQ2x/9ZuJjBNBJGOi8jcEAVFXkiNAT8ELyFgsj7e9qCKhZ4WdtN9lR0PBR6hDrWdk5kKoz86
jg2nJPXx/coSLkaO2ttyUT+SkIyaIMi6zruzTzcnxn1+xI1Rf2RALZgna4MAtP1Gk7ZRmSbcQtDP
5NLQv/JIDlJEacjwKGz1ALG3Ey5aIAXaLpQhev+ZkYL0gxphLGh8ZCnEpGKdU46+Y4KpgT4djj4t
zhZjqUBCSo02ulGPVAnHi2WGTUC2ntP9AW5VW2r/uGB2m1+8AeoXx3+XDsT0zYMsqYw86UYp9too
eNA1KZtOV7MO0XpGBME1N36qVQaioY2ox82wKg2tDYvCMdKsX+G/9fgLMk5qOzu7HxD59j002gBq
aQv7GSZl9EG0fuqXRKpiMpHii+V8FatTcsiY3X8r2qPggXS8TzlXz8yRhgz0pz1e58amZ3Wkk1Yt
djBNYCAWa5CZPh6efdt36cFENy5IszObEXbNOpIpp43FJV8fm4YKMcs9pVYagTsaFkG+EZw0oXfY
A/ltG9S7DIZaOhes8Advy3jsOmFOh27BYA5/Zm4YfIkFKDwWgC8Ma1F3axFzfaUSSoNg0S0QjvJ2
3EbVvwSBkk7Dk2ichMTPFuBZAgP+zaVHCPDsY5wX4IDIK6k7E4R9aUQUeLYZHPcU6MOOzsoTQvXz
aedepR69nleuDGhE4GtAZ3IPt+6rBBNDFKrzr1mFz2K+Hpyzaq9f7Q9nIog1gWAmhZu1Q+S1GLvx
XThP9dU4ERyvV250xj7vt0epnJ8i4F/+hNHpNe4fTESS//GFFqv291IPmlxuinKZCQbHJ0FI8fk8
n/rGE2Gm67bCeg+4TFK0kMjigV41ssGxDKvbDuXMXrjpvgkNGF1R7RKKV9Bz4p7bj5ZD7EBaKV4r
1QoVuZzIaUCiv1nmyRQ5DYbrcjsBb5VOEsOW7O4fgEwgIeykF+9v/V0KxKJHsL8Dpvj5tL+bxZ0g
KJ6GXX4kZitqX1e2BYw0fNgzbWi28EcDRoXkBgTqIDpluf1BigNLKvLxuubg2Ib3n9bpKOhrRG1c
D1o9atw1JCSl+cyMY3D/1GpblJeMLXKMwsbYlbvqywLk8LF9syIwI4ZemDknOVToIKEGmsyOHSPm
L3R47A4Zj1njsM8OiOzmmaS91onj41/qh9LB3gU2+yS9UYuBzDgGK9kPFciR5KN6n2t6H6c8o9ow
QasMfSaRg7A2/Vn2ZtF48XxKsggZ5Xw3NHmhDpaOkLBjOvXvLd8Z/GeF4wVMmjhQhc38vKYMMjbJ
lXq4Xi+bKccb2S7aS6noBeZtIOLQXnXHeWBgzY0CbUepe0stg8fsvgdxJWKsQGeVVa2XTcNtr9JY
xHHCpM8+YVL+ACmfrKAfPNh+B3Rvmu2u8AiQ8/M+TEQZvAg2yKG3S9UOyshNL4KXJZpY8wrD4qoO
lFQyrMuIAoU3xf2OHjzYcwjJNRoGI31KhSsc1ky08D23AJAdyM77KskQeha4eKe+vuoaCl0arlz5
9XHpa1pGws95D+rz5T3l2pL1BNeJSSk6pxkyMsOMRZaiH3rWc6aJvKUBI/ZmFvLygXaao+xEcUo6
nRwZ7NrpTAZWZlq5+xpjRQB/2kv+rJ47MWD36RS7vISK4ogsiPbuwNFBtTSSkbRJTNBXq/e3FTnp
avoMkcFrc8CWJir1kPmRf52cUgr0UkTEg7AzUmE7ebY1SEeoR0LjNt/y1o0nKAxaDkYM9NkPyxRN
JRGbQfwBBNR6qa4XL4HkXLKEQlDVSZXz+GTAi/Rz7cqgWJceZrb4E+VpCL0CeeNCR1jbaevAGF2K
Frg4T6zWKqAJDYa9cRGWphZilK4UHni0MIWPJGimbMV0NiI4Oat2SkNnLTDuzgrfq9bdM+M3JUmg
sSaTWompTQYAAeMcumDriyKW20NwDlkxoxx3LsfTM07i6rFdNvu69YkgFI+qz8A8CsMWyIalgqCB
s1psI7jVOhCcvZLbm/u1oDX+SORqsSFOEDV2Yyah4pZ+aHqk0rANFQSmEEmRRBr/PkF2bQEeLUvy
kCoSuFLZ9XaP168pjMMG+O4sGwrleL3Lp/6J70fECs5pRQJspHIULsxU6KTXfJNnh9v4ACB1YYK6
f4Ym/AkaQQcM6mc0tr3Z7qifzjoAoV+1mwrvDX1e1b7mf51M60ncNVgLpVHgRdi2w37gxu7f7ZSX
kZ9hoQGJGnZmYw4k3H5Az93m2RhoHEH3s1Z+DjhHhKKQAo4VR1zvAMSPr59Ye6wA1LUYN1GUbMUL
T4EWpxpZG0edlPVWh2TJfyJGcVJtKQGvADGH5/Wa/YedWDXkY2cx2EWlX06CGWkB+ikOlyesSUhI
v1YuVMK8lk45eIiY+v01mRZREbZo3X+X8L8g9Sy6411KpqtHJPYRcF7dd9IQtBimAW22oAc2fiZ3
l7pAhClclMphqkccQXPpKu7911jtF4u91XKnkzjSTzAMzIgoPbDoFf1RCDF9TnlUgK6bI1pCKjK4
LvbNY0Pz9IRodXcO0puIoAUJpJir6VY+C5Lj6SjPjJDDebodTJqQWaxb7Ai2SJujzCTbvksw9cOf
+9mIb7+N7udO+SUAbPx8n6L3CIhArpnqeTKJN3AeWtmXvZ9N+EMBh4L+IK7Rl38I+o0GQNy2IokL
sMaKCBSDgR4i/eG8YDOFCXIdasTAMtatUM46mhCMe62J8FvdH0JU9fJBfaqeZYFumL0f5aWFaF/g
mIwJ6ZChsTCbxaUEmjwuLvc/Eflt2yqJMdFGx5OwxGs+jxo/tGljVujkLoTCvnMmrWuhaco7MjfC
CxcKCO194l/R3qjJMmfYg216S6eF4O/8ZGytZnKx/TwYUM8XaZDAowgwzFm90f7YtCrh0bU++e1w
QRnxb9OUFab0h83Z5g5ZjjXtGg+0A200O7XXKGAPLuEZXvr58aspjdN/U1LNmOzDcd1QD1P4pYMF
KHunmYDiEvHGcFqkj//Q2Bzhnx1h2xpGLThya3cm4pMXZnR2UrJp+0IhDkS3BfKqez91kSetkmDr
wRLFSyCJEWf5JzWK0udQfk7sTB9O2ICJO7Hg/ToVEY/qsso3ZVszoL/stoYmuCI6VaWN2RAic+zS
EQZ3W0BBlT+F7qbbOcdpm2S6JomSH0PXaKbJOTZ6SgvsOw11QLkTYK3RAhQVRzdgXNSLJcciKBtz
YpWT5Ybj0bUZZ6vtaLxkoUo/Y5vyW5lL4lHIX3x7enOM5XBahMj8QM3bo7dEQFi2Uofhe9cz3724
8ccczWjXNib+tRJb6A4RCu8FcJtWcJm5k7rAvQRIaBQo1CEOumZ/nvMZo0aGM09vGsel+w4Sfqau
iv7fxBuKXRnOEKfdrBj7gVSyIR0iSJNVqX2OAvux2PZs2CbuNMv1o92UJ/8+5OD5E1MgqtycJw32
FYUlMXcBj4N7YgudyN5zyItnotE6dRvwmvLDu/XlAS+TPCfaj5SXNT6PFfhqhvXhenu+fhfezKIy
e1sKKjISut2N6I4M5zJjiaEmHddqPSEgbPg8lga5mQD2oyfQwN/l/VcK2K5VD3LB933OCuLvSKLW
pN/91M2zZC3Bbhp+jVG/BZlBDOdj6U+g0AUrR891XwpzmylVeoxlQUDWGdqia4ZuR4sCP2WcSzQR
Hk+/5vFQf2tpfs5uGYt07MEj6toQ/wFILkW7mB8wa9nC6gx9LYyL6oIbDw8+xLrjPXS1ylGzkhhk
QJzy//Y2lrVV+igRTWzgQ5wAUBDg52C7M75lA8/+mgc18NMBCsDhGSS0NeViRwIOHh0CykkfXDjS
lKzSuCTJoY6zXRoUs+mSLO9RZJ17+qNRiy+Kh+qVAVZDE0if7WTAs4eNvzkpDZ1/0sAaHL+TyUrs
BaCFwfhkXLXlLM9AkGfXjkeYczy9kyGXJKNqW2ScOk1J2Fnz4WWpiG1/py/D7fyralEkKKvCB8zn
W9FIgOqPMXNOMkXIG/VrzcWA+oFytqKRlx3oNx76vhRbAqpmCSJDrirYRfKaMJRg0PByFUOvY8XX
H+9FxVV/iFYQWqoV5IETOBE+BXoZ5UrPuTJ9muvgaCsgopX12tBmbrQzY4uUabZk2EUXc2ckersA
JfGBpNzGP/JH+lpGK9Mln4njIUM4Y+9NGIL8oVFHgeJKKD1npG58m/ccWW4jlnFesc5Zu7rkSFsX
pGKkvRpUbeVh8kUymIGJWJ8NtDYJuq2MURLObFmc8NFlrtOKh/js+7ZTu265dPa9rZbjoOyVln0c
Erfx5yksD9PEp0k5Bzt8YL/PH1tMHBTv9WiBUQQTqYVaSwLTPIdqxwQtwPNpCQpK+T/GTfRWCjjo
aWjh+g/v3rg7YCjR5kgKvRn99fTrbLJ2OX5F8L76FNQyaC0DF749zGkDLcXnhgMAQP5JbdWydfji
1WO39ATUigRFvOBWq+gPcoNNDWtlQowxLg0+F//yAE1u/0IdBKyw7lTs7fVsc/FaOcgUwr4Gm/L1
SwGOSRQTmPGlkzfu4Xd2SQXUKLntgPiU8/8TWCkkFjXU9RCbcFep8E9lN2lUrRq3/3BBUbOhQi3I
Jrsro85gbrqIca6+bRc4xX6p4w+eLYV0NW70hk+M6kr5OersTh1wtdqg8HG0XOLScQq1CoWX16HX
kL2GXWfLVYCj3V+34fwtI9cAAs5Mfp53IqujzUvXk7O5u6yxiJkKjOE3BYpEM+2u569FfsGKwGI8
kEQQIMhKWLPS1UE7NibLQi5FtwxFWkZITwaPfIdFNEDv/VUkV9UykT28SsF2eNrWEc+PH9YHkv0A
b6HzSSPWfJ2Xhl5O3SAkalx5dFE/Z0tBtfF61K27u59E1x8IjIXmufe3lraTFNGCuE7ENHCycjBm
aWDiIzlPVFcChz68q6s8gIkufnSRNST/BnCYn4EvYwZm24qANz290U7FHNWeBwTizlKvQNO71N59
BnW8jng9ZMa0Eudmc5IDPAWyhWVi5VT16pEv12TTK+nZBqNlVo7Fxc4EQ4jsDN4eieZrmtWA0zqb
6ybmOTMDnlQ2F9r4hMl5l6DYmWDJnTaU0JNVy61by4YvQVVYmdj0L1VbNwpDwfSpz7c8YcDsWhti
nMN1I4KPK/zm6tNRJ2ExvLu2bouisq1U4m7rGlRI91HPlhquXgTlfrpUsXe+ogGgCLRX1QUrXeK2
AhEjzXmPGGqXZ9JmB0kLWdlkervQdd5aAeIQjjy+O6AWYp4G6pflexvmXD5B8V20j+lIN4DSIlpg
oNza52w9fDhu4AHDh+PRhOB3TedUg01svcun5+ccW5jB3XqfoP5Hiw8sHt2qS4kKUW//IyxJ9APJ
HSLgbawCFqKJQX45TWZEJew4uPVwl2pUjGJ/tv9ZdnsU42OxXTb4f9iGxRly6KkEdzQXTkbwg44q
lvF8VQYbn4Nnj4PGcGUIVM63z19nSfcKwSdaM5MdkUOEKTLZKiv/AgvEbV9KsDktBnO/g/46XA6l
PHv+rzOlljv5KSLhsEv97x/i0mje1rB725TgQy1yGcWDKnDx3TL9pMA+NEUv9h3FnDf8pKK3hVeM
+0Bqth0kzFgrKl4iON7s7zKk5r7QOxLgaM7N8LSwo57tyyUWQ9N4oCegI8RA9furqdYTD1Bfzx1b
FeLUDwZ5iZq4dgbP9KZnwbL2B/YjRzhwqVTkamp5XvlYPoG96hdMZ3e4E0kB+M3wwCafzXuq2Ht2
buvnt13Ufp5yTF47KfoL6vGQ2kBtIdROxoca990IL7Q1ky+1t9uVcDR/j3hYE3wp2cnV8mhKOrf+
FP3ZmI8p4o8p+56WHqcxvI3ZHSh8Gl3y+papCw4cSGHfq/P9GACgrRC1XAXuiKxK2WKz7ZvYIP4t
aazgzSfLTLdtCWojC8E7fJybitgRbFTqycErI/1WIfyoiiLkA9u0Yd2F2Tqro8D8YAlTHIQspPwn
EBD5eT5EWrbJ3VlDCRMlurYigH8eNwQLIn7GLnzg9pyVqIQLwH6v0sfu95imCNpoz5P8i1d8fihw
RWtyHY4+hhnmQyA4wD8JgkcI8U1XzL8RBWywTjdmSAhJbm0gOU2aRs9jb64cBjCtOk2fEWgrKFx8
1GQXkNQ4sSJuOgw5+yocSrLK5ogAwhVrFfjRP/SqPCLdU/E07GDa9/jpL3ZLC/ARn4p/0t7tC2E2
l3DgZTOh5dMZtNltGh1Sc0QHYmedHGS+aI8ToL6gO7HyY1mjv12IJgOmmOJ3+KaaQ4eBTLf/e9Ad
KxrrMxz23Ha6vMY8CiTdf6nn5W9IgSEwamh7d91jqicD3WUv+RJvX7om21Z/jCwQjLsqydooAOe0
x406vsXqfWz+E13vGrCVSi9FqNjczcY8wt4xofylOoodSvtpEZxVMf05CK2CSNK4rlA8IS22mafz
caPnrg3YknKbmjiimo0NfOk6uHnFg3MCLzUef6ohrU+PY3QDgNIcLzTWOX75gb20CfR9zF6wYR4T
SsG8kZNx6PotPsePGP+BlGLh+heColxrg81TIy8RHPnBoKxti8eDddAFNJ03dTBTTasQ7G96Bbu6
Q5T0TswH5ZBlXdlSy/6IYkJCIDNixxkfBo668u+kgGVY5bDplz4yOvyWVkWbfzc/42Luau7mKVWT
JReOk3f3upqvP7meh5ScUnEhh/BoEimvOhGJS754MphV11CVNrgXbeuMVDa6KhBEDMQShswux3K7
XzyHnI1lRy9R4Y+s8tHiKYuIsbtY0xv6eVDGfnW+9A1mL0KQ+PUhC3/gkJhAQ4EN1p9rdSm9Cff9
ncnjPF22u2FXhSDGkLDo0Is5s2LLMEcAjaZb+it9elE6Qmrh3M3GqtK3JfXW5p2ncP+QbgA0/l6w
RQSMmmNVNY7EjsHgA/snGT4yPGzLo7cLpuC18NW7uNG3Jsf6ioye6J2xvPjjUz17BvC1wEM5/u8v
P/1rl7UzkejM6z1JOcaDG4vt+aCiDgVgs8VJS7G6/TqXvQ95ymxlQa3NPQ/eUZx6kKIGdsZrxQVJ
2KyGRxaO7XH3asHwlJj4AcmIY7R1iH7N5ZvDktbqHxCaaJd8Wpfsxdyf1XmpzVIudaW+xZQ1yapw
RIzElsoIjyFVEvbOkLO/0KGEtJfRcO+5efrWgR8sKD3Y8EuqHQtDhfnT+LZzJ2FG4n2XLAstOoVU
L75aIwbZlYpiwwxO0PpyIRh1nfuZ7XG8jGo3Tq/J2VHNfVVRFwZGIWZ83bu0d11d6UbvzImb8LmQ
kFfCgn+0bIJMY68z3TNFyX/+4xddpstafPILgbtq29QVJlwy0M8CVkLtH2snJtXZmvhlIMf2gj27
hDfF4xSg3OgEHWt9HO3U9XAj7WVrpa3jyzt8a2lrR2/mGOA0zCEeKB8jBYknSzxTRDkBa/g58FMf
gtzJtu2hmMQRDQgRFopKDekOAX8+/0xpWrA9C+buFlg1cAIRMPF3Lux6tfY//bK7M2OU+WuFnUHo
RfCkR8wL6dcvAeqFzTJn76SCyHg9CYaAg2o0dsOZ2l9pZGli6BsjRHPEGIUL5whFQehVDX2YCq4D
QttbkwBPoGA5UJHW3sUOKA6qXYLVN1TE/CxpGJrFTrhFgpCt/GKGEy/I9tA1Rb9a/67dLSboskyx
JynEu3vp13Ajv8Nk3LCbV0QIS5m4eKDwN86aK5oZHPxmjkKjRfoIvA4AToeaq9nu3iy+URyVwB8K
xwBwMGN5CK/+zDgdpq3WVv96bj+HXsRzCIRD4ktjkolVMoinUQEBgYY1zogA5kJ7KAq6RN+GX8ko
cVZWTMN9To2Dl2wYOyqjjKGCr/8A0WJzc2d6C9Pa+jMARCUbiQppfPEhKKa4fnqmAXciGHuxEPWd
V7EksnEs6ZuJKrnCwONtrU10uPiysQBjgXywLXcO/lhaBdsjobyqgKHZEu77Sb9KZni0ONpJtuY3
fT3AIwAQpkS9ya1KbrKrxSe8uDMr2jGiQOaJYiLA5c/GckfeDpxkB7LpfkY2N1zU90jvrlRyVUmy
NiNpSOrTsqSzLO2kVoPQL0NJzfFlh6wYGCkC7AFiKvRqJxIfT+8pimpMpdI/FlyvUpJqYCYVjL99
uIWn3YEmFWfHzspAT6PwzKSgUy3X8pe4XHKabJCLnCCszcudwiDf6euW3wFWK2FCvctZYIuwHTha
u7NulLIF4XcJVxezUo2PcO+abO0Tbqs7AttOILR7azxvm2Ek8d1D8s4TmY7Xhz2QLOXnr74bG6sD
NnjU3hoRO5Xst/Dwo5i+R2vkZR9brSrfUJlvjgXWsxtWBrtMxgSmdLHtCh100/QwoAYLCc5PwXOA
9MyTXli//9SUB1NS8ejm2SPBEI0ZQDtHlEaOnXGLz5B3eGHtQ6QV9oTI5t2252g3LSLnVE22DodV
aGjsTOMzmvAG9wstQ3eig98cVLLeDdaycvDtpPJDCpwydFSHTGKc8WcXjDp7e3uNIUqLZFz5eT+h
HI2YvEiMi0w/zD7axn2w6SFj/ZxCAbLSgaMCt9/D7Iiuo6dXviJlwKcA672/8mY6hUfYkh+J1Ai4
JPQa/zSJGt3UslCRESxIz5+PsjFMVA7ZNft+akswEiHbCux1KBXAf0LvgDnlewuLbm2F4jr+TcQ3
Yhhq3DjNn7lUFAImjLyGBsKd5t6+Z0g0ukpOW5ZmNl9XQgdYti6g78oov6peQL+syLlhmtq88MMC
Wy9LMpsMeWE8NNesYNhTmSmVH7rKe042BtNV/wAaxp6YtjiNIxGjV+EG5UIScMXJXtlrZ1VqCHw2
lHZ8m/QIk/ZOAXfUMetlj/932pxg3QbYzxo+kPA+kTz8ZBao7xdQ/MmBdZDHzcX2K0DqIsSmgV4R
qsz8eXQg2mRDrU6K9JUFxGzySjNxctlp9F8xtvj0g6Ysvc+j5t7dx+oNBXA0xHrkhQOkPywYPQg5
UaOz7E4WbZXbXqSG4x8kJKdhUMe7LD1kdGiv7yvDT576BRrQLpY3EBoosEvBtJzpTpN8c1XTZ1PQ
T199DfM59V5k6OFcKcKrfSsyEmNMr1lSYz1AqYnHoMyrjVSeCnhyf2dizpliI7K7y6rsllZ0FsZs
2AJ6fZeiQqZYUn7Q4w8UK+KrrgZq8+pRfH/y3mEe/L3zeU+8qirUKGiyYZEWRMv1HbexK7galUVs
jCm/8aMT35SPhJcxw/7FbRm7nyfG6Yc+G3TTnUNOHvPvwwFv2l2tRbA7Ylk7b9vUP0kFQpoVjare
+W9W/HUU7IHipm37+6408g94U2yLwgaaIiHPFWs6eZJAMqUrPOFPwbNYbqpzllpz2E4K7O9P/s47
O1hg4bjGjCm4whJaWLGHEl2G6+aibizqtkqTiVCq+5s+FT3OQxmT2MBENBX1jXqkMnjVnA01HVcq
yQEqg6gqlD2rbOtV9Mi8HYnB/C4C+k0aaO6dRGB38Ayoq9wRgxN0q0DJ05Oqh4VAcX5hsWjKP/Aj
ejFg3BNn5vyX34kxpZ8I54WcJWlaA5J4s4y3IFbRNoLDv42M6I/RdUB+Mg3AN6zoGiG2wgeWLLJZ
cRTIcuwOyt+2LDv+O7A5jaVi2rn2eZxKquon1WoSXfSID0Cgna7zmCmvQ0DDnfU4qFOyP7EV8Wmh
ugT2IkudcJFcxfunyylFuT/OTY2rS28qaisVT8N3m5GObgw6TWpw7263qOoi1vCX3F1B9q5jjJgq
xNBtkJRZ2aJ/BbS8IlC1Zy7Bm/WMns4tS7S99vwguQ6H7zE1fRiNgGv/CcSN9YTvbUSPVldPPhj0
6kTGkY4k6C+6q/2lfl8bJ8lR5VJbNoBVuugUSAJSJVdN7IjIfnrIBFOe0eblwJMq5xxhiS1HD+30
N0mpTRbVKYdASorOdPnFYDns89LnBMD6zU9Xc4Nu1bxjHwWIHYSTOTlUTsSE1QpltdU/3hQGAkEp
hmCn5jwtUG+EOk7Y1qYj4udd2qJ4h3K7QbDNUMepDZPV9R1mqP0bfQUSjNT8pm0KChQlZ+l7XuS8
w0U9Ng7KxkXGXfRNyQsQ2Y1oH8E1hG9ONu/IVmvSiLDmYYLAVyvOn+VE0PfvWG/6XYyisrwca0A5
at6tDWa7LPB7l9y9NMbxPuO1QY1BrRdmPdgBIL1KJzik4LCH0AXtzH+jnodCT0Ny/73yw0vHk41g
n2aeUljgJ+E7sz8uKXDXSzWrE9RL9V5N8HeBx9Dl4XUa9gxYUx1/Wzc7gk9XX55fjdANEqwl9OVX
tL3GzfvHR2q2OUq7NJgpOtmKIMiDg8KSUK2Sfw5VMI1Ms1/AqvjxRTNlkaf1Deo5geqLij3FBMAQ
nlOB6xFPEGFu0YLhMLyolIJlx9RQTS2tjK34hQChMRVjKBDrtqAe5gSzJqwna52NB9FxD+WX/Xqh
wWXyaF2aQ1gBBrQnQ22OhuCr0DRh+sn7NIsG+svTksmUYEooFgyRIBt2WMqhlZvvLBe/cUVJdK8U
E2vPxrc9X/7nbhlOL/IK+sdUv/zGTgyWG2m4WQTGG4UC1tJSLuNyC5VcLaQrLGBmT3lWtEOW4b3x
PoGUsOYifhPNR9UuEFYaT4cARBmW0YMtdlA8sr4kw55qloqlJv+C7wpSOfJXrrKQGoy4y1z7erwI
TyEXLQcrwMg+B3wi46AMz/3X3DFJiTVBzmA000DofzMKHx1Lr8Wo28Rr6dwn7BY60gBq3lWOE3rk
80/ZfHIfFrHLO+qsblFPBoIXa5as2VORCSsDaMCzmSbhlY2k1IKwJCQA9PT03N0S587KjZrr40g3
KY6i8ZVp+cHID/E2h8iwZmtelmunl5NUceJJeQdT3+Xb0gReWko9DR553BTZWbH/SSVb5sfx9Nvq
3XjYvvVRm2UtJcySHtZYAyNlZK/DOCDRZ3rfWFZbSlNINQ01Va9qADZh3nhHPa4RNPxuI/N09hmc
wwUMQPv11KsOeLBIuQkslkCR1OPRfwnyRiIH9KrSVkuphbgLQnsXs8wN7R/voXo1dxnLHP4EJU5F
my4pH0NIEdc4qCoB2EriDQudS8gTqV10DyFXg1DRhS9lmXkWMXmuIXCPSF3ni3mKAcHieYHf1g5Z
EUCnlCS1ryjA2Lcs9PyQkUn+0GnS7US6abTnr4FHI/Vuu936ejlXTeNczLR7Ekoc2L9Q2PEG2Th2
tQSvUPyZ/Uo151okYSMxx6FBxIP40GkMH6O4OKsIc3ci/21ASc7kYnVWvPgIxaS+fIWWbQtMk+KJ
uJSW38Eyn6CSwc4Ti4o2STcqyib6egmnDe2SFe6oIvBS8fqnGYcZf2PzHUCeqzVAILRafsVE0zsG
F1lEWf3J1vPT2c8OanLQ+Wqv3NpQHYnM/I+ry2L1t1fHMiZC6bB4JgL+iY1SZgT8hKpGXo1jT3F3
E+FIeDMw/IJAUjzUQqM9hoAkYeFSVA1MX8INqNlfPogzsuG1MU7fWQCeGNd2AZUal/DEw1jYyMs0
JOa80c5yUFmmISvAw5qWPZoaZi9I42gCEXgi+5V8J8rbBtJEmvVkcFwJltTGK6sQ0RzOfUA21FDp
bI2z+LRpSITmDA9R8SP6FZ2aPBhefaIIFIRiFB+YYysw7Hx7EvAOU/NprNxZ1fuOfrrKI9t8zIo3
waePaQ03LPSRtQLRdnirGl42plhfGGOKeaVUKY9YQNs7pcGb/GxBE+PrDRL8VMZodaX2qp0qfn3M
7VyhjnJU0aSgfNd8+TqGlrC4kORKngQc6LiJi+0iOBO4Boxhp2HdlinmxXcs+tnZE4j6vCpshVVh
io8ma8El3MA9mIDDOadjW6sCbSM/IEbzFBFdsdbmkIP9q41DG0xoynwltHjFrAzp8PsTbKpvzhw7
jvwwhCm4wkDI+AqWkGNzVvIeYF7kd+RUK1WphmSaphORynSpBi4RnandtIhAJZToOM5V+GzEpb9O
la0kOHxo841Ml+xLlEEyUjDZZvucSzr3KJE2q+MZ2AC7xM223Q13RvkEY5T/ixX0RFHTN354cuBa
i2vsIri3G8gOiJiqW1ZM/JGF4EBSpoRJ2QLTzO9VafMO7ym4zd7wfxGiSu7I0iIDAw+o4Ea5oNJm
NMNRdnTtALxmBekWGgu/6nIPY5vT/7WdnhS2f0QWyilppwP1/isqGu+6rRYszjrvBBETeTq9K2uL
uIUwDAuFN1vyW+YQmvGjuPq1vcXSxb9iJsF/zlm9ZacJG0amDptRMJ5vdvWp5HfF0F/ghqShX5eG
NeG5MciK6GsEpcOjpYDdHJYIak+axC32Xwo0zCkqDU/ZrMYQvrKTGqpuP8o/QxoaYg5FnvSGTTwK
6HGdyIxjcQQNT2bSgt3eak02yYT0kU+7022D3jFh8jmQ9ytf+DcBx1u0xDbT8F3VUvOCDaGn6ZBw
KDzQ+zHyWSjMWEonATqci27tCM63W7+6Wf4olUKQY4AZBDWEUWlEZ4vtqY7smtKa+urIM00BfAiJ
jaoyjy55k0FHvAywkToiZUSMlYHzIzZQvV/+gmce3mfHrc6kIKZSsyOuObSTNkxqwtaD3lOlEev4
B2qOq0ovvi74zj+UvUDmnUBtxGnuonUf6kLmBbZ52N3KrWDQ+5UmOBhInZAEp999Pk5GfGe1+Dod
T5ExLQorztNZgGr9BOCq9h6Obw1np6ZuBjD7tK+OnUh+Xu+YRtWuhcS9mRolcMQpyclfejLbZ9fg
ZVYUZkSnIxTn+rC+6pIrQMBsQxvNEmo73oOQ57cvzFo6wpr6q8tmoyAWDbkboJ6v6TR51eeOykXg
VKqis4EwHUbZBU39tFLdaKMr6nd6kwXq8HwwoTouxXRleWPGpeAfZce7QvzRciAwlCTA5nIf9iDg
/yurZ52kKRFqRzLcuJhSQAGdg8Im/yacj2TYFkKpPsz0KfPtZIlQlHzUxHVwU+5AOjWUsP00yHAl
2Lo2x2BHjVSWHUssuhSgyo0i9hUJuvtr3Zi0WocZzXAJ3ifZq229f+V9jqohkp74QIe4MG04DVUw
v3AFQg2y+2TIAZKMyls9SOXyJY0+BE3yo9dJuLcrQCzqq9XD4h7B/BUzVqP3Qb6LR87H4QGs37g+
l7vf588TZuxXXYgYOUPeFbeAPXwXA/5bqKA3lOTRvL/vPAR6l/FFg0SXeiT54qCd0HnKZGFFtkr0
PeMvPCgfGGzEATr3WkHocfZKWaYRCHa0NyXkZeCRkkAefAa+3f35yNtQ6RKzSBf3OgkrwoQYqOjZ
28xG7i12wZuxaDA0s67SI8s7q8+iCpFXfpOXKkq2AzkWioWAWxC8fhqFDPi4i4ZC7PioUAiIutBI
Nxb81UMJcsYciCciTz2qhHD0helt06uC7zkJnkwaAoTb7CDjzyuzQ1LiG50HukhK/GjetRJC16Sr
5mTAEqZ0n10HWGGDizkKA5ylhjaZNXnkmz2Dcf537+z+w50YsKxArbLiN+OtsCYzOAF5cSAdlczA
LqQHB7mJllEE7tNsxmr//sxPGbodmjCowBodOZApQ8Cgolwk3TtzJVuSBqcPB50DF21E5nImObfX
vqFrUg9NyNIxawqTXAIkWHWvg61WZLGSSxMPj+Jd1RL24Myy3Sh/m5BMp64RAHq81w6omBtXvgyR
oG9Gt5hvkWwnZlpyxKNk1jIe62t9MIAEeTCl5jT5SDV3i8X/MoUzPoESoKuBNlQOFz3PLyN7W2FS
+omG1QR8hnFeuL48Iz5vabodyO520BOGW8QDqPgENHGcAEiP9vmmQEkoDhaxdBAr9U1Gjn75xJ/A
BfTl2L0pNwzeOqmnIUMTU9CGl2g6rjKy4LQHrYDLGUgJ0IBX3LYo3jSmu9FGKHBdzkSQv/bx/2gU
IQZixsl6eCTYp5LbmUrlMNYEnnz7xXyxpTuXysNwlbt5q2X5p8pyBrvSIH2fBzv+iPbAm3/EUDVJ
5+qQcBzByCaoiXmkUNwvxclWqJlqiT8pRhcN20RnNlTNA4CbW+wIcbM0S1VhlnqAlatIhzTNpoPd
vUauAGi1KaKdZ+qmwh/Xd7z0MXig56I/ecW+QRtov8rNLBHXyKIElS4SX0O2eYKk0qFs3xwzbDwN
jR+JziDxp71B1j+3vfnT5hteBCreNViulkal+erxqLzGyy7MMQ5pjoYx+R73Nt5cpoUo8o74RjZC
X+9Zier+mut1QKI6rkWiOWmwgN/iAl2+omQyHpIvzkUBZgC6TEoI9V3oadwOrn4pGsNrILjbc2dZ
m3ViYIew8KZ7z281Dbzt/FwRYGf5pcD09xpeprT0n9fGqLvOQqTLdKNEl+k7NGxQZdYVcr22r9nN
Zb7yEfsURb6lcTAZVznNxF6u+LKuuP+S50ENgf6xy4zq7yZSoaxI8kXPbBz4dQiKR7eATs8uESMw
8SLJJ2UpstNItzJ90GrsR8mXrfVfLj6P/gFuusiQdcDrxsbgSeqfMaurYCycFX9SjKaZeKQCazTW
ZcTOzWUnfnVexA/bCS5gVBnwzYKuCItagwmoSHxIzZVgHqQSFttcXzvv3SevRe8c3i8DViuijeM8
8JRnpgdC6wztEEv3CtDXZjLMtxrF+/LQq1xtl1jpdPqrjbm84Syi1jquYtPryErSaJo/3Ddb0K20
fCnHl0+Kwrjhrs4bZTeLFLe/3dHmsQIPi0e7zu7Fy6rh9o+fo/8HaftubDGtAop0bYoNQbXWtWI7
HHsAQ/27rS05aK3xIox400qZ7W4SAiA5wgr9vZFZRJnA7Z/rL82lUNToqIEHO61ZrHoABtJiCAa7
Ampom0O0/L8362/HetsJGv5sIbtVweCwBr3onkGU9wKC6mUWrzPL3duCKtJuj4+mCLGhQU7+xcRD
FvQQDhMuqR4BSLUftbOTLX5zLr76j6FDoWH77lvaGAYfjUNe4Vh16ESgK3gUwa58VhW0v5KiSMJd
t9GiLI68H3nZNsg3wjzBwSggxFYCl72bjCblOjNDZaxYOA1CEF+LoLsKKKjk2+19GsjEzcGrGaFI
pKS8kmu2g6jb44Jk3a/3Q1M4xNYehqhkc9I6ZV5ByZyrRTBMTN3rBY0vmJmgjuJX2he2LTPn6E6O
lAuI3dFOF8vRwt2agGDi57+fv2Vpv9FFYZ13ig4OalXDMhA2msevlPF2E8eqJDf2SGW/FKwlCWdu
PTBPVKrdg4SIoJSsHfuewylhipvuXDLUTZpgrVwgbzvsWRh/rhu1ooUH+/OeTUdMGid6celRPUOV
E/QvSMa4LrleTsyr7OWxh+O2NL2SmB6cJz0+CnG7balq12awGKK0SiY/kvN1O+NTi9TJc0Bzt3wF
PoVnj3WWMhbW0olhE+eiEYIWF3UYIBPr1svhx77E16m2MXXLwBrRR+OAUiBjiAUkJau0dhXKAovL
Q0800C6PDpzrHZ1Eej37sjazJW+bLymYKbvCJUfecUwBCajBHVJWkoJ/oiie8jPxOpplv11G6fWI
NPUsdxrjm9WPxdMJusnhWmENxcWcbY5NQoRnB8FCmXYhbKtszTPPmQ2/+wFQX9vQ5Y/ODfqHObYM
4CwX37QKGsYGydXAMSlElBQj4elayqmVMYQYybtFprNabY8vRZJC7Sgmd+ALPWezxTmM3GHC2/6S
NauED0JWcHsaSTxf63v6ol5K7IsCzyOCrIhOFmezhNG4//96wNO8/cafV7KogM32gvOZk+XAjQaY
5TlHaRGZnLNEf/2WvznTJbVNnGaJeB2UzhH1dRGn6k3iApMz/i/toNO1H49H630bt1cDeZDQcPdS
r8yB3HzHdDXFb32mOVsvZ4mKHSXNeaDBKy+m03dLA036bUtX19qZqSMQYeYhfTV7A3ibgwRFldRl
bUBnVNJD+/d0xPV1Pn72veG65iSCxhYTcY7e6PkyBcKt9KqVy9yKbupA2CnIimGwVCvKtO8LyIAv
j1MCXDJdzfUehLAR2H25+EvvNzUM8z0JNhIB3WiSZ7Q/+b9c3cZvROgkitrrBLohEmDU3AuPoGvN
UilrUgpZHF4KjlY45hI/X7GxVoXiMemTUII6qdyBbh92AN2EgBP72friC2wAooOvSlr+S94CtQKn
FNZSDUM0EiFQFvXU0emi5HJ7VMroP3/R7OIvfMyG8ak8WIXF6glvjI1O9h6XpCTNRJLWGkkALBnE
LBUprad6fNn8C+Hb2gFtNFT71BV5XZOsTLCRqhhsnWfpc2jonS3aikdR1HA3KcvUysU39BIoFkPi
4fZak8x5gLuy2jqcMHZd7T2rPROXB184rPXC3yCb5jk/o4Bxv3j2+PrYJjZ9gIGwF71IPN81u8TU
L0LC5zyNUkjKCyvOeA5Bs3t+XXq+zUbUJkGs6D7MF2bKCbIYr2fPtnxc/+LYnW1ddq316d5977+r
FjHebQqONeY4l4T7fcx9RXUi7JTuY+EdM14vINqmYDHimDPQx2j6QpkaAr71B7Obma3ClKgYPd4T
RJcnJqofjNh0lnnfHOv/culIZWX99tDSYlTqbFCDewK3K2p6cIcKWdoXg9MnjkJNpfUZHHlQybiQ
J6FkbQu8f1uNXVy+7fxSebCtmpmldSV8+2yvW0K0Mcg1AlOseODykdzrArJkzqi2O867NEK4vsBG
6d6zd510F8rLTLBAZ1tLqAaLC9RC06NLK1E3+nOerdMAzmaheIewz5HHmuuupapP74sJvCQeg21J
kj4xFmV7ha0mVC9eINMF3OfOyif+NuYDicgF2zSZWELrfL6uAfn+otE+yVhEeobAgDAUVW5oVYYZ
huLKJewrVPehuH+C6dbP+ep/vI3dINuXC3TLx8kQlYdAXXudpMG54OusKxm0Int+m8EBya2BFQVO
VPtVu8OSfIuXADb2qPs6ShCvksnfYbuSJea7m3d7w+42w+Z9OOa7P6ZkPMz8A/VVR8nwpdzhZF0K
RWXtE9bPMDbIzig15T5xM2aGLINz3PYZxEUyGkw7Wh82nK1snODgGFxrdOHi+3QR/ULs9bmReCCH
al4Jn2f39eMHdMYt8EPakkyO9FfreA1CA6uw46NV47ZsDtqbfoj5OWYrvX1vRvUzrIS8o/htyhsC
bU3Fuxvwb2W6HPcHCDxbAhcm6318shfQgmPv0B8g9mFeNqowhB3S/WzaQrfkm1PJwvSW0CpjXaXN
JZQnCY0ePpVrnI/tUzQn6C85MNtVgaWQdD/kpp3ZPOpEjQSC+xbTPEnDkfzGg/CMOhdApQv7nZqb
GqCMDicPvJaTeyRI2X0jrcupJnltYR1mT84yWsJCcn3PAd+FBGd1cNnmUmG56q63WDgJ/ATlY6a2
XfsQDZo8F3BiEI7FBtj+ILUxSWKzrzNl8iMPiDUx9mPqvsEfPhS6XEVQZx5LMhsGEy/PGIvN9q+y
5JVF3Q77lZitf5MknEKwWJ0t5rymMIhI/f9AmTBOvY0XOfCTXIbFdePzkETepuMVpMFTwixZj9bd
rdWobzu7PwWebpggZ3zsoIsoaVSE7oWnPXrDG7SWc56RR+eNV3uxoTivViIYrl8HqC0hr8FWgoFe
12Y7UBHVtMxIzL6plOp7G8iTk0KrkXF78fLc1399xMechVm4GT1t0orO6qscVbivLnGSoLZvElPW
EoknkWIZ2IErw7Jedp4vPzh7B04SP1zOrPGOq8nxZgvgVHXsYkWrreJIVH2UAA+YNWTOGvrFiwHX
vHHtFlrmafAHLB2hKXX92IzshSdtKEaOr2oCUgAx4EcSCtzhRVGzYsOrhjGPG0bRzS51SkAcw/gT
Jd0VW4HZJo5NVtjleip0CLphK7QLiaqhrgSGNnYeSNnYSVyX077fprrENRRoByN60sxwkgF5I1y4
suLg66oaS7n1gNkDey37wl4Luvb2XzblFEvhd9a0t9EL/lzuYdX6VmuJ+KIZ78yamrc2nFAY+Sst
eMd7YlWvM1vYVRz0/T+gnnGkFc2+391MHWVwowBsTOTRJu47nq9Neo6olDpvS9uXYAvbJ9Hm/Jsw
MfR0PvuCXrhrTWVorgPgT8iVo+fLTF0zhsp75LU0cGf0lfkXB1IwzOefa4/WMOR48wOa0xg6NejS
99dx7yWavLSjY+dp14bRqH0jHE+jB1Oc6ExbsHkM/NyY9eZbKDK84UrH1D9cc7Ne+rcWz5cbLv2e
Ule1fdlkKTr9/io7iPZigbqskjyLI94Zkk6P+RaPmNMlDnqWd2VTrSbqt6wM+KVEbDULVzEGplT5
vlsHSWz6QK0KtFdhwC2rVdin6q5gpZDE8EdXOG2sVZT+zHhDC+w4Jszg342R4U7uamGuraa4f+yB
YBqCZEvOIowEvPDfgmZnL45Vwnywj780gDgAD18RUf1pQtZnpxkK6mSERC/Snz5TEVqN6X4dRvhU
Ro6wEx6A296gD0+qvx/6Cr8zitUUXe+a5ESquMDJJy9qvgLSgA3Bd7KNcLVt57hV2Gocqh4YPeFw
Zq6qgcJw0nvtMs5DPQhhy4wn1O7N0KoCGidRHj7/kLTYt96tOh4r+gRw+GEHGCaQr9+vQYjNoLiY
1GNb/mCpWVKEMgRnOrXAsbWeam0UK6/i2WQ8uWT9JoKaytYue/vIKTUi7xYVz6J/hf3tz+ZfgIeI
OJIkEBZXxUWjmXNAvFWHriox0u4DgsJIfnA+4bTkNfuzsRKosbWJ57eP4i9H66p6duGzYKk15q6L
u4L6zJOoIxHp2e7AX60nmDoaGVeC0VOCzv6FYPpmNsz5M1BevFjk8Admnj9dAfXTzCao9V+a4of3
x44g8pe4LykcxMzxRZDBgIjGKrs1g03ffKhuV2hde17y0IjEM5WKumPdlfw6GYS3Oou9ZyKQ6Mom
SMV3JYcZ9PRzIfomy2TJtusrO+DswovKtv5fd7HcKZElbtIV3J0Y8yYRgKiv2XwAomys/+xBYvA0
7Shl5G/kD8SRA3Yklez67VVb6f8SBKxvZIHQjHG19mQTIauV+D9I2wE+CBhSsIruR2WoNEQiUWBD
BAQGvZs1cszlJ9PnuHyCdQdtcUVBl/5v9DWcVdgsHByJ9fySxSspaV8FacrBmb5Ix8DTmyWDTpOJ
8Ki9Xsy5FJtlZ4Ey7AnbZR0jWR/4JT9GqwFA59nLzUbjHt2sEQ6pGYPkYWuZ2v/6yd8E9TKYLsU3
4FVNNslfUEVJ/YO/YvyCg85o7r5b0BBULx00tU4qkf2/1YhtGoeCJcxM77HOnY9XPkzbVdsYGPrK
yisNClkkKiRK1GY7eWUEwqE/33ooA1Y+jIHHmE4rt64q6+v6V0ghyM/40TNIuJdFrXD+wrHAz7MP
CPlGDCkcWtFD9Q7h9VQ8WyTOwQQqDzZ6DIdebwyaTbznc66O3TItY92sYFW5aqcILwDyUDexVk50
8N2vIs45ciXo3cc7GwQwhOqZvqi99StCSOOhNmvLG2r7L1UMAD4kH4rKINwlRD8RGnuINpbjdiHj
qzJCNclCVOHEf42t5BIpXuhxAu/oys5w91hl5RYhhXz50WVTxE0q4OoArcJkQN3geUpY6YzPMnEl
3eVi6zC3L7q7MFuRgWeZ5wqERenaKJrLhm/DHzKw1HNdwJvkf/8huaQoaC55P7aXG/LRrz3LbZVS
qAOjf4/eB9d54buyywQkx9MzR0TgbbSSHf5oRzUmtB1c0KrFyhmSHsEP5MetZ+imNolLLF2GxhlX
r96Iw3smh4Z1+ma/GwEcAWIytE90Pe9HvOtGunazqg9Oo6+DgBi1avy3GUihbmHSPrPrkn4CUlWq
MmG6tNHQSlJGjmXpi6GIrywsbdGKDr5kStE9uwCCbYM1fX6Ta2HEY1DXmAVhkLaluZvHNHSorJMk
Y/i5s0VyMhN8xR2oeYQ6m/O1dX6a5ytGC3bsrU3hcom9wSQnkP1C902mhOpz40Oi8E+F17tD+VAl
blBITDnH6ktT/+biMxRAM95cNFgiGDqdIcC49hRNSEKY5MjunwhGauzPRPcJFlDmVgKHTx0IMNeM
4PXUtiHs+FlFN6aLwARcdv5e+5gap05g2lkA+ysKte05/3fHdYvqrUER3ocysldtH4GVUorGF4dx
+i7pjhFtZpBRAFTjhqpmZ4Z/D41IcFx9AfEA5OIAJvmIRCck9QAzVMKU/iPmnA8a2yWrpnVgxdrp
lg47/Xo27LHCc3RFkCwTKBW+y6f9IK29mkPdXC1Y1lfl0/xDFZv6opITC5ALxL0HXSAWZ6rwPplY
jUK3v7nrngATNKV353ws92AbF+or1xCIybKZAT9mztNUiqQso8eNb0Lp3kfZimo9Cd17sby+W4U+
19JIog5VHs7uuhYbIznO+j+9EAhUpX1aZ4DyAonYydPlZID54yZLV5RgPfCTPP2kaIJuOWrcAh30
5YfrXP+cWf4yfdnMn9nz4wZqpUj46zxnt1Q7y6dl4Ij9eK2Er4wbjY/15uevmnNdSxeiwhb6WS4+
TVWcovJuUz6y48kgTT9Fc6+CXLmtLM6n4JjrmRyjKaviWbU4GQIWxqir5g5aVpAU0+hpAktcFbvG
UXjFzAl7CMuL9xJ/JpakVVy2yYu99nn7ND3B3HRX5IdVaboZlB47lQRpzDKKwerNcYhyY1egRpV4
zNveZyfm7yykn++02UM0Xffu9Y+Wc821T5eEwp24r1IAO5Nxn5xjYkOdhzViBejA+UyRQ1M0CJTP
wPkI4mJavznea+CzWMbQuEhaFcs4o/wNsAdqrROHiU6BkpMbwM96Pww1Qv/ZfpeG6dUQMPwBUtLO
H1VpuaE8nhgYXDeuHLuGxsjFCrbJo9+V57cuN58DTGhqxq5lEep9m8+sjcMZKIHVyWSY9oMNi7ku
qMFri3ik+auhTy4+ZjiQBFqoKT1eiciNeM3/p7Ga8eX9UzSD8A8LreHgOJF5bdzb2krEpmjw5nO6
P+Y2RVODP3VBq/2I5AI2tHkp+z/4uEEQSYtaHNJ1M7+nbOiu+9I7Xqve3rg27TsV4AopYzwye6XX
/1ISL+U7IDkIPttwuQ54SW+blogtfznt9f8rXkrQ6Mu02hOPdgZzbpWASbKuHfPRyhXD77GLOB75
3uWjPbGLDCJovJG51DTl+FIZIYZXQZpI5Vm0ABFekIj0JESjnuuPj5Q/8x15qa6ZEjAxQ04yvB7s
hXglYEaXoScCtP4mTfZG7EvL9Y8HwmHiwTFbD/JpIzQZFLHvgA4cjFb6xTeRSBjxfaAEQCdx4/Y1
R99B3uY4eXnecgWhiuTKkKWBSoV21tpHe9lTBtUtV69fo2skMaNOqDdNGfd/Dey9ZzpmwX467X+M
Vm19trA9LiyydnmAEXJeMziEqinXaWx++7KoKuKDoi1tdAJYJYRwIzlL2+FuSDiqJzzjwVnICBZN
r4ELGfLYZIiO9Q9TUDGSDhCTklpnwVCtTkElpH2HeI8rLWOoHBSVhEv0S0wXIS/hqSIwmpIRbs6T
L6dOWnkdNIspVBncUfIUzw2njk5itmCBDL6AQLTNGCSSlgMSI+ne4GDpS//Fvvf0DqwoeL7ysaPM
zzpCcADy1D+dvVuq5mJmTJhPI27u/oO+WeNaicuO/k0K5qBxyNFzfNzSpVHbIqVN4Um8XVRr/Tba
QymtaO/ns1pU+JDMnsyF+YG0LtklRQRaTtrewSHAUNiasdMvFwkRKaqgd+lqjuLKg8TYGkTZrrGQ
UDy/1UkEGa+tgG+RRIqOIOo8EpvnBJTXGUC3Q+FDUw25cN//YAhYD961elk0Xlm7i63FSMAoXFVv
VhRuk6JfTL5P08ua4XnrMFG3WHeGA2DjUr0do1qnv/JVw+o0hB3b/QBLrgJ5v0UrOv3bOngfP3E0
iNrislkT1DziaCPGvI5iZ5oTU7czcSw31nJ1HTKAEzcgcn7uaMvua7NSbiHnxoh9iUc3jWbo9p0h
KSmOi74ABSidYPPOg8b/QStEgvRfQCvu6+rkRfA9LDeM6Sqe7wYIw+xMmAmtPP8ZJtrd/NG4nyix
ZceNu8VW13+IwEqhWMBcF7ocxL7d5KcMFQ7UH6Zq3hgpyF0+H8mGVTzM9y6RhhoqAtYlIqPvBdPm
AZIhOD3e5rbug6ryo1gFMTH4ABC3LNqGHU6na3hyTCWG5qRAG4IHS+x6pkWeyMU5mTOvnGvUB1A6
jE/ORULRJ0NjSiKJA4y/c2FOSYP8NsQLp9sjg7Rjblwjg10AYPQYNhj3j83CGfybXHIwi9RK7/UF
p4wGRGc+GjAP+Wcf15GCgjX/47h1tJzBfTUKAwd+S4DQelQSxkuQwKf6hqY+LKPVwnWJ8hwbtf82
peBiEefRBzl1isaVcZHadnBj6QMvaxrC7uFPPjwEkvuoJmgu1KZYwic/g+CusjYsCtglrvcZRiHI
VzYAgWA/MPe6YY/5ze6NW/9gr0RIS000V2SCBs0DrfRQLadQAHc5Ley68mO054XlW42DNBMC2fK5
C8j0tZFg9zj10w2XfWt2eibr3RQPxYa2OYeibHWb3nOKprnDsD+7NmC9jTwfaG9nA7CPFtee8M5Z
M6XeP6eywucywKOjS7/4mN+k09MQjXqwxZltFZl4bYoZk7PwKZhUR6dnlfC5xdoxmFYS1H20arKO
o/CLRJoH/w8y8hHnRQy64ROeSsNBhbRcDsW9ZVqHYqYmo/JUdgUTcQzFcPsRFmI7z9+du5iHpIAK
dEuwMndg5HpNqGy+v4hofCu2ShxnqWG8+yZgGBFa2rG3iRgQK8678QiLwISPqof1sQ0cUnlD/cpv
R2cz55DA9D280KZAT1ZNMV2S3EUmk7hlGI7BTqcuibzUelR4RxRUiaI55jL7DPzyoBsPJ63QCtuO
ZHk0Tj9HIDaQF++fxfxD1yBPqaldCwOhQty5vmFDXdIaoDuqyls0iepo/IT4UDatCAvVvmrZ5y4H
of9tIYh9AWNbIkUbp3M2CCJjqget2VVPlDqRgs3RUHzez0QvsHfjyR0c1ubsdIz1pfXthOqOezAb
4/K4FAI1+8TM1CIjulk38qzBS/nRjBa408Acb1XNKGIQbu44bpxZx9YC2b16/Pk6hTgWEkk/oIg/
g2t4sDG3vdlpqNK66cRQM1jFpSyVgVC0so6hrvHkgzwc2GNYqJoVfmjWKCBmFxunld2CUltzacIr
3pKK+gSHT48XejkXgUjmYRKVhLA4/2bb8hiETDTBl0BOk0sceYZdF4pl1GH+QQRIEeQwHVEpYiFo
WPyq5xomBS/cCza0wbGaKqx7QCybpgubEvG/rIfyGhOttrL78kE7j2mk1DluQJUILDN/9+HBnBeK
KGSiG4n6ipYJy01jn3J4LeedO/RiNGZAOjIbbKW4AsAtZdxM0xY5g3zG/PUALk1mk9Y49m9xOKqA
lymkPOT5kSF2bY11PtH4QMGfZkP/t8lMhXeQ0mP/XcAbUOI45UUd57B6Ro4GXOAHvQnvdprglNOR
jwrq4ZoCNj9dkCL7rkxm14G8ulnMtShk0QbD/rMWrQr1fJIWX5RqhOJx9Bz14rKfDBPlw9hL/CMg
3bqNS/CYspGQAV7eFMXq9I//lmntPAMre7xWWIbRImsxqwwUKKWkVR2uGjzxMhdrZyvfGZhM6VCP
EFtG77aQdBmlhzFGgQNmd/4LOysXfpWtsjrtH9ZQlvBrm1+rYLh2ZYfvf8bLcurYADCZeBEkhBEq
Pe18YvGbZziE2IKcmlD3s79A/+hE8RSWdFSQVv7PMdTMDzWkKtg+K2oFGXemO4SsDSkwHDSjGoUT
Z/Ux0sYRXCGS/XaN+yZ6vj5Rq4p9cBZsxA6KfP09FChzabCj/mdS3aS92SZayv6brhJ+m72Ga5GM
vqYaP+bePsyuB9FZoTFlRq7+ufFheCJde7ixozxGg8X7jVzTRsELM0vJPgJ81i2Jj9QG6/1DWqaN
FCwhKkYJdpBoVj+NGVIdbte/oS9Fw7YtXMk/5ytR3VhHwmqgpn2E4U6o/1Cf2TsJj/BWaNtOA0WE
YQ3qu4yJzgexZI+1FtxfAg8MXQ3us4x3jm9WtClSc8O0AuTI/HKOS6ou2DOPbKoFd9V9z4OiyVAy
3ISBUe+gxAYT55z29yUrptOZ2feN2CWUWJCytGp9wBohjcwn7WvAYzozLkrNSLuBm0nKkDQCINTZ
zp+kOfsf+uGAU7Te1t8xB7aILbDu2OT3gK94E0bu445PTTIGGmg8lrEBf++a0tIdQKG6CE40JJIs
MFMIwUNFA4CASaSYZ0mb/twgE47MIojUHHMggJzmWhePRoC8ySkIil3Nm4asOcjevWDC2PX+C2YE
bOkgyd84TYdAPCNmWkBK32tJdwSqguB5FZ2eLJN2yv+rWJ5D2+ai9VJKIz7vw7zLdW8PRuw+5RgL
L8YY33j0RMEiB3htDFZxxc4k/D4xoG2amKK42fbge6pBVUppncj+vvYdW5echbrt8/NI1Dy2yzZM
wknfP1Y3w7G+4zmF8b6rWZcc3eopD0xdQ91QAaaMSeX6uTYsS8M1aqFvKthTnVyYhEfFSXTLaQdo
0kOP04H+coFnDeS2v33VU/sKOVWHogaxwo2wt+hyo+0LGtZJxLec2He/feEVwKy5k0xlmFZ3v9gx
nVXBERV9A+01R0v0U8VoDsY9j0nZUyhlaWFO0XlgcTFl4VVYL26xGOpvfYSTkFISYCvQWVXTT9SC
64fRzNwnEhE2BqAJLihsxUAuiEgCF+3LjnMu2uxJnUIpSYaRNWrKPs8Eohdl4NfFOUOHYLDTDs82
2n+GK2Y0AUchC9r8uJ5INfdr0k7m4RCdac3vjmIaX8cIc9cTNvDE4koVYeuxMndHM8oDoeuBEFrL
pHDH/bcgV5+OCt7Jy1GtiORkpE3WQyrTDgeHwdnoKA1SyydjssF3cNlYuDfyJZ8A+X1fpLELIb2k
wyJTLUOKvOBiIzEOk8CrYpooFycU3K1MHR79WVkjnbHhRSeLM9fSR64mpwhuNqdd24yCxiejCtbT
aDTpAIX1IEZ7pPrNUF+0BCqN8g0NBKRuWueCXTWX3r8CQ7ZbUL4tMPfOhBjbVENhxGm7HjSIbJ+S
IfC32Di71exQNhyD+97Zc+XKjn0sCeIG1oBwsGCdvm4A/trm8Bfh8O2hWIZwH0tcgHj6PLaDUk+7
AyP2Se8ruV0rE6Xv2QMwQYicLwgBAKDJMlZCg+vIaS4ifGRXJHOGWcgyH25L6dFixtt5ZLWkKUWE
hhwCd+56I0cuo9KTPTX6gv5RL4wSVtRbSZOwazLYCmMUk7swu2HaU0EIyq4pRCGYxanSiZGcYQOO
yMDy53IsamRjj0VJfB6Xr7Dg3OniL4im9RhKU5KfRjgV+Gxl+IGLQ2SMK59Peg8ibUX2aAF93IEK
scfiwF9EDJ5Fk9sBHyH4Fr4pxjt5f5uuWSW7Q6n3wEdaNPVHApI9j1I1XMgnFONjGYjeU9fbVgzY
VkJpVzDeNO4oFP3qsV6lftNoi+/h7PXMmx0/ggRTBbqrk40g5J2qjx1bcxHq3DkBgzXZef7aKiqw
/u+B52tQDzeNUVqD3KlVvhsAvQsQiYwg0tdTa50jjNL+JDmJAa+ikEgp3/KyPW5w4q7yve47/7Gu
eDjJXKidB8ZQ6YxmSlTKPR8jPA0Y5v8Je7oMye0d41AL7n6o/EKxDUPcE6T6/gPK3Gtef3Dzr4Cn
gVdXJicAqMi0sfU/d/HADg/YWsRFqTwyIWbtpbqDfZvSNpS7a8tP1vHYNGSfT53apKrSfR2QOAlB
c+af+a/yb+xXBRX5V83N2ioTi8uJfotE+f0reCgyddx0oB+gQHmSTwCjNsSndG+fOvOncHMiLZMX
Ppy0byI+RTl7Zw6JRlJUzpP2MMIkUj9vOkl4ny5QGcHEzOUfhn1IvmLr3wtS/UPwmfRpE2h/9tie
+uhWFQkWhNLGjIB0/JvJhvvHJwdhaBdN05OE9IgvoT2Td7gobpMc1NuL7p7imEAzRD+NSX6jXNoJ
Ygch+ow8CCIIC0PvBLPEmrcOm9HopUKLkpoT1zuUWcgB+ccaBS3EgsW4EqgOwWhrAJjtgIcKwRBD
RwlmRvifRRo+eWBFEEPtBThJmTu9QN73PaFcWDBVicF+211Rz7yoDYfbdLln1lQiE3KwbDw2LNqU
q9a/MH3ptUFLR0RDZtgKFQ40n1SrPwJh2u4TAMGIZmObN22TU4xbEARCpxI2FQRjBIx5tfQyojWx
yZvMojX9AwEUG0pv+933kRiGO0xn/b8rZAa0RkAEw9E+gzWr1oCl8hb1w3ixnMkVodxC8FXi5ZwZ
XXbD3pg1ASyweKV2DHifSwXRsLiCFMhFHZZXPUsUsuhVFLHiwvcPf2SWIEg2pAnVOgVOu9e6XnK/
PQKbfa5OMqbwoLf70fXCxThmdDDWdEP14RG9mb/TPITSVW6wN9xW+9hE5+eN3upVavHKj3lZkzzd
KKyMepVe5ndMeEs7UyAePZbkQ4TUuHzzfto/rrL7IK9jFCdH52zFpGlYE6jqcWRjFAsx5c8mjS0e
8L5iQaNr3cu3rBq+YOKH5Hzm8rXmKXyFvjKe2AJFrllOw8lDSqYbkfpS2DQrGOXroZjd1g1s03+M
vkqkKr5vNjD5tto0MVRvQaMT21H07LNzgMujacfSdo4ibIALQL6/C81Q41gt4qj/NM6z3AWaYS/T
KgSD0ZM29cQ+wLtXJFn7ypTh8eT6VFkG19Rft8ZSFt9BUjBz4cbGgg5LPsjLDcOU9QKOJY/kF5Dv
C+E4C8CYhgwqTlVBOzThFo8qi8znxNgjrvgqlFNibqmpcQoxuv6ROROR4Zf87V3zgxiHukdElIEG
mt1NRjln1D9AeW3b+AnR/DG4WorKuoipssFGlg2Ti0wPtMXuA2XjHBkYj6qQwkYZrMW4SPI/Y/5Q
cdwTJ1TB1eWGisnhrZePdDiAjMoCgFJGneDatd+ZtQEnU9zL9pc9bY2YtMziU7y5zmua4xOZdFLC
MSK8GZpjxicVzQZ8MwVIA20gpZlbQuVx+b/wcN5Oa3/bahs7wKD2qS8gqrcssp42iDbQvc130eSw
TdChP6WFEAmnrR7BchBuNPDsGROD53yXpQrUsNpp9gLnNyPZ8+piXitOLA6VC52ur0Mu/Qz8qKbZ
vjVlOZB9rpBWMyqQ26VvpVSdU7UmRR8PsCcJ6lUBsFuvWLVVX8oJi+63ZcJSPIZ0prAinFphLcws
BaX77VyGUiJjd+/NLpOiVh5ujBrBN3loKDBgc5iUolErNVysuSzH9G4T1EJbltOxB+tM9xqzl51Y
5T2RJB+PH5/dawNP7+vmaKigu85F2gfU7Ch8D8gwO3zl8DxX5BpGglCLiwMiHRhh7sOYDiTjxcio
Sq+u5kGesCgpv8vRTxyqf6HqfB6j7heAY3FWduJQRnJ2IN7H/DLvGhJe9kKHNB5sGqCWXPX26bwe
zpOdQoY39sWMJxa5DHhjeL6znznuXhHrSTUEWPPu14MUwEj6mpHTT2SBF4aOnOiGsZ1bI+wmZK6t
T86vvYcJ73M8COS5QCPrjBliOlCSNR9SWE1pMoFSaFKfnjU0ec4YC+mmp1Cbpgimm/nWQ9Y08/hG
1EoZ/yarYYeUq7CGU9BJLjnMXjrlU0vyiYkzJXyhwAaHRunUPHosHT/NDU1gmq8+0SUfDQLK0MRj
L4jJ/cESnt9pzz13t0q7I/3J9rK48qup1PQY405GJFwqMRLZE59A1N4H4T6pxp2MkWCXUF+OObYf
aGFc2/ccoOZlxH1eldQ4tuG16UdM3NmunGIs66oqbYOLWZZlKCtJZ11ZThsgru4kuORrcVKKvp3T
+SgM38kAmAjjbNUJ4gvz1OnZxe65kJPEkkbI/2gV+WmigNHZxe+dNDZoa034zt6f+qAmtV10SUSk
44MtYM9uUmcvzs3YA9HIWWN+5oTL8rPa93wYNqa+cTBh4FGRGzR3rAJiJdmlVW2icUS5/H8jMwN6
RG6qzoukx0v5g3qLY1oeO3FCPHZB+iELD5GSYHVlVJc572nxXfFv3H2uZkeqeuYC5YfD/i7CF7+0
lwLpKtgHYTefAPLm5jCJv7Y/0Tv87y07UTTpUMHUyI1rCmEQkNhRkyVV+ZsH9Nt6D6C+xnIjxO69
JwjCOKYnrVO5isHOzKKRVjJKNkIYYDC64KNghkwnU4sSeaReIRaDHTNtCFLUEgtRHNJ2wktFu9Yr
dIl8Uopw1immlqnxAnbWl1EXho5cfutB71WDVTi9kmKB81cwT82qo5QSd+ZnE4KdKcY5UbvUyK2N
1Uyu82GqSXnVVUUnpvUmuNcH/RZdZAA9CWk9J8JG32eJT2orX/hP63RcKuXQGPFNlOxMs9MoqmlK
rgERaKXDrzZr6tmMa0PFHZ027/aTLlVOktZ+oT+zrfFlx3V5Z8FitrMZdDNt0K5sM69DhZNTNWmD
BcW8lMa3JSrn+BwhK4VXtmTqjtGchjJnP0uXKHitOyFT4arVuf4yUPEFCU1YjhByyJaa1X6J4MDv
lAFywfltHqktzY2tK5i+ThM8GTU3V0yaAsbDU7IjtMm2tQLU8SDg0dnUwFMy99sehU7889bHSG5L
v6wSxatVmHHOXijwW2TfPYI5e8bdDn235eQD8a1sGVs9Zi7Sztm1650yPOb7ric9tfFk+pBYJec1
8nRQUajT0t5QP5dJC0CqJN1zbCJTy+NvkEeaWMDfjxxo4wcloNZ3eClYH4VZfTAIxUsleBHP8nK/
pv+boVGrNLTNKGBGlOi7QryHdrP3I/DWPV/EQbV19IuFTAPSasa+y0KMwh/sr7j4RoBXa8odsGgI
bn6M16OnX/pn61fkRDctyWT0/CLFqAQYm31BOd1EVRa2zYnz7x1UmnPkbFr+zu6Uswhv7tzATv5z
BuV34Z5wEZTKXH8qqz/SLC+c3fNSUIM1U9firKJcWwMqv/JwWR11jxON293PxEWdTxZhGyBzckMm
6UYO7Smd7GRlMoQs6bX3zBAFGf9o/erkhj+cNXFBgB70S77OF9oakL2VqAB6TQOuU7VCUrQH8zt4
X6yJfabjTLtV0CGw5pjq2I+52tfAECstwOzkrCDECmKLcKkMECd5T5+FWWRCLOQPsS9sqyWI352n
YH0GYzsVZpYeN5d1xfTlmNvA3ko02YRZ/MMXC1ckmWRZ3uRK63f1hUkGydJByYHQxAsyPfjJyatQ
s8d1j04h2Lln4bDS7Y1EyWYPeg96DF1q9j5ZOA4KaC8gRZgRYEnLd/BE/q79R//OupiVWyV7gCdd
P+xFagM9zTbF+5VG23hwW/NE7cgTvdGqsE98qjDzj3dr0eUJmV8D7QVf34WT8in99K7eyERMH3zp
Hrhp0kZB6HLjXrtiJ0x/tuw1AtKGF4XjyXb0Mkcu/BnkdjXlnlTHc1vthJLfYGE64F+DvKkg3TT8
c3KIvAcgLn69zxwdouz5JL7CgXgmZ8ypo81Mld5pj2qd3ImQvFZnmEzIfZ2Wx+m6uwUn/j3SBzCn
DnJ9m2uJZrOq6lLH76pvCwfT4rJn7j8+1Gyt2UZfMpKnGa7a6LTvWMdeu55hS4qQmrH8onBKUTcn
5Xmt6piIJaWp/Upt0L3eMQWRLldrYEKFR5082r+DP2SI6YFTOtDUsXUfyekbA99mFm0Iu+ghj3QQ
wpZe7ezZX94tnx+gVikA4QKja0XZr0LIDcZsEjpC8RXeaI1mKzg4DQGyuL4OXwykU5SUqqKdi1Bj
wXHIPLdphdFani/oyvVhqW8jNnKgArC6WkYh8ApGuqI/XKqfIFpurEpHgsB7m3PjrRupoWFqgTrv
soQ6QN+IqGB1yAKUQDEr/V9CibIzO3oKFdFKV2fDCyc7zvwGt8Hyv8/5JwaeR5kdw1K1ZFM7iNfZ
a7rlhxFFrm1Tu72cgpYaO1yTqra6G6DQm2376t2B+A8K+7qH98cqP7SSE4MaWnp4RnS9ynzOGSZZ
SAn515UGb/efzY46FrbcAZgcaS+f3vQiWbDcStxgDogddfTY+qfm3nerIJpNNV0dHy7vQ6JE+/6J
IUWYL5lq2Ke2oeZAW17AN35tQlAq7mPeGovFA1el31BFsg7kOiwCC9IAf7g88Dn78JpHbkLWACRQ
BE7XLtsU84n0pDn0pp8ELoplN3olx5i/1urGkJA4eketh2mzFRyH5D+El88soGHZ4A1U4f7kTkub
ttzM7px6J8sTH1HwgWzQznQ5oro+x8btRpUKmiqQHsVzhcwSq58bEbJGAg2mtGrfsD5K7uz+OO8V
rVvTPl9uHbcyVQ5jVYGJYab41/EKlIxglAz9OuLXT1E4xtzd2RVadUvykcctFwMl3JsTyDzfeddH
8L3F7T5KrsI2x0dbyVwkxyFsEqOSU+i2zpOzFuCSXnwrD71/QLnfTLUKskA/ZAKqnF/kQa4/okok
NIkucF3MZ4HmW5AMWJ+ms817JAqIqVsyq+/31en6H/4BflIiX8UaB9veC/MHLdtGa0xXIj9SKNTd
axYJRT3bJHmDDmcz0LfX8hU99C3VrzFobnIC8ulioWo+XU6GiVYDv96vIVdmA0vwiFy2CqDI/jOb
wJazEumIGFyHTEkNy0VsVV5aNOrXnv1FHPRh3+qujQDUdNWSSFSWWZEdwLrhCCkT+F0G5kSLEuUb
S2T8f8+Xq9pnAblCVy8NxV0BVRkLxeD2nhoRRt/j48/oF7WON2Oh3XSm7724snG6Bfmb03sZsJKh
nTzHcKfxli4eDBI7+Yd6aiJygUJgMiqv9NAmbb+3/7dy5RDSr/RFlqxaFaVNWhZM08Tv3td3PrVn
527R0CM6o2B0jB+IaK5wZIpK8R1ao14GacwEaSBe82/Bclnrnj+USTC3Cwj9LJZi2XsSfX18J3ks
7a2q8w+CM8Kic6aWVo7yLc8EPSMy/BKGXjuLvKj8+VKNCgq+U5+mKfecu3DQPRNpK6SSGDhWV13Z
riR0u1mAxOuWuE8HXQk8pBzrmSZHKan8Lw2qvblcCXg8BKBhT+HpFObI4Mfc7kablL5XSFDC+z7c
+l7fXYFEocNKdxCxFsF58lLL2AnjUzfwe5BlTynzksgq/ndUY7TIIIsLDHFD1WzVShxUUFYOE1Es
eE/Hcje3/VJw/i4efxku8pyLULkeKbGJkdGwqDQinOuwXjpwTeP8EPcG/mj403NVnMrKfuxzaPfr
VcgjzkHgIb5RHiioUbD5+BpirvwtTLQFQtBnCsR5fEKwB2/zGD8omm1Sy7kdLi5v2szVtose3bbn
VcESrUWlMSvBxl7xKLlFQF9gEazOz8r3ajy3BTmdOMupIaoB5AldSC7S8V7NQFa1YXStHKgh/VVM
w+bd+S2pQ5QGx3t1lHQEXhZd9gG42459X9l+18f3zRpKNfuN2mfGkUdd3qC96iKlV188FHkpc5rq
nqpplERmHmGGltOT6953KU1OZHdnsBDD9wx/qdiV+wBZF8cOVcI1CQeax+KtdJwihYOZ0EckUbPY
sdqRUPaT+Pb2C8xqh9B0UxcJuvHymKzKLxzq2cEVewNjBpUIa6G55/W0rLHbvmM3YTwZ4b/hvvEA
bdh0KODhwc9e1wupHGqMuaY+4maWKKYbuTUwzniegIwDFWMdsiTruymqvZmmmndvVImGAUDQeeR5
vaKP59ILbi6CRhNgGxnN0yvbT0LLHdLG6FeY/IGy87XIqM+DwZ4ld8AVo5QvOUio1VyeS/XSBMhO
N+GeArAIlJGnq37Ksb29q/mmsKpLA0oNPTfkw5ZhlMP0z7ECMDZOFM74p47rJzSS3e0Sr6XbHWS7
CniiaSNEcYqS69gwJ2iDfbWsauyGrJbj6TgiwnZ5CJ4XM6dFwg4Vnzd9uUZan4CK9Mun/73uiiZT
9a8gHFhST1rGhJ2unwFwJzNUzkaENZ2esSBeV01U0yY1YZ9/rEnWv8JW998zwD/NvjkPGkUGhNKI
nHgKsdILni1VpXEig4vQ/0dBPRP//LZb5Ksig4J7tYF3G4UZ64cQF5GhJfZmA5fquUKOT8nDKr4U
6e6ETYsGRE06fIhUMMDNTO3wAokm0UMyCe3S5vgS9erikLtD/h4kAqL/95JnxgFaCq/OHlipQSMf
bAcVV4fH+AXWHDfLoHM6hmVegQH9wDMwAXrWVLiLkiIW93mQOfSwzw5BD5WRhJm4cRDlTqfJiit7
NfHmlaw+dCoENHoKEWt47r455qWm1hj5oSGRntA6YwC1JmRkkEqxRp1xjhlME/x3P7RAPSj52W+4
g+EOe5RNpcdHIOSl4s3y4OkXCyaiFk6XQLg0L8/mA0s8VN/CViWcmpQ/6UDhU452kWs4zOue7rwA
/WY3k+GVSMnLBodDoTI3Ah1qWcYKGPjyKAf2yK7lZV78fV6JyikqYS9UV+VkKYSg30V/jTmlhW4M
9TsKBYWAdmnuQUHRrtZs18kQXUIzrOsHS0CKP2J9gvRZyX6yqxmEMPfkaOnlH0pZpEy5N3x1gIyg
fiRH+MoBnwpY5SH3/iNEfcR0/PunAtQhbxn0FN5yZwQJwak/XOY8IdkhJbgptuPnJv2cNTqr5wtr
hx/nuByWi1Ap819N90CKHZ9+xCMlypb5jabOhjaiFvRlqavIWh7vvMjQtk21ccOKr82PTUGR0uPH
5/xPaEhDRfeOigRAtQ0xYs0pmfJfFJ7nBvGA/hdYkmV+lcv0kk61n77TbOffkRWTaqiijrQnvxcB
FnCz/Fj+KQ7lapjZdPCdSQb2g5+LJ4lWhtmbcAo67UFKX/zrQBxq88qF72QZi2i4dWX+p9SD5Qfi
zO7JK/bovzqBJJhgrpwc6+MesPTZ6X1mq/JBxA6F7N4cwLGjkc/4mv+F3CG9HBPvm1p5jmJnRvvz
/aryvei4vphWxHnsfq7W+dHDQj1skaA6FeCob4PCV6jbXncQcK2ncFYmRZA0aOZ/s1uvp8P3RRYY
vqWU8bLFPrZr47vEu0GXI6PRusnn/IEYXOmOPsd3+2DHbNWWvSnbqTBgXTHYZH+5iSpRYi9v84Dx
3nLhNyWYW6bBcRs4Zx8RxyrSO3eFMH/dxbT94W2uX/lbya/BHVz56ouWAZfy0Kdgom3zPwKGo3tV
q7e+Li3JpxCOXj/S1D6WXvdev2SGFfI90TApSDzcfhQJaoqikKAiyocaMcfnuwlp+ZlXjflt45iT
l4MhMkZf7krWxSTRVoJpCcTRDdJz1tYUZ5P+cMnoXRKhYfHAB0YcWWGw4YP2kNj8k8g2t5B190RZ
X0VHZh2kRTDoEaYFkTWxlMd5k4vEXKSJ0V0Kh9FEkJ0+zg8axzhx+B2qIYrteFmNu/4sWMEyicAv
Mh6gbfR2kyNVoAd5IhGaPfEJ6ScfLtkOgFPLJWoIJcQBbOiniFs7IL2nGbT5b2NplCPhQqR2HCbo
pRoxFC7hl435nU/ugW5wKoURgjySCtaIAP7KNqkxygQ85xJgWV1U37SFCD7cdEwFflHwjF4UE/RK
2dkMm0Zo1MLWIwLG6a9wEryD1aoWR5V/xhbVmyCr1/KMXWYFI8aWIlfICD9jwOJN4xNKhMivjkwh
SuGlNXNWeM9Hdq+skN+2DPYjIN40WK/wCPoa8Zs5wVShxbRefCN4SRmEceTpaCV24dpQuzGF1/Ec
nKlyrquZzT3LSkHGHs2kel5MhN3HKHKkbeUIJg55LZtL22rQ3cOmlvedw/NCSNvU9SXlBlppb1+c
VwjIiOE5zPjltqZizLElLeEUTJrvBFOil/EKEuKQ2GZ2x7hL/Wh9ISVla8ef2t9mOCfXeKbqL8CP
Bw10+MUlQppbz2UOyaGPd78yO5vFQFgSDGL6n2NoIPNdTx4yHNNoaL+4OUhQC4J0kg1XyXvsJBDv
Dk4grYR3LuwlMsAKZ7GMuDY5ftUxXGBZZcNm48QU0SfleSdWCwfSIt9/hPGDVKigEJeI60u4siUj
JW2SzUeJQAN/P83rqyc+Q84efzMWkcLMQ9KN0PEQ23fhZXtjfPYFvSA6x2zmla8kGbmblwKmEjhp
dpS4zkPAEezLfcnOHrkDfjIe2888gvHQO6Yl2sXlrDDxE1rgTJIjq/fAh7i8HDtPKbbfDzwxxh17
r+iWz8a/LZVBxlRc/TpPSY1ucxEeX7M/fKQeN1xrXkSdCQi2KMxgRi0czbUCgiPBk4C2m329o+Yg
WkeWpK6GOG9stUpPX80Jy85LRHEIhbbfloJAvPty/ns9yW9QU0rDPUA2msgRSzc6vLO5qixsJWK2
GF6j/eI3m8UF5F/9XLVkYVW8MXlGMN8giB4b+egPYkj34u7nwCx8AsQZdmmQhpmP8xNPZWyE6mLQ
eLXemutABTwpzxPGizUrVzZrTRHHvSqrccUmRBG7mfHI7s1jnHFXP6R+kfCKy5s16Qg7AbO8DeMX
jQaxeWwlGVxostQOU49B3uEiC40b18YgElzaoLy/vuc+iAMJ5H5Sh2f7CY9uwaXm/iBFJQ0uT9az
GbxOqFxu+ehyT+3I2d6iY06cT4GoTBuGqHqvmbNTYzcSiwCel33mIF5REKhTzekzDkpFnFwWoaCM
jZg6bXeLrFscUerl5/2dWwG873yWbEl4If7rn15tj86wyc6JM2nVAGuhM4bf3C/1xNfgv2+AmyDK
Ji8U3ABBeef4kapo92d8JtBUnLd28vGT8oiGzPx5CN+M011BEHCoUAKimx9mFjyp4orJsNHsqp0h
Nizj+x32VBCynbqWeDfroGwooYbZE/FAlfLnIXxqnJPCI0SpFgm9+n0TDq5iVsyL7CdnNvnHS+Yw
FDQiiuh+vGE7tVcj3g0bT//Y+Lz22I4o+4Sh8zWIKio7pV05sev5Vxh7oydSEfdNpUqcixy4rqeH
vOt/9YCCe9c2GZeyd0v3KNwOdHS1gIUChXpf4yVwzL4kQC+wG6c6F0a3fNRHTBGzO+Ye7SovWOX8
0CqcinUWimfMW1Btvy6xpwmkr0dqTHeP4gkEwvFer1QfNShc7EUoySAe4pXJKoorHHyAtxBWRiq9
/MePvKA8xfienH5iHda6uuxnNYYzLR3irlgpVZ7ykPlL4PtPcW6azCP6l3oJGgsCgL+8WFygncPm
dme8MGEeoNHafUilFKNE/F5+kNrP1X57peNvyLUzuZzFMmqAS59k9goMmXcE6EKs8eCGncJveg1l
flozfZUMPVOTSTlct2SnosoN6qqad46kxg4aMdGQOxASetneYfLENnpnLiDh3KcLg9SG+lIUf+CP
XDoS+YvEnsXKMbLNM4lTjAOM7sUbiFmLB9qa0RNP63Zvvqnl1PBLRp1tHovDW185+f2PJxv01ghK
txZRWZJpfJazSRcV9EUiP/47gR0zpwqwSuTIS65x/d4iuWLhCmiLrmO6oVglaqpr5GM9p31MJ/n7
dv9US/FR8muk8E0jNgi8NY0KelqZUUkL0PwESyqelMQfi+h9pY0VhYM2t1lqzXcsGSFR87ewQkej
BdQNoUIBctD4yupTwUJc4OrlnE3/VuYljctflHvuBCjNaa0grwAxHsuTuWKoGO4RoVAlD8oRDk+x
d0MLi2HvODKGgz1qyxSxHfsCwZ/xbfaQhCGwjjDeyp8uC764D3T+A6lly6S5flFmiY6VWhOoAgE7
cAOv7MPxS1wN79N3pvX3PIl7Hp4Hc3rg2BEWR5CmS5gFyRT/g/iNr04KVLY072qp2DNvUWMxAlEo
bUWP0baGJNa3LUCOhYhs5MtiYJyKxwvuT8rAtwwwaE5kB7OkwUVF0KhEdnv9QD5HfsKxjxCOKW8V
beHUTPgNjfd+FF79cTm+Z8bi3b7dOuKqlVzFkYjpvod9TaF3Dgaq6WC6Cn+zrvNtZz1plKG+btr9
RNwwWo0YXtAnyGCvqIDLFA8flVJgVudD1uSeFtNLHuuqsmFC5iTm/8ykYkpR5S5KMDAPIeK4f8X7
zSfoG7aButoNRmTzZ7EOGpXlbcCCMePF+VDNEzvhjkPLH0kfoqfqMVQBttVQVn3eIZ16AImBdDTZ
eJhqI6ysmabZhLfguh4az8J6B6Ubwg4l+IGPbnHyVzj/HDe7ZCh1rwVz1u5ieYN1KyuvIns+7X1f
zu8ZIPnc02sf3kkFFXXOvyfzwBQkA/oZwXeauE27BOJRobVt/a6N4OB0qxShC+t3ov1LY5SKXdxS
43FHOpKQgoDBBPPlcYG1+IQQ9G530zueAMHx2mmCx198+x8XTMavOS5McL7CdNxWzFCZKX90UwU+
BghF9siLwnEjK1MV34945y0II05NtcACG5+ucgCfobCGN2wgjC9cAIDJHF3JZDXJx6q7tjpJH65p
dGJCCb37AwQP5HCGmDcNDsChjbQ9TOjRYB0WVBrxtP3GLKLIej41vcRemCPyEuP8dwWDhbpJhhcO
GVnZLbxOt5n+cQ/Nm4ezI5eLRaa7JJX0VOzmmXlAPEDQzqNelph54bwzMBRpoS1x8RrfaC0ZA3PT
4Py4U6adqWuThvhw0JCytiSiZqHiu2RXulT4bgy6NW1md0MvZfyr2Yvhb7O9gDvMPiNDecsUxWp4
tp4YjOXnUFGCkjrmYDiNI0j29lX/gFKwb0SSaaLPCeRTLwa7VEYq64J6DAOMcnpUsoi8z9LAPgNE
jWueh70t2QVZczDbJ7to9OqHNetb/Mp5ivMT0UKe43d/kl+46i2d5I+Warm0GRQqly6hoWADNwzj
dUY3yddhbfglxPl+bp7JxgHcpmFS+yQnWdYYakSUSX4AZCdHwBp0LLeTmYHqDiuXnuXONWCT7meZ
39tFF4KjkWrSn+82pYsz6Wnvtcv0xoOHuhKHpkmUMY5eRsPRbaWdWbG6XcAqjKyh065SsOk4iXTP
j8f88mN1TcdTGVgssPogl8NWZDtPpeV+5sggp3OcnSJ8NOWuAsz8dP4ksO0pWYY9mlmob3iBQ85k
xICZ+65E947qZ8m1lwPrTItcMQZ0ulYY7u6hT2RJSwMDlyspE+6Ow7ZGInOcjz3VI2GdBmnv8I/N
lBQYd5Ktso8fdTXoROLINGeQKD6Otaj+Qb8njhcHhTWmnPt0fkBnn8USTyB4bSxy5TB6ALynYjVJ
GcFEA7rClzsSRkOpsO92x9gGn76OmIxviFBkLX88S8Se45xgQ/C6RPn1cRQP4Rc4IwEBsqQIOayy
+svVgAMfrYNJY/Am2MxtPgs2p9tRkUtNUpu6VvuUs1pOLl6BRVERhfTx2ud0EHzp18MWBNxv8KLU
CiY0IGrZzZpyj4a88C8/nXR4fz8yT+uSOyu7mdRnrdo2NIWDFE1FeJwQtcEPpOuhz0sNACWMp5Et
UIv/NMIhP+m/uPWPtL6HMdmAsrmyxz7Od8+uw8jKVyspEGXbrjztE29+16I2KilqTaV81UCWbVty
IO1dWERu1JEEVz643+yJjva3Otr2F41F9jB2p2mtsdjIzCG7ui0bEkhXuSb8S1cELkcbwD+0sTTW
y5HYbQ16Lp7jMkQFsyadh+t98KA5sgT8OK85mGrkGJPTsJFjo+YnFkX+SsoaA4b0QN9i+aaMM+Bf
cUxcU/kNeV2rG7oGuELr9PB3B7lVWhfjHa5Mdl9YasUAoaMy2GFMFFvwv+jHknGhB+8B4K1keUgp
JgGyq0YVmJOfXSHsfJ3DnOqv5yiMm1CB9lFYWpZy5n+uOIgMTujWoRb480Od/ZsJbTpJyjLPvKcj
uMz/lthno7voFLP4WprCx4leRznPkLSVfmF2c+L5zMYqHBZ5WnJtL3f721vq0f/vAVv5jiWlgFoc
syqOUyudp1fkQUqgMG0KY+vLvuzpqOUrm4Nv6wEioOGgwKfMAeZ/Wrf/hc6VWVSLQjhzOS3FB/CV
+MfBT3vXSKZgzeRc77VWHwI2SrnySrKhpsAz+cJNMxY1Ykz9Zhi2kWnjqJoLHY+jCyCZ8Qj8BNDE
PV7jovpjZGaOMdCngKF9YWwPPB/ei4Pm+3omF/HIZnojpjH4zzJ/C/AaqYmj8S7T/maBBMJtcDP1
yg6dEYBjE6YiR0hRWjiKpPe3EUXQAfpqy1w6bThhTPMG43sW8DOCvVKRuEXbNwtql5vgyTlyEbrR
6hzx37TGF1+mBw9jmCZgAEg7GDaYo89PVD/QOyfk9lo7ckx4jk1TF8j+YpNBJE+6z+fdb8fNJAGc
I1GR7PKC2hZHrLxYLw5jK75Bn/J/0xn0y5XrfEagMabZEL8kHr3eGwBbs2AyqZzAb4L27EHBPyiI
QEiMDve+pcQqpaWSxePsaqy+6DuHx61C6dow8GckQXEyJMMJyeD81LR32VKWFpph53Mk5Z4AIkR7
DnU7bxud4NlS78EEb7nElkFSIBq9IotlRrm2pzFcgb3hM+hflRiIN16cDGI5ExFC+b4P714NDLTf
7SFJWFCn014SI3IUEuHFhE0DhsHR8aJzb+hyHYHiwogc7BmdsyHio2IQS1YmHFbsQ2KjBweDaaaU
U0VeNZDR2ufCnD6t5u63Em5OBO8oUYPHNIsEwoUAOKKMYZKQ4JJV6qRlcTED7iIaRR57b8maSdXh
yE5qVZOW6FQjb2AUiqTJXlz+AcL4PfTS8nxYjQ1Qx9i9z42+Pj/YEL6LiEwZ7jkx8nym6Bu/f+D3
IPWADWQmnWxGCbpwW0Szu8qlFaMSX6ppnWjoN72MdAmtazlO3D41FLkilpNx/WCQFCb/ylu9DToL
3pXEfgP9Ca317TqFJ+y91mzm7mcRT+oUa8l19EeW5CTVIjPXrHup9rFvO830fFRHb4o1g/nPySxx
SIJwehuyIDUf3MevSW7dd2eSFRKRdxjzopQFyPVAfvEBRlEWdcTAiIRYzXQA5548sDstsF1VemAV
h/8S9B9lTHwPbX37XW+4FukYDr2reB3iQr/VwUdwow1bZAAhpr2qObQ0LV7Hmh5bemG811voXeDl
HKk2A8uoaGwSbDDt1JMj2ULX8P97OEIa6J77I510zkwbETS3rs55WQf1qVZy0cGLFjqtK4HHOyGT
gkIJT0fENVbkpNCwA4OZkTl87DDmJAfeI2/jpKjQV6CR1Q+Fc2NG+uP16SrM6Xh1Gw2ojHx6R6+a
pP96xZWqrN/d7Sj1lS0BtIadyzLjcoF61XR3UhIUsRLtn5zOv/7bLSiVW+jNqDH6+Iy6VTxwhXaR
bj1ymXplazaWkDg0YuuYwH4Ip0zbr9oDdNFvRE/tn8Osr3EmHI2g0wEnsT0lNi5Ye/WrlrsgYCXN
QrnGEEWPvhu0t9XjYLlqwHQ0bqXTVdePvQg9Is8UQ4FY0SLpeX0KWgihzUqAC2Kg0M2/bYXfdB10
LE8JC7NiBofjDZJbvIY7w3SwrEr6NiF34NrgHxNCPpzp8p/eSfN0JtECL8ht59V4/2lwbCIzKtvC
yU9bG3bkYQU4swAinVM1HC6mMoWuJ/NQaKlvM4h5EhiUYbUkOEHlVXAFM6G/7HNPCwnpeTaKbycb
Xm9gSkN9cVwPOxPOWym4doTAImynog2ucjEmaQEKoOz6Rw8SmtKER+6MJztCtuzuHd5+nObLvDgF
EamQt+o7RChvf3aA4bB4z9CndxuX7hce9Fgh8q+wkDgHc/+a5gbZVPvQ+xhBYGTlXnAdMcsd/iMj
NPskhbRkX0k+ledrJWXqHKVY62Nailu7mLbF90/pzbGS0LJ1ke1IuVMyQXxUD0/fpYDVj3PMFDLf
hsxEaogNy93N19gwEClk0nTbi47nNRRItTCjjX1dgFZxzrVKQFMKv0LzxUfuIUFDJ+WPWiK98cPa
L1asfdooo79NkVe5+oiITTetkuJLHOmjBu1pMf9Dkqrmct48kFaU9BmaYqyNFhoMBgdq9lWySGh2
O4EKkkv+oUm1UotgoqQwjyio8JjgfQNY5Aqk2zJ2pb7sGpB+8DBKFPU1CKkDUIhNBVBNI5FDrEO6
a3TkHeVFcZJumbSSVU7iY8z93itlRnHskp8tdiuk+LLeKW6nyZNirvo8cMviyRJSiwnpOB0c4UdC
odfG0fJv8hAh47c15Uzc5hJLZVtyka20+ZHodfBdKlCmIBRxZZhLPCLB9VSnsCDCNLAC2bqa2EAi
u1IwwMtG0X3nMMbJSR2gGIPsVrGIlErT18A495bBMFowLIq4AccVQqhvQSwY3vXEz6kIw9z1xRQu
PNVuHSkxGe/YWBeH41CJi84Zm0jCW7vW/bpQBzrgg4Pi9bDokEl+NJNdu++EOxr/614/kTFL0SMr
GJFVRIaHE0KSeUgqdpa9rdJSmh+Ug6n/vd8WfuTyMbNjLNlroJinjYXLq0wewrQZ3i5kbm2Wuwxl
ajpnddIV5uIohbbKBzdcwmM4lPoA7Pd1dakJO9MxbuQR51vH20147hFKxDMv5FtlWIaq1NqZaL6y
zRRL+lE7pve9LpOOACFs+WgnE20NQHEKamFBUVOuCiopVqZLyitemyfIP8EPLTYNagU+XhpDUKMv
6pakt6G3dnJ1U/DeHBT6FgwkDuBqTAcXMgXHT82SRZZdc2MrEZoayjW1LXZwtuJMKftE+2Px983c
7DYTzVpOdk2TSg9F1v8ZcZx+7n0bdlmsjgTDcMo/huFxGYdVRuIXJS2/WUtvBKs8WPsbv7XhNWRq
eIKcxNlWrvCM6JLsvZ33bnPgaD2IDicuFlEYbzqHw+zk569Xrc2Unc3IGJZ34t55S0mrVxIyu2jc
UF3FWns8g4Xus6A0viTHTAeQWt8lKxdGcVaT5jT6xleg3+P9vUEUytZCEWQ3pdRxQygRf8AK3qgW
VBBQ5jUA/lYVkBbbaK5ZD+CjNJMl6Ha7BKsNGxumKnaMEkqwmEv2amh+aJlrEQ8ZKjJpD8R705gj
R0bGE8edThvQEtctdz39wyNEIChV3XRiEige+ffOW8zfPX6YyPqTlWhcOqnpzv/45VNEpaHOGvH2
+Cypy1FwjBVCbtFjERJ+IliLTVMgRSaz7o5Vp+zdBo/diANHTbf8vWsuLcE/owky5Q5yp2vOvvoa
0oGC2IEkGpyNkCQPD+kVve6IxyIj7SPBJevrURMXAy3948XtmalxjmlaWDu0tU3VV8dITWuSVGlg
nCvQ6DQhwd0tvHgz8WEeFPmao2j7DGZ7gP6HezW//K1b30nJ9Mav38p2PMa7d/r8mgahqaZuF9zy
qwuIDYcMhwwBC/+hJa3t233STvoo8WUyT0vtr7PxGgj73CjjtbWS9M8BUwP0s112rrLA0Q9jiXA7
L2dkq+5bMhuN81rwSHEGe8Yf4oYDAyLWzSahqamL+J4E1w5fmeJbZu612e32Sj7uH6zWPvVQWJ+8
36EromBbx2vx9bZMxZCgEI62sXQgwLzgHV38ZdTITCFLINZ8I4XnJFxa2tgBI8zc4R+H27/3SeId
NvL3ziwUeW8xWXcwynHr3nf+0gD6lzsJPk5DoFkiqKhrCIeKWf3vRKA3umdKQvux1GwsVlWaLF+3
k5a6vOb8TcF7vFzY6JOd2z4YxYQjreMINyYbMtNeBLurodKDytOKW86nzXBNzOJLjawftJRLvLDQ
SqHSE+sE1tUPuA8VkV0u5lCpNY2/Q1iCxOSW3OFhDzz55ElQBvpkgeROykIkNktiFVjYTJbMijAw
wYEBJ1LQa0mOgwLWtL4wShIs6Rh8bZ4oh7Laon4gsYxZSdlI4c4d9UM14KPH4iIIzGxLwUICEQcQ
Gkt/fNR0gipIZwVWZ+tNMEeNTk1m+WyeuCbPijxOtKXiGg0xvR+9m+dvx9TyRZRmMtaShhBDwcCd
7XWgYZRb+tktsHUQ1Scyoxd2eznT5HOdRk6WCtoup4bVwmnnb9owLBtHYljw/eiy+Us4Lv+2rM9z
umdPdr4n1YWOL5IOazX/7XAOeOpsBEfpcoOuUMZ9lhlRnKtMh4PPb/IO1qd5PWkfxaA2La6+Szuv
WIcgIwH3hA/DOs3sCfo6tJZc7M5tQ9cTB64bexA/w6Wsyep2gK+Y3luuU4fXpicOc+oGul6/98vs
7d6FyI8sHEPhJ+nA5mt86laR106ond+1J0dP9xy8px/qffalvrS067R35+b8WdayskdwXLuo2oCx
RCaD8re7zcf7AndCh7gEUf0LNEIrMRA1hPO1DOqvZ2bq+K7p+K6JUfGZAgnhZEYxJNv84tRxvNPn
QrgplZdcE0uJ62nTJOngr00TEhGYygFUxj38KW4hFww3G3vfa0T9/Jvs4i/JB/1mejICKdLYMkpc
O1LyyL+srGtR/OFCwrg/0yi5xiaBDfNuIPa3Jy/D/QuJS0aWd5ZY505KDjCLlZ/gfBsJQSziz2a3
ZispGUus6P+aAj73VY+Yt1HQ/kFelnM5xgWt5a7/tGXlqvMzFPYNZBDroNPHgDiywSSw8hQEy2ys
6n/Ck1A6D865BiLylVlJ5X6lXxqgLefjDWcTnxTcfmMF762Z8HTks+0uxsLmyXBZTcjaDA/P9UI6
HgAKJ+f0yFqj/GE+mNh1WdX0v+q5Tjo2pcxlPWHGi6bzyKlYjl0OZhWhV0Ft/o3Sa4tVFK0mnF7w
eUgpjj8oxZT+31xlzVSIidshsRZjqcTApn1GGRBSz+Pf4Rq9/En43EqonUNIszi1NKcbX+iIlSsP
IMy3sTKEk4rxYnlReERhmnrJCUu8VqCthK2/LO9ZCPp+X8tvm6Pr8Ze70Wz1Ho70TDSnC27cZpwO
IROOE/NKHQj+P3dVk9cgrLdq6q7HzQJnpckIJOI+GW2PTNtR3eOJIOXorGga1VgeAH4iIzWIt/SR
KWCaeEBnC5RmF6JQub7ianTXGQM9WiRJB8yp4B6n9i64NBObkKF3XYQzgKhJ1mlNnuyhvqqY06B8
PFzT2/KJXshFlBDf3y2x2tGEdSkGj7NY/4ixTV920NzG3ari83ekvXDxFXD4eQShSdrHCUa1e6zl
VFgXuGrBFpe7pZ2r4EQWS9gtYjxko20oGAKGhdHtYWempw8Hg3UtFk6XPUg2Wgxv7Wfxojj/g7mb
0yTTvYhCWOv567oUnU4rHZOeWkMI99T61ciR7jRrK6l39oo2edfohwQmajDY2PDbcVzkE5GVTNhr
Y0+qnnHi6d1qAguNQgMervcgLxnZjhgmS++zFP8xQx5ctGfvMGLpJJgBA0gt6YU2T2Z7oexFvtCK
J/3AQlE7BFDLIPoxSq1p+JqjIUmgZz4/4F3feg6Zcwv+kXY4u3xnj8o95IRDplvO2brr0Gbifjet
SbXj9u7Mn8sMNoYRStmqpa8uGk8CguwTb3kgSnnpHPvY51PlZltkoSt6wtT3JQ05WScGAEhyG337
fwYa5CcKvu9k82ZH0WkonRqAmeRt6LxzSXhemBckTB4Up60A9k1EWSHpTAWJ+CVYnKIPX5hrhV6l
DJgTUoc1rxg1386ajgGYWYVDz8CwAgjYYrTq2Gmu0J7s1n4dCQChzAgRXXQC7zE237ssQCCKucUW
rT7zXfUuVCutYJlyd3xRSYdP/DS3HKFP0zAlpxMVE1cYwggbWjAzVy/nDxdJzfdW5UqgsrYdD3O2
Lz32tci8hgsIm+uptbg8S2CJ1O57PUNu/4EFR5HkLIqUAGbZsIRjykj/FMpctJDnKNX60uknP53T
Mv2s9FwL54RlQr/zSRhSbicrkvr6y7/LtgfkOFevwNi77B7HCfieGJ8QmQeqCs8C1KpPYcq/R071
OydhZYS6J67rDa/aqM/8zys23oM9cp75d2zfHqrYMM8Z/lfY27K8a8SvfJM3Yu/Mx3QS7MHkOZWE
jncVjmkCPG27H5KUxNShlht6ReoOSBE0mo9tmwWjTmhUq5GcI+6c4jmD1yIXD0w/jrPlERBwGjVQ
g9G9oZtTG+Vz/Hg8cCkxQwWF0+xjYglOr2o8a3toP/NSNQ5pOFfbyr163oAmkGYto7aiZev99DVy
4wZMMwPUQTRx8vxh7seLC+AE5HrYl9/stqu9bCWWZyqkRAluLBXEMyBqQUIDa3Odj1LXB1+5813r
XgKAe8OehZ1/SPea7P9Y1vvkKgYHsCmLJbrze4frMPucQdvO9jTHpopManb6qmIiOaNw6wHxMzzZ
wAd5S7TjcLU5SRlrKKB11PF7QivuynSarw7fqSVc9sKa5daY57o4Fw2gK6eLn8ZO6+ruyNzIjjCW
ZMWPmH+synZJkg5O3S1IZwnVN0MSbArs5UvaRzfGySvi3TR7bgvXXN3l16rTmLLsVsxOnpbKPChR
kZYgH2X07RejGkYSDh6qYu2LDx6TXPbbOUCuOPDLefCHIbGNCBgaKSxNIElM7+KENap9j9IBdMTz
6DEfo3GRzK2j+DBafDzzmEdtHvRxa9cua3n4hxpOv3SZ38pxhkHLGRQfNSjyXjD4sErP6ScPIAqk
tRv7k3YAVW4wBajzv6UFLfRnlxGSvLqRRo27Yh7/kU1mjgZQpbH41P9D6XAHoS8IVF6TYUkaX0AQ
UxVeINPUCrlYMQi0CZCtrfID/IccPgBXgfyzirYJPkt00cogDDNvhFaBj8ewrtD78E0NVUgA4+CD
mfFT46pW1FBSvVjs82JkqdhLQQVs8PyiUW+WTNpyv33ZAXVs7kyYx22l6md/HUxN6k2ZIDaFjXsX
AU/3vCOsDrBk7kt1FwD+zko9o2kxovcSYar1QwzxT1UxWt6qcUxnyb/MKqiws1Nfw3KnWMaRXD2l
zrqdNr4zM+iyeAujGvBJ69TO27qI3UuugMxiGcfpe9goC/rZP4QLpwNpNItuahb4X1hS8Zg6FTz3
zYQzGIXZEFbIZhz6S+UMDu0jcSh2T+RwVDsublaxS1Y1pfsYj7A9QngFYaACIz3j8ntGQb9Oi1aQ
zlFWTwpMFeV6QoxOTxgf1vpyVgtwmbbQUnOEV/tn1TBzCq+zh/XGxs2hADnXAz0LQj/h5LLXk3iv
jBlV8IyJtdcwdeEJ3HC/6Xp0kXpqNk45zBzcnbQs7HibirGYOSooXWBGMKRUG0aZZOccZmxO3fE7
GKANvnsZx26dUTgbQYTviUBPWzef0Ox0dzerpsbBb5cbKwvAvYzXlDWS1zChomgrEWUZr/rR1A+6
vPYnPy/Ds8d6x0fC+rYOLy8sAnj+XHBAWVNSXuSp0iv69F7JN176OZ7lxbdAbVd2rpvmbVxZJdld
k54JiPOdIUZRM9L+fUHjySlYA2nkGf3Exs+fjcuNpKZmIJRbfdC4UPFz4MnP8oB1u4mgAGd8PWiU
T6uf3cIiChD5C8cLeoz4UvcIP8s+RlkCPVzbf+ktyHBiukNF1y4V/RyNCUwrSMIcEGd9E0+7DecU
oT0haFkoW9v/I7ngKOq6811Yvo603WOiy3Q98UitRLtcv+Ahi5WE8QTemU3Yxt8GmmqRMSxVKYBJ
fVt45m7g8D4+Nb0MXABl6zYNM3vM50FvbggYf813EYtgIyi5BUpzR6FtKHkxzVs2+U69oRbXymTV
CYjrnJ3P7k+hhSBAlhj4rjqcXQh/pe4kcIxhDZAdQU3MPs3qnw3GBGBo+QQJhPNTxNxSg+2WEV8n
0xoC5DZ8YVPNirpBXhRZT+ENJtRSWBOdyI+alUDfwyWb5p9chWkdARel3LiUiqpHMQSMbVII+kmV
UDVlJEL+nmkWgvee2bfkQ/R5FwfitWp+YyrPYozNZnLP0bmP6I0WR5UZLL+X2m4AEpjL//KnyB+g
aWK3JtCnRy43LRqE/dQN0Wbn8cTf/64DHu2cPvA7u4B0XphSUGE/+XgXUoclR0Dt4imhFmnPVnDO
8vvzdpb0tjfzMFOFmkdtj/lH5q/PjraKL3oet5VcAp67nsPC8okzOPWfYwPVlhllIP6aDWWD8Vjo
/srkGKADRD7OjoP5cdouwvUuZynse7tY5YChABQ87XSEvULS+mgShkOLPKz1zvPx72tErqKgo9kn
O85E7rOj6n9dCL3zzKxYD1i8iFFBZXz05O/YlSA5ZkaB8lzgJzSWt6Cn9Tv5VMjKxD6AHy3JJ4gw
xRw+g01xo/w5S05qHGI0FNHbG++ppa/lHMd1cOxkFzcJgqVd9uEVVLCrhpnKOfCWWs26au6WoGD9
pqQaK9vwu2cybZBZo9PpASyFB/Ilr5ZUso8bspPENf/IeOcWuXj0iRC6xE8ldL65oI1v5Z8JZnY4
hHz0nVe/N1H7COqt58RL7nd6YlyA5o4Bet0zM5ltBFVWKydZxuvCmo8V1ayuSzT64vndV2wFWFtJ
U9LbqUaAKqoXrp3x+Wf1cYOOVtFfWEYw7T8SlS6+di2ZUI1TpKPIpU5+pwdIW88emFacSDs4zgVX
3WxzdLGpIlp5rp2VL5MV49u8VMmlqUIr+uJ6D/uVh3mrMlo/aXbDTzn7bJqnC18RhT0ZwK07e3xZ
b0vt7pRknFCtgDfsfUeWpvBfUIwFjwWiGizqJ4gqw3FAlX6IvgAWgNVR5IK/+3NbOEfRmmkj6tpR
UVBtkXXhc8Yiwua2A8W2qPN6acXkbfLybXKx93zknn5evsucY1YhoPfHqttKX3YF7MLkt4kUL4HU
6Orzot2e7gniEQ9eRtS2K9Alwcrdp2fZ8O9RfFMZj4WzmpZ49nGazGpw5vICJh0dB4GcQTByFW8A
XEXl3SL/kcL2QpX0LTcLK7MwV0O4nnAXe0TnJo+VmO4zSFPQWNDlPGTEIJ2YckzwNXhbJklwz2O/
laVRHyocgrvmWKVdsPu215DhJnoPJs0dR1pxdaLsKEpogWLAee9hrA3tzAFPsMskyqtsBlox8LAs
53AYkya2O/NUV4Qlb8fzxfeceXbqLchDH3pOcWY/xzsR2uzM1HtHxi3iIVcLVItVLlfnKIqyhIes
N83xQMhBvHXrP8MCHt71yK5k+oEXeS2032YGxIl49MNi3/elRvL4aH4OIITWe/B1ZP9P+mzP9ePC
7h3u0o871BmMncfwgFQvItc0VK5p2k1ly1Kvb6p+dtm7aB2aK3rfePDUnsSwZCrmFzzF/oNSEdWu
5MnOLzfIf8EcdjjYVyR9ozBC4d830ug32ko7CQ6WS8xpOL/x1CXLmnHQIdd99tzQl6vIbEDYCQDu
bfdSydL5cjkKcG/kKZKfbGvP/Qf1J8fpPh1p7b3oenw/neCm5Kdn+mWAZltxXarBh7GUh+6rgwn0
TY/BdQ/wsPMzoCJQ4C5lulUsGjnDxQbPFasd5Bt8YLJvTMJppyIBeQQSIi5mO3Ok5sjD96vfuezU
iDsdYf6No9uLQu9PzgZIQ2VD6U4ghQdeqwzjddk/+KSh/3g5twzvdQ2SEu3riqjemaRwynnlQp+j
hiGcYWKERFTrWeNvllam1maiMTwwrCEZn0RaWjKSeielBl69Qd7an8Kgj6laIJbvQaiYbT+d+9Sm
lHpkiuGPT7q0JCIwCjr77XbLRZMWP/5xKaIk07RKHkqs2Zo55/pmq7ru2mOGauOfn4fHITN3q7ak
CExVrKiaUnkT19uWP0aBq+F6CK9j4vQOY/4Jc1GU8iR8QqOatuERhsrQh2ZKvnOPYDKzXg/lEBWQ
S/UggJriTp9LFP++YZysTvnepnJ366mrVC5ucr03yr0KrNcHtthKYlPfFenXKcTi8yQhA4HB6Vjp
tVLgDDaU43/Vpr4FuJrzGERQK1VykgkHQccJw2Nj/1NyCgobsz43kHPoNuwsRHDza5iLiqqajIFY
zQAjO0x/KVP1gBKD9D7ypNkm3hnappNhEcP/MlguCv7LWiSu7ZmfXXqbPL5BdaUwECeedf3GzbfW
j+LEpbRNg181t6Z69mk3c1j9TZcAVimapXq99+7xKbWEuirxWxHs/m0xvIYRGuX01wSqLgU7EGs8
1AvOsMKDlSf8rvRNJYj6+XPIHB+a6T68k14/8kku0ViXNSF18MWqrb4Jz12hG7lTicBB5rPZhDZD
2w3E0O+4odI6LN7bUHoYc5gdvP/HrUBqVfh8OA7BUjBnBnh4XetS7GKO7Aw5UKiuDeh+Nns37HFB
BldDni47RKMZ2LZmX4QXhszgEPrfplu7zQno0AXxde8I/CkhoUrTAEGKWOfyyK9+FApmWJ7NUpjL
Xj14EjgjzIHYTFn9QmyfDhF2xQ36VnKCgNRqVaeDHe/k/fizBxsIPD+4+IuPrE9v5gBe4EaphfZn
Ty/ShjCnBGSsRYN4l1BUMjPDEgvSKTpMjqaa191Y25JykzeoiECTX3xZ9Ra90T59QF7KmreD0VNl
Zgs+ji5NiYa3aqwxWYIhYrIYPKM1JuVHZTXcKT8NHWlcuibLcWAswyy2eHHp/pSK8er3roL6XOHd
TXWNuhnZPlqfDYk1Nm6RLVNcy+iHefgJHebj/dS8zl6LiEU8PN3sgXsuQGQayAM2/ozQugDwXAUL
6JIjkoyEdTllgM9qNaIDUHOwNVaK0mZNglplSlVdGRVtNXMsyS1trwxbDXVS5ooyq+7OGQitOyQb
xjA5WY9D/dM73lhDqwYBY+9EdXjpscRpHn0bdSiLfl/bzoaxeWxjk8j4NE4J4MHx2VMZDV7eX7nQ
Eaku3qqS0RXqZ/H8QZU/8SL8TiarPULwbuLua3w6B6OpulvBVXLRRDtObPPP8Fmfuyy7Tkn9O43p
iv3MQbQeFpr1h2+U6n6Vc7lfEONWepZGJ5g2xpabYAqf87njx5RDltJvan9l6B7yDi0BPkpXKzWv
xEkP1SBfCgZm90Z1CIgl9V18QEYi0CdcID7e8K0B4XbnKCs5zJppXUKTLxs4HCo/1FOD4flakAxY
RtcY4iYqaVOSe3DXod+d0OTd/en7vMkVNwyZcTX7opABbV6npWelKAY74z2zl7N+Sjn/aO2PoSRu
JtPB95dzbwaWMCWLA8q3A5gz+gDLViBWnwjAc6sDy7k588TXd/3neLuVlzMIFjCx0pzxKxFfASUG
7/tx6A+LpxbAl/ZvMtOEjPeRdl4+jQshPYeNxDzzbf8WMzbFvvA92aC1rgO3UMHBjU+nXx3D9YyR
WkZG+Mp5D+MwwVthmR7CL8SIYLZzGmUp35fBzELTwWAB91qvYKnPEyvTV4FVTm0pkobB5VNKCxzu
7HI4IoYUSAdgIxDXbig3JPxJ6JtIdxFSDB3PVPHYcE/BUz4+aipxwSILXn5FjK6uA58htfaaiweR
02b39p0+GsSqTLDqV5IJ26JA8lzAhPF0JvY9PUvzdLqbVpyE+gJcoxXxAbzXrcTdprKhQXwDLizt
wLSsDjRLV5XZZUxJaKQxCoi3G0KTP672MVowoD8RWMcS+yOgP/HSWNd9lF8ETP2sHpnfnpeLfcsc
VZlC7HK6XQOaJdiq2ceRj+GwBW7oXZ0wgLLQrUA/4u8y2ObA7Nnp95FnKtNEigJQvhSsui4kkpYM
5djbJlQTl8mCaP/eSdjSd8hglgxyEWeLqiGSHRw4NZtEGv/MX0NQgKGOaGycllC61dWqa4JsaXVL
AI+xY9kAtxqE4RaSfuYtmw8Z55a1gQsLi//4BVQgaukqjlioWTDFjVaAY5FcEn+C7zxHl7OHsccp
knWX0vio22VwSaixloJvxl+r+qm2Ic5g1pEN/ugsFBaJsm56Pjda1giyxH5XS7B7zUyKiPtZwwV4
di2pqCqO7ybHa+UGFtqnzS16GCJSd48UJQ/Asi6PirAmgukqaljDcs7u9GELFV2WiedEwn5RPfn8
3wE10TgQ+RHr3h0Mz7WWFUseLNqtNHRKvEURmCCU11Kn5d80dPQ4PAoLWGxXTXh/Uw/BVydze6wn
N4546ompneFKp50LAFm0hBVHtg60cbZPAx1+qpkZsTaLaS7K+cW6F40wCyt/MpXUmJbbEsIIG01U
sSlfu64l5Z9/Vhv5AxtKeP3RQNfbW9xuQfCuQAhuh+igMJxjR+CqRxDK87zJG267eY/MNYL1fg6H
rjL76HgZPvOmgd/pm7VvpuUjjLZdMgFPU1CcEWVNjEe/2SsqYDHVG4wYwioSfcGuG4lRi11ShYX+
ul5XAM/blQrTkYlGdIXhmc9CiAK7D5NA3sViuY5+/5VK0A9VmvDwRzdR8zA8iN9AFvu+X3U/5jXz
sMvL7LN2yBci8u07miea7fVxWcqTmuLiug8emADWcJZzI63/fupTeyCOBfeYNZC8VfojBlzKMz7V
neutub+mhJaZx391lQYAFgvsdBrPAKhLnl3ARmy+w49+othqgs6Yv8omPli3rUNBJRsw4zQMsrtG
mrkdczKvRFXH9cKrpQidLmkcnavESnsfOb5csOO4F6LKHEXW2v30BciO2E7xAX6asOi3OuPTKcDK
tB/FOeOOnmnQmrobJZS3tmjHJGCISL9svzloxx1oqOC7Ib1yzXgR81XPdGX03LnuVOkDwFJwEYxB
He/pvkxNOorRu7r4tPxgbcnxh3oifnLfzz1bXk9LTXXPiof/9ekCpLc/uLzdRz48EvrCFe0FGF48
Bw2SxBIDUDB5e8VxDBEkvtMgeUSigdJXaUpAGqLADnl7Qos+ZvMBcX/ae4a6c1x9euGs/u8SArUA
eh36FiqUg0/Hax2vK/bE5EX7rrlIcOabGFQ43Dr4CqylvWHQlnZS+d+pSJS1j/jYRSzARCImHFUI
Vmq3m7wy2HQ0fU1O5GIAoRzwlEmQvF3X5woLa0iNIvll2kh/Y96JgpooTBPIcveUP7ai+GjsTxI9
EVHLbvdF0go51Gid74aV8h7vJfoE5+wN8NCsY54mC07ck2TVp4BW52EC36sVfSaPP5YscBX4YqwJ
H4JZiHuU1AA55ginU2IFgQO1EbBZCoyLmEslrZZ+mh2B8upXThguzittNt4Pz8M1VoR5xEqakGl2
3YiaFCWN5xyQY4m64etdl8lvQ/cqMylv8GrniZ7vRAaTYraAfe89O5JyKPFHzVIjpQV35Qmi70AC
/3eo0texF8haAsKXinpb6HHVfzYC7Gy+te0pkUB94Iv88yv+qW4IEIuRX8StuUeXcYVYQWiovUT+
0tSV5wSEM4KqtnDIlvZRA9DY/WCUK690Sa9JIyJ4MpcoxShErs6Z5He734wTdNWcdUm5W1HzodWK
bNYrAn9uE2BsZq+VIwXKZygz+h4J7ylHLMAvwQJr++wTKhysukUlgfBjUEyi1qnGZY9e0q7XQgLm
FaLcEVcVFBw0Ngx42H2hch5h/yC4tC3V+KS853IKT2pJK+Rr+L6GwX3QGrgw1bwNTjqHk5KNOZMN
ZZTdnatonaUrDpk/7uRbinAsGYjQQ3/m3wIOIjXLhOMYZyzQXlmmToiPKjo4ZxUu7S9FbO5HSwR6
hODJryb3kwkHvfMfUvZRjm9b1mIcPtQ/XyDQz+Y8s5rpuP0vaQGg+npzusDB6RLgJ43DjpQCXpD0
sGwCgSn0EzK9w9Iah6tCbYhg7eGt2/HE48vktRv+dZqg+WI5XBSvZmFOU4Eh6u8IRBCkKIqsPxRE
kJgoNjatmtwpoY2DhGE7VMqZV6S7PV3Ly2plG6Dq+pgkRI5OA/0WVcWXhXYzqxE8GGLJgwMeFVAL
DijUc8lDAKAr6jlKZ8yfZt15PfhvyNGp76fjCzB4YsXXeJxhTk1j56erwmAGllSqR1iBym+7ORIy
RgqSpOIwEneKNOKUesJ+5q8PCpsyJG0wiFFl5xd4D4OqReUVz3Xwn0fvxmYULvB6PYGpoOQnTupA
FnHnDb1mT6wXvf+JYLZ5JN6cAD2+SGLqbsNH5HloQk+fRMh9PsbiR+CrV79AJkgpe4WU1RvVC1Zf
HX6DlpWqhsem7/xHiRe4mdWNfYvIBjeFaJCjQdjxtlH6tjpApmuLvFkL1bO82Ooq+amZvofulH7a
Q8plBVDAJFL5gJtLu8kaqiXDn7+RPa1qOwzdISNN4iwoTdqzgx3/aODd8xKzbjhifJVJ/0FjG0gM
eGi9p+wCPr5qpuFXKlPfxT+eU638ZPkSU+tyFr7fG+tQQsInBgAjrtyV06dv9w8qP7tXuuOqlb2Q
SzOPE5NLMXkTsDVxLvZG4BzmaWKg+e+FaUZRbqvjptQ1YDSgRcIXzmrdArb+Zz/LpvNKDPYQyDTQ
cp81lAvylghs4Ot7RfZUXFEYIApvMUk+K87SzCPRYvzALAJKQuKdHZ/b20TQ6cfzepRKpr3+oXAT
j+x3G2C2/oZAg7CJKDvEICmxd9KIxVai80wMFtSQLjzRcBy309zH6ZZLiKjBrgpSD5Z0Gp7fXCRb
YftqpPry+LpFHI7dyODJa9+TW4X3Wji3/BEmTARhk1rQO0Xwr4x8eOi4XpEjqLiBoFT3vOkGKTGy
jOFB8FYckj4a0z47fwaIuHlWihz1TZRl2jXztalR7kPXr3iG/hz69zvy1jVManmcd+HIDdvTdy6Y
u6DjdkOCQw39grlF6MywNllT8/ucVJymYjX1XgJpNZ8gkX11R0DV2CZ/T4hV5vlJhPV8eFeeEXmI
4PKSYCM+yJYs4BVcIomYmaPix03tBuoqP5b/GHXIRMt+BH2dGeGHgtyfOMcvnZP1O84TkcZ34WOB
/LOx9P13+d4e49MifyMVhgn5f7Ryf+34BsKJcSZLZ0l65mBOWdJ7/J+R59VVFTu2XUb8LUuK6nVt
LylnKTwpBlhMROt1DuMWmMJxgkJFY570lBbviqicIQJf6JyxZ8Kh7bWQNcIEzvwqVzVLxf23z/Q8
CYhGc4YO8epqe9v6KEWA0bYwPkCeeSJEcUy/b4VqLq0H0gj2lYpkeNNlUJ7IqI3f5tunC+ilcFjg
87riPh9gCZj2VeQ6tnu94dRor1OJbeupA6qYgh2rQbsyYrO6SrMYZpHRlQn4x9sm7Ex/pRUcmI6M
YDje/UrFTwvm0dSMf7VicCVluYktD547y1VZb2ziNzTB/MxdhstYTuLDwT9VS8O7V/GH6OZMdwJN
xUncadlSrvvHoBpEVPf54smhRMc9T75IFGkSc2HgGERguIVd6aL0ejYZK9V506iYaVXC9gdeqyed
Gj5Vmb2xE0ZQ2acz8Qllp6Fw9/7xUPmZc6cJEDkwAeawQTwmQH5+Pe5YLQspRSmhFGtcofsELCzs
zJeDP3BLN+tsbqt5gwEUHzOK2r7p7vAjCasCUK7n2Rqp1KB9WQqT+rJHeyzIHR9+xNV54ulQpyLB
+RgJRzNCWm0jWDHXf+xVm/aMT0CvlOhcpRkzXP7ywK2Jxc7pnMIQlvkIqEa+TgH3UB42WeS1RSMU
3jkkxDCD7ETymKTEFJ9qlA+QwxmM8XxU2RXPSp9dehJpQtv5zlOjn0cj7fcGsMEnoShvDXStg9ff
qxNobqjPBxijLu6ABhQP/0p/sZ95HEF39aPmdIpE8MdN/GWFy4Adjefltg4vt6p/TcTt90JT3sMq
2ikv3+l9lYS7kzP7+UMi/G8//qSbw3BP9Sf/Aq00eCZ+Q2kERRci+VxLJn8zMC4ppJrQbeekFm1T
EjTG7AtKTECPYtdHeKxnWBHN/gMIyPkWKLmQPmlC9grUaq+rVGg7OvpedYQK8rY5cWy62gxkfRMb
cVlFStdfpxRENpNu3MKm87fG/wHtmOHk4UhPGqrLyMXS/EG2ocKHyiAsaspw7vzXTm8Woh5MXmok
Y6KIp5aFsoggDJs1jctA0mgR6oyxdq/eNktlj0JqREcVvpQXB2x53cgjSYM0a+8Qb5eXaOMqSBXS
NDvUWw3ZUVEG++yJt5X7WNW9Z/6V4FoN1I5+lixKOgSnz6Z6iXsz2o/Rbk3ytsHKfgoydOjOr1rP
xAIv7cEiMcYkRw8jVaXu73xGamqlfSSKczlGPD+8mlaqMFsLhuYgEJCLEm5mPx9ecq7WH+oTaS8x
fV00dPvDxR/3E2Czjkm9jNBwxI0/DhNlI+rWWMbMtPwkmR+awuB6OrTiLDoZMRYwJ2DeU6pkoEMt
5uVc92tiFT2ORZqrxT/cf/35ibdOxehkM+P2P+k1oAezJ8Kp8B2NeNA8MPXQ9LdzEAouUgbxKdkK
9Gis/njH3usVphn1HGCBKrRWUhqdo/hLyNLSclfsGfMFTDHCqUo+P3zZnOJeKSNLWZ8GIN+Cuh3S
FlKuO3rNC3Amr19G6lZVIb/CtxdPpdDdjg4nyUJg3pmcAb14HozHnUAPuE+wCj9w9w7pIoi6PD+F
axklTB0BfN50CLgWufT0IPRaOP7RJbRHcCsRTxnRZHp6JTe6kvvtd0Zz+Z4+i4GMyIeOwmd63vg7
FQe7TcnJdvTz1+DmVArasn3RgrHfOYnQs4KgZgtnuMXvktHWDNhQwz9cttOsFp1vMD+lPpk6lXKO
KA6N6Lni6u2VKu+ZGMkZ+Sxk/3YNLQigoHeivcBfz349ZD886NZHXYRz/7sriKTCcrO7/gm77Qef
78RZKtMeH3Z1leLAVg4pBkAuJABslytQa8gSFRBcZLcs4WYtTD6vEcKQIIp8O42IeTTiHxrUWfBA
4ff9jGGQuU4MUQnMDXd+5A/3yNh0ZWmNQ/KcwH7QVzgCAaxya0DZjsjSeRbY9kzXSo4nnKJxTd6h
ovBvK4jhVcHmdk7NevCwD7i+UKhEehG583uSOXEiosQE5ahxDOSngYoaX8pyw6LrxAdSJI/JVTbF
EfMLR8sExG/J6iOseyxDkqxSTOa/hA+7y2FjHKzxCBUoOY5S0NFKcXEfpTsYuhvRx7Cn8lziMyTN
Nz9YRNKj/RSyfkBUDH4r8LGV2PsdJh1Xu/sTEKsXYCqtK+kt8KXk+FpkD12Munm4yCGwrT8FT19R
jb3IikOYoVogEho81BFvJ3EVF0QJZ8qEJrIOvQb5cKRlA2HXLf/SOVzKIJzlVpvnhIOcP3KBZMdA
apvZRp3eT2EWlGbXHvVAGWoj67E7UnmjNDzcGBZQDaEwVUiiXeAa5lNR6ZsCwi+RiUx0KD2KrHoo
7DViXEje5uEmdBn+lPnB9n5WAtwyXBzYyzVGndA9Nr1bwF90jgzp0gD/B1E8eqQt4kpykqmk0dpz
Wa4RPNKtQuNwqy9SdWqLWTSwkfHbsITa/mKGIQtIqKmkVPyppVBw7WCHgEkb8qToBk1GdjijYFtS
H9zydRCEUqwU10zvEGzDqETzF+7zvTrcRgjhVn9AyPK6ekUjcfE1oQO33boJzSiNlTggZv3W6ul8
ORyTz+DOw2XXu8uve/z9v1hSYpwy0ssk3o083CGHN8O8wJYepMtzGMEKLWhK7tLZHl39Vs0s3cvd
mBBs2drT3qlxRDBNIsvitqsGOwGMuZU1NfW6LMGxuE83g723worLZ4/NixG8LwHHgjODMlkMGtru
PwvEnWG2RuiRrpqGCF/qYEfPIoHcPStkqmGGrks3EWprCOMiI9E34oVUxn+Effrc150eXsYpOyLk
Oiy0Ndnfgw61GiTFo92ObXLh9djniQM8cmw47zOS/rmFGOAuFU1/iNib1A7ZjGOM0Airxzenu70s
u7pCmTm/rRLjWryLZK/+aG7CVIwfJ6XcAVSlLQ+DIA5mI/em02wjlfOY/h4ADFe4BlfgTqf+hPoh
/nPbOygLc8EIBOtl36hr8dqCcSNd5S2MsO947faGDEk3q+SmNFBjv4Qv+o8wnzCaCbvyCIBpuVwf
cLgX/HmYlm5M6z0qxjhH7Z/Oav3twPh0tKmOm+Kt3Oe4AyAWJ34YhVgu1W90xuBjgkoh1lFK1ZPg
82/+UPNi6YrvaeOeTiBS81ZyWec9N9dWOH5q+KlXd+ACPXdrfoP9DYyjjUWvwg0xqGxtu4Lp/PO7
RpcVfWg+80VtH1r0WCjh+F8Wm2m/+rZP4Fzgytp1/nqwvP10t+5Yn9S0xH9vUIMF4YcaEXstOh62
Vr6qSG62z/Xp1emUgl+iQ//nqyMFiGNWbQM3rzW4LP0uO44dG6ZJmHXJOpCBz0qB2pjP5DHYMWMi
03KU0WqwaTD7n20XkgZ8OYt5x+oKQOgvkeMQ2X175R3nfXVnrPpxL/P9ZN1ZE5UIE4pxKxJ4HgNo
8jB+s6YuWnwXhiMheXygRTChBGA3Ew3AeVF4FSR4uJxHSGTheG1rQQETK5lup+KSdWbyGFxYcxNf
IGSTXSY5IcXQWa+16kQl9WevlZEQIiH+22ifdpDedIz0VWjiRVtzSZA7NWDEml2duOJoBfG+iOCP
aSmEz5OnILT2br09xE1ZcbcI/YOhz4NDPiqfvUTiPQ207AXaA96TFWnPA7f1cVygkLun4NOx4gPf
UYMQ59H9l3H266xEKfwPSF5EecqbxqgwyPA1utEYQP6PkjD1jLUptdTtWC5xn67omz9S4wusioU6
D5BcnFDJU+mNfUqIUml1JpGB6bBJCe373B7orHLqR8W56MiS0+AG7IpZAky0OnBgVeO6NaPLIu5I
vxzN7mKKYyavMkto78h3wdTUGiwkK0CHanDp3LtXSDsZas01/egNlNqpq5mXnzXLAXrOFO7P2KTY
Nw10sPvErcue6z0M0jRAq8uhw5IRA8RClYswDAJuxZhCmIOanwMsp4+fJwOe5HBZoRu1mBiQrGXY
Dcn2jSrAHZw/qh5/twpXMph4AqjLZzdOR474rkOh/VGHCZftho53Bu062YTb7ciRq/YNf1ry9c+n
MoTU6urrLtMihtQVoExeoYrnwe1/sCQ7MYzsfoMjNAX2Du0+1gGF87tiFqOMkUtKiNsOKLFLIV8K
EoU+D4FpwzESlAVe0pJYKhDss+RuUvk85GeX6Zt0LEr60j4ize676LtDNdsyhPPMDzE8ForTOpWv
JLxnJHK6ovvIsZ3m4DcBwomD5/1QBTaYMtKAEuE7RRw4ripjXtow40OE9pAHcsBIwZl0/4yFXeqM
93rUQbx8DpGtzSJZVekUhqz2Yqc1B0OILUsIOfj2tIdJUCa3Cv761dwa+LJNdPf8+Lh4CbA1Gl9r
+vmFlKqSoiA5M54EPuf7Bzdb2zemBkrMrk19CJFqMLPDuDj1dIovOZr831qiPxyzpzc2gwnPLQp3
JUOw121OnCV6LudRSkStOLA3ECZ2yD3kcewIhd9ooBqtPJeDns5BK6tf3ugEfY06pzHEt4h5pabD
uS29HtkFfw+Eipywr3ndFIjfHnsLPSHcaO4fmy/UPqPhdOsUSmne/G2Atsf4UHM7eXHhU11MsPtf
0naVglx/OzoHjCSt/ikMFcWsVQ3AO3opE1jaJV2sNccRYO1couQpZnErh2JqiFTZcyr52ivVPOTt
e6aWutPwTKzZZtJdJlk8DXX8aRf1gt0u/pisEdXVhq3m4LFE7cLVIVTMmjVhvx4vXZ6ujmsO9SOd
pHhYUuSSn2GY1R4ducDqzTeJD65YgjRpOv8+ofAIP4icNt0dIjIAxmmTsIMQ/GFsRJP0sHUwwudK
0xnmB7aEJn3uqIOzK8RsqxstZW936RzltAsONNaGGJfJRPgb68EKf7WqXyMQcg4kDAPva0oSczAy
XhKSI/udywhm6egv/kPDRfixcCuwzgTmolZm66db15nfrS5G+NZ86DU9PfK02Uu77f+0+8SRMRTl
DFv6Icdrgd0Z0TXgfJM/CsrRmULD3HFztBxzUZuo+KTuPYn8QBXJWy8kIWVl3112ppXQvHon27B1
boxytX2xTxkpc1CT/FKtYhClbm9CWIoO6hMALXjZ+7l9B41YoHb4LpKL++54LOIsHIALC1Hc128w
cU4k8dupX31G2mvV2i8F+vMgEsomcqMcYa41n04oxEX/SM2Kvi8BBRREVWHVO3QvX2YEzYk6NJP6
STn+QM8eAdGWpPrbmWfsayml9KL/gBJ0WvOKoH7G9oanbQf5QVgXqedrED/aQvJKY1HbgPblGWJd
36vwWcHI4Gnav/vbIL6I2PZTHxZFVzaKz6ZJbUnBT9vHk4yadMnpDwuNH4Xb9bfu42csPTuzjSHo
Ef37XiDlTSUY81k7a1BIO0ruFPpr12nl7MrFNwhieDMDsamYpxLZW+93XkXgm8sX0dvYf2BGXm2C
lnTY+MuWkPZf+m/62itODxrozQ613WpphTwJfnqfcGVuKG9NfuKCpETf4Y3tuDKy7hhF1JcIKHEJ
Qiey2A0R4y4eS7mM2momX6dXOL54oPknVDXSaLGnVVEcbBzpt72YGZ1C6qIj/UkpIQxqn5roS8LR
J8m6YsCRkcoLAXM2vkwGgRZOWSDL6miqUDN2CZSnlqztpysVBPsCeG+f0g9kqITDqXFz9aEWdVme
tnqRr4SBlRp//wPPQcZfemavToBK2X+5sC/VWT8aWb5ni2G+tnIIQiuBYqh4FgSdDecigPK6sCv5
fU+I/Q84OG1qqfI1/uq0iKJNbWHWm7Zt8/mD1HRZXjwTrXrqEmO2F8qALA9/cqQ0FMSxBWckAoA2
/rDvXbvbfdbqqZxx7CbdH/acBRvtS8srD9r6Nb9Jhf8w1icaNBxoG1T0y4UdHyCmwO+PsbqGMXP3
X1FJmq7Hj/s8bxaruc8sVXXtcyHI9DbLgWvOX+1+JpkvHPRKsH76vYzMtytLpEZRotYWRYhCM21B
6MRIBZMOmxS5rF40VxS/4zU1x2KzQXkeUrcFoCm+BMlDuggZhaoGZoadEXi+FSnpyp3z8/yFPjfx
b8lSQXA9Y4n3xvXI8MStIumM9yb9VxO8WC70xKmMlCXTsKn9awrlKC5r4mFl4bs3lsXxMtxhSdD8
nmD0HL2Q8+bh08E5QwW6tLBRr9TzoKzp7S83CPqNwn0TasJPk0+WmOXk58Fr2PL1Rg0ir451sH5g
JsgJ05YCklAXWEVjsbfUf2GZUgKsyyto15mavzCpV18//jFjtq/Kldyp15vckYVvxi/BgoFTVtAl
atS3TX3InPeoMDTFZJXhsGQ4Whuv/vx0yDEp02oIsJr4O5MMP6VWlxzvjlbM0tm12fK0iMXZ4q+j
WTxVeZGM6umfLsZ/nQoeWdW9x59IxjZLbuNFxdja6riFJ59ftvoLKyjUNCz2x7Rk0qVPg9eJTrF0
cb4ftADEeTmz/rbCGgC/aCLFGxOoriJHsQNs/KsDtWz7q5G1LrcffN5dagM9fCg8WtRLJZQGFON5
HzmU/QOhuT5Z2JSZi8MdUa9zRsL/liVvvXnQ9d+1J3pleCtQT2URtNtkWqPcWGKZD2pBRPc6t6j8
SfRuMe+qug7Lu/dPsufWLBix3w3HkupTyPojehUFUvA9YtJ+D25FQN9/c3JfuehJgMpGjQ5IUCpS
n4OaGoRY02hhaknfpjUCVB9qrjxNiLc8F8HKqE0MBaAgkT353OM5Boe7zX/1E4ai1sZY/0BWEwGe
l8BtVzGN6Y8HRpDGuv7dgMbVmD+PxpowUv6m2d2MOjl9FDpfQY79zIvMG4XATgfC02AjZ5JU365k
m0U1XGS3sdQC1U6HY2kohwxkNP2oQFF0CohRoyAVTUf/dC3yBxeS3H1LnSVitjwCLs9UQhTxX1tn
6/MCq3kib5lt/ky9tFghLjfv/gQVAXEPZ7kkqi84hx+MPbpZoG5Zb8vu91SRagFsP1NsRVZaE9M1
E34icFOWYxvIFPPBVOd6Mmt0oYvajWBpAM5sPaVOpHmTUxeXGoKB432lfmN5VjLlyT9wjWIzpwV/
oVtQRKjwr+jc8cjYk0jcTVA98nY2YZKuFnQGjt7vMjpLJrCRdp3EYLKr2sxkPqXGF7XoFqW/nrWT
sx0ZWMbQKhtoggGynhOqdCLbqQYtywStrQMqqyN1DdUQvPb/kmUV0sK5Y9nBcec+YR7nsJKKzYfD
m3rCBvYejK3U7GIjnnI8KEU9T+JGq4SYg48u4bx6D5t+qwVPeRyvNt1h1PMGDEL0sGankHOGPlNN
fTb9M1MlTB+BVcc0HPbAIzWPXCfsMdEdGcj53bS1UED5UHGaeUU2iBNIyUu4rK4EzQ0UdgwpW0Sy
bFiyJnsgK/W8ErwgM/Gc7o3J4FYGgwmj8VagmFPD3PKS4GLYad3U3CUcnwGwgGFJ7ExkgVBzxGvM
5pvHmEF3dgb4TS+N5tWSEOGkJVSAMKzbHB2ciQb873kkSiNBIwW1UstGiZ1wW6IfdQ/Hal0t2S/T
UdDQCQ7++BJ5wKLJkiluskV6BFi0z4v6YJyZD6XPaCNF0Cb3xG9aq8KQE0rAlk3PisLuHOVVvOhq
I2Y8BBYmuJXmZzzN0M5GY+opaBwTOZulf0ELpNLU6DQIhbq+o3blbfx0F6Sbi7Zj6fmJLuD2HL37
3E/WGI8l0rimAVK+9ORyWphtp9hFriL07aRMvTLld9M/fAohj1x6ZwyGM+BDhHM9irzR+6x905kR
C4qnHPvrF1LL1txLcFbnp7yQqqEH7uHKZaBbazI2NPECh9QfM2q5xSAjattTGFvXe85d/sI9oO7S
Gnq4iVq37dn25S6Yvrbc2sNJL3/dBUBrZttwafpgc3tc2QmgsJhsp3Bwn+ZCUmmgmZPvX9WDnKH9
0237fy7/R2DS2VwJY4yUgrLNqHlgHlQPTSTyimx9oV0UuSLG6+n/FBUjixtOTh0JG8OIKJVs5XDv
syOsNwqlzN1QDVwGCIivHXiTp4mNLSXDcOSpc0ZVqZ8DUFVmqfjf8SuiAzaxKYH+1JqYUCGzHt8u
PakGOHzbPzUMznt+TRmY+gqpHo2n1LGPP03kb/OPo/xvMWz9LT2sxZ2uidnTwEmJ4wUNkR3WlIjH
FwyBpPaGRpu56clJP3Zu3AuDhR2iotTFCiZxSW+xjslggdPeTHHIphcv2vhE3RIzr9hK/NC0kJb3
QPsHWaf5G8F4mKWpkHQaxNWGgnH8Ek1/L5ynofWTX/LabepbT5U73llq4IeLxCW7Gy08Wx60ILXV
ie7IoLxjgJ6FpjB5XTLNnD+R2IeWEMLeisVpaREqPYqzIOPiPFeM4NRLlHGQqICiNCO5jnEUQhVu
zARD7R6Fth+jyM4SMORlVfXressJyKIvq+bdYZFHeeJpQwi5KRoJGzD3xHANBcvWOncTRWmcRs7m
ZHpBQMeOC+PJcl670SsAAEEQvJnIPoCqgDBPUJaPLvMiLy2k255fVSDvzudcWI4iRi/NXKDU7qf8
Xo5gZHWF4DBh2xxBuYlfxOPlXXyoKT/ZU7FhsZ3JmsGbgUwEBQ3KvnqfZWOZEbEC+t6Fs4zdk6Oh
tXUYqgnFQFKzszLFvg6pyF6NGKELE6DMssNs9bWlLImWarks8hVFhbuTPw6//7vOhzjUHUrE+tnT
jjAls8aYmkc++nhiWMK8h+ySmUZdqmtKQ2MmMerqtSS+N7b/FHoybdSgUsO1z0Ga8xlwtJj6slKT
o1AwsHaTkySjDzFJ4tfZ08OXvKqzAQfXzSF9OpcgTbd+Vd+mDvki/uG8OiYT0djZdz9X8mKO4AR/
IsEhhAIiZVitCXZiyhSSFG9R19odLh71vyPJz/XSvAULyswaCgMWj6ZQZY88oavQA7pU+kEuwZO4
EPtcvZTpSatt7rBnwDfl0DclOoCVDwTFNVNTOl2muqOBGWkOGlz2CIoWtqt09LJYfzbv7CjwlF68
OkapSQO0cplPdELq3o8RHNJAmzNheE+Hg+0XGaazs6Q97HVufGHmVmgAqa2R0c94HyfherMuo/m6
d/jKdD1Ppwda2fLG3YaN1aaGj6BIIG2ulZaYaKNKsUhFW8F5QKteCmfK+IySZza6pICB71rD9jDI
6zKHJZRZxvChHzzULsFoPzK9C6+pn4UXVw/M44u+G/IwpPeNEUZVwmFMbK0zVw63b8aJ5yFy9bYa
CZWu9k4BSElbq4HEsPMsNu4j1UMK1HamxCJrrx84M2TVjq28FwBh2qtB1Td/SDBHvr/wLRzul2Qv
T+GcOuky/hVqelZqubtw8uY+2C7X/5B10y8vMqFxiZw6rZDiQDCK70LP9SF8FQHE83U5/R9e8+29
CRK4UlONC3DTlOqZ2eq7E/fj49cLppbF/9R9Rb9WHNkPeCRLLahKQJMtVj+EQmBlG+yV8Z5vldpS
/c9z2P0l03iy7tlMx5e7ByHbqJ6ImfLkCZorKrqWQ0eP7oCGzf7wwJ8jwjtkvzXWeMCeqn7phu0f
3gaqaAfbFKkTw3Gy8slvsgKTbnbfTXfCgeVSWtIb6XLY7TIFIu/SC10jIQUCNeD3LCnuaCqq74gz
NL6VqBnz3KpkaYgfgW7sb13735ivKhgYx5ldrVuz3/F3bWYMXmFVbD+ADbU5twPj++GD9foRSMU0
CKfXfOPsvFJcT7Lz3JQWwcwV9rLsDyip9J1vJWqBJBka8tfeN+GL+OGLxnJmiv5RaT6FG6QADSoD
DXonj6PB9EaveRvqMByRokKFkIN6OE3G1TlbcY9nwT5ku55Rk/F6hKe62JIVESiDlaOVk1PVkShc
AruyXMDR3ocgFS2evxJWaej3l+SHdxu5NG7WsHj/R7L0wZ3jBWvLkY1kfuF2+fJinCWfQw7CQiqr
b4rosG8e/qU4eJNapJsF8hjZYB0ALSReDHVjeq+I117fKZgfGZXZvTrx+98ALWNm4rrneg3/PdS1
DWrfB4xRcEntI4m373lXHKXPagCQ/Jap0Swdp5SHLlxpyXQD+uw2uGEoDFAF3IfsKqE/3DTY3J2Q
IelBlkO4p9jT2zZm92CcAsdqWZ5IXLLLnZDHABsrYmfx3hp+sVMyH/5VFhjEPSA9z8RCaBR0bkzD
G5H+9gS8pKUNvQfUUm5z57w/k5f2rP86sCmFBMunijjUnPjd8qdlBhzFy3ujRR554HHGgCbOeFuT
iG2+gprGAMMxhR0rBNdYAfnjJfCzTsFc4NkKdDcNSY7b6rNZBrYCn5808W6A1Gb6YfNYWzvm3BKL
PX89RXPEJGnMGv7CdjUTq6HYijIL6wN+lJZND0YN6PoBgyH1mK1e6s4y9ceYcri6LlT5+4mBYrxM
vLqXK6HFZq4uSeE7Avu2VGYkzbdfJQjH0q7iZPdR+BT4sZYC7L+2FIdDs/uTcRNEwVLyb9F07CBS
D6/d283lWxK7Q/2F1s8IVzQtM1IGUbPNcWDHJoZQ6ihSt8sILOahYqVHG7avOo/Dp9b4WkAZnVWk
IZwWhMLKA6UYaba6Gn5NnqyCwiLdJcQsTInmqC24amMV1oJC7gT5oy5OnxJxEsehbSqzwvj+oOL4
Fp3OOKfyASWhkGdRRbXLx7gTmuiWT+Noz9LplqXk+q96vM6jPaVf1tOrrsleZ1zSoyFiiMTFRi8W
GViD1qbaUL12OLf2Bip/wVd4pCH/REVOg/qFleOtNq/RAbZmS4tdNihBdb5klA/cdF3onq78iNTI
tV4hx3WNfdTFb2i1Yp5TbMOeZwV9a/icLyroJs9odPi4LlG63aRtVIpo0MHQMWZloEvLE3WnHhPI
mAcq1FrypBn7NfR2+Gqmki05pZrPtvJyUB3KJyolJZMyiu4V+OEGP8LYNwhJ9pr3+aydtB2gtMjw
ow3yO0RXvt1tGwTXSnYMpItk4akbHViJwaAR6DeCp7Yp024OILJ8veiISrFb9VwXupnMNswpWRmT
kYTRKtZ2aiHuSruvDEGNwgjtg0U2zYReYuTPMt8yRr3hUl2yOJPlZTudljIIIRgzQN681WoEcscr
6GYbDUrnN11R1pJRjBe/C5hZGvDXFPXgA0ujJBUZBR48PU+SINj6t/4crxX2a0ou/MveaATbphiF
CRDivODOwCHF6hEstJbPeHqTFhEv4UstitibBrU+YQd+jg9DlcOkGDnBWzfNB+pC9IdNOx0O6tHE
SxVnidntNXN135iCxncVxY4PaJHxeqPN0y6kaljfzg99CKrJRUMd0Jz+UOv4uR7GcTYFBfSL9+nx
dTL0WUnZHN+Y94U/ctvAay01SrasANTfxxPpKL4FWYk3wP2TbqiNARGdKIqmMeLzVf/LejLQgHcm
OszAs4hyuKElRr+B51u0JKL34+sPOiP0MqiU6HqlTWkQMF4ENVSqS1U83MaBn5Ti0eWa1s9BQwJq
aMKyYVe32AALUu5ooNVgZwJTRcyfzPqp8u3DnoMqPce4GEK8n+cuJsSU0wSgb1eKzX6ycnLm0CFt
02MsO6WNv3Fr5yQh8EpJvEHaOESXuSxKlciqw1RZzn6//dsInL7BZwzQDlgzlHwv0Yglp17NyuPq
Owf8WHUYF8KAdzEjsrTI9o4YyWUEPkpwxiOnuShRQkZ1va4NerwmUXmWM02NZ1VsZjVFCVuZ+vw/
0liVAd7QaMBc1AJYMwFVKuqkwm29p/tDIQW6x/EG9K3RNR/TcAK7vXomm+uRmi1GVDoh7q/K5BXS
69Vt72yeOtARhmwYDT6YOge4r9UAf4wPAQEQaAFt7iOuVpUJkaHtfkO7oKv4/E9u2/8bMyt4cwCR
6g31IvD/gIvNTer2mr9XI8fpLMh35+yf1QOP/afCCptRoIcvqBeAH219UCfV/gq1mH20cWTEiHt2
M7/NfcB5gSn6vAydjV0Mb+MX+gnVurZCMMqodVHhPw/NogDGWt/JTuP+cW65iGf68Ojgvje6m82B
ZtMo76SWK8pbWY6A0flpIOotHtzwqRg1cZ2KIXuPlq2lJHXrGCQiiQDBgstOFd5x4oHS3P0BZYCb
B7YFaIE9swzc8V9SzzTjfSO1IxwjlnEyCcvX1hHDwbhu94LWeAkVFkRDOu7UiJjbxq+YLF6rz+Pi
KiR1R0aUMgFWrqF8IIrUFK3StCHuyGYtNg+tfi51NPuz3pDCXxnGW+f+XWCLPsRP93+AiEHUee8a
T3xxNvtjlza0jy0jULrc2uNPVxNlmTlbQQEzU8xJ8CREVMdZ72FD6iQ2UsBtf3jmSJKDDU8pXFJT
Egf9GWxXi8zfYjmOrdNz6Eo4fJrtj0fR4cT/tr/YOH+VFedSnhEDLcPTCXfz/q2cgcOlLjQiDQls
al/lr0k9ZOXjvX+uNK/5AwFkUHUuJxVLoT4KbXXkY00b60vna61HsTiD4VtwhwtYNwvKzY3f7BHy
bXPDFh1mxhufHS2nx98/zyXEDRQ7O/wjk0HQT+6GQ/gN0UCe/gRV6+ndKWDjM4WsTs8sT+3d0tkS
+cl92U5g3Pk6YM5Idj4Srs0e4d5Up0RWoH4dZH3HR2zFvbiZXupAakjssMTfoMaX5RsXdEXXdp/A
nRLqOPLekDXa9YJwvqEYQaTMA/m9fbHREWbPJ6nZBC+LQ//jqPiHhkGH1/LuH40Nb+wkV8tB9xlo
xLAPO3attAqNi67JHE4AEXJpJIoGMWN7cFHaPV84FoUT7wSFi+UjT9Ejs4CJVJequMWOIHBl3PAg
YlpLl07D6jwbuEa3tpjX1MUKLVYOs6fXb0EFP3RkvfywPuU5vSAebYYk40nJkNVLYxXpsc5sHmRu
44/T90AaleaDhUVHGuajF9lJ97FUHBe/gf5q2QhYJbmQfggl1QuEapMhjKRY2ks12YCoFgzW1oB8
JiM0EAfG1qewAdT1F4uiHnr5D8aX0vQ/+dWe7psyuPGjdecgntuTZy0B81mSs2upONC7ChHHSmVG
oAh09yaTJVwpMWpT+EKYSbsZ4PQxPH+A+dpiwosLrKZklIPG33oR6lYHs+U4h7nbwduvWLesnA1m
Y6zH/8V9B7+GNnIkQQhXwW10jmVcy9HtFf24+tc0sZ27eZ5qva4E9+JvfMwbZ9nX3p/kXLy7aRNX
i4jdWh+e28AlK1FKk5WDRBlkRT4SeS16v/omTQNlE7k7nLxsr1YkyrnG6Rz33vPrB0eUfjdFp5xP
rMv4FfAFUXBUgHL2dfKzKwSVNXdA3LC8aUHsU6eherkjAZcw+zyNr6qNlo2PmvZq+uJYgBheU0Qi
YC4W1iW7jzoEVjdvV8RHKBJcpn2cE4Lt7CENkxAy+TZgrRNryvVHKgXS2AkU8esSAs5CX0pnlGJH
Zr1TdtOUTjAlI7dRmcC+oBXtXMotNgYSjwk6whdXppaS6xDd8bzF2DPYN7xtVLSMPIfPiOega9Ba
5B6Xl8NrtBr80Y3Hv1p6Hea07x6X65DM4atK/HWlnrg8ZjKHg1TlDPVvIU08n4aM+qfRYUz9ASp+
4bCjFbwRzmVi5vsMa0WDay2NAD95tScFKXnz/yl79+Isk5GcFXW33CO5Ejxd+szyTstI16c77uig
Qv2+TIE+mG1YRYae2kqsDpLbeKxdxqdiTX3Blp7pyB1+hvLoX90sKx9CGVuw2C3f+r5cRQzOwDDL
Rl/+KJJvkEM5e9LNbxHiedhwz1MMm+bwBLzzdUNUUjexjQEcF1K1xaZ8cQ09+5aPjwdudJ+dpSRu
uqjgtOI0Ki/PkZrWrTnEfI1fnXJSqVw7ZaEYHoHX8oY4fLXjhAFKQR7z3Uv/D/OZJ4u2uZd4C/XV
uRASj0ZFhKhll/XzBfF1FCRRwk/cLS3H5TDAplaS5f3shauilLOisUk10EMBal0D4c+qlMQE3XSU
8mAADaAUN8WJ+Ok7fdRMKWWbVI4gKDBpxXpK65mqFIR0uxBn4CMFvxBQgVgmiikWN7JymyD3JQDj
ThaYVuXgQFEyquQnSVIh11Wl0lKnlCPfiLOtxJ2Mug7YykwjQvEngNHD+RG6ZDGiF3ftPO3QkF9P
OZikk0ek81WVYqibuopQGHG34nSlMD+pidLhpumaGgQWUsXJeFmyxtdzhkhDLPbddsMImdFW7QlI
LQWoa9IStWqq9SjrJx8Jtj5OWjrCZc4xiA/kJTvNBIkei+hlPM+PoqhPim9HhW2NQkD+A5FdWRH9
ka6JcXa3fe5olYkAfHE3CbA5wMgWj+SJYHpbjWKcLnyohTDcBvnKc7Pid73wv31P0fCIqMvZEU1B
s/+QGhATS+NkwKl58l82/kxD5OwdhjbVZDCwqs75OOGadieVHYgyxBUeXqnsr03wFzx4lskBeJ76
oTl5d7QHdJH5x+qzyW78iPsnulvKZoW+Ial+iSabCgTF4WZZjrX1eff56J1j9f3HB6SjYirTd41s
vaP6VBPG2pXfZbVGNo1rk7N0VlbJTXBcO1rDY0rrApyxuwLib2tOZyi2O4Yr+cyJeTMtQJY2i5lq
Wz7wVGjeabOrqzR91FAoI/tmYMTDqikYRaJif2OxCeG49fx02LbbivW+/qy6Ikf6cho8ND7ITNEd
ersA7Ivgc9fbxWhARi+GIRieXjQ73JGSoCyT1aC+yIB1/+s0f584gmXd2cXW7Ks86dDGOIPPz5IH
+RXMWLG1OliSYTwCN8p9vMIlf369+Ip+gdtCOZt5Kqq+UagsJMqgz4rnSkT/meD2pN9Rg/OILpmj
bW8Q+3J4ANHDmtuQZo6u/qCOXNvltfXXvLQdKfgjhQ2swc4GyuBk014nUbE2mYPCAVS8SS87RHTP
dG0uS6Gw6Sr7LEvesOq1TMQAyO/y3rIr1sy5sZ7WEw4bR4XkPYIE1SkwQTgXFfJU7GeWuoRfvjDb
MppNXNgQ42bmiaipCQBRLERewkZOQjKsG+ocowQTPVLFdosZ9WedSFm5k4P59cjGugxx+3uHEsVr
yJpCuKLI8mhFPeASFaVmgB+5QpS+V289DPi6pw5UI/t1bna03ZRy8iGf6HZhmLXe2uaN6LTmW+bz
X+wPiVwWhjU/MXUHOAK5D7AaK/05bhfOev738bj2h6aoi9hBaZt+ULxWjnWKg2j7OwylLYSHUAAb
kDiWAzrXF0T+YF559P6kk9LNbLP2cVAm6DQXaPc4DEuHj96FgWgyVoxUXBNocENlDFDe3Rs2A+pQ
0CsTBie/5qIlnnJy+bdlyO9ncc9JLx1tkCh4CfERCjCVGXK77FpVhxtBbjt83j5zuIPCBwNTiU3o
45vo0qS3453ljPSqd32Cx8JFsmkaQ5yAD9EDprwsezDYnEAIXGisp1u6EWGYy303J5X8S3jhaKRl
513Ro2o9+Gx/8Z3tR3Nvi6WJkIM1HmRv5jer1t2f1tT2ZUVG1GEaVEIurGExg/MRbjORSATagGyl
pubaEUSZhqBVEOwwT45UvMMh1QVFDVXvnfoLe3UHyCBYRdAxsoLEKp84DJAr/6YQ6g8Xp2uDOuC/
ctUxLsVtqdugEDzdTBiaQDv0vT4T2CgqOmIqmY6uTAxMGs7Y255bVMxPH/Nuvb65jYON6RPD4U6i
PGCtuWI35MEzUMZqryeFwYWYxculYNDVwSHwHx0LRp0F+/klUh60iOt3j/dzBVa1x7k/7pU2MtOt
do5JZ0TnMQkQC8atUOrWlQoueLN7QQsu/41JGYRtEP7N89wZIJzN8t7Re17VQEgtMX76TaTVJwB9
ZvQ9AiUR9eNTMDHWzGB5O/8fcBnvcE0CnYMJh7+B6Tlug3erFFCMXpxPYt5CicmZ+FA7HAkATeUP
Obl13C5QozkKOCmJZoSa+bqB/RaEeXyDbr8ird5zAZo31Du0qfNHCUIv+eSPKbZp6leR14PYiaX0
gaJDDYz1gTsQJud0DqRwY/mRU/l3sZ9Xy1Qo6Q+phxfRGQ2oxbUnKXTjRlPmTGnwfhn1Ij2uOe9G
XzEPVKAgFaIpElEHLeWb0KjCmUcPTfKXH9RtPqXh5k1NnFt3S41WfGxJere/vvLTQ0sHos7kiYnw
lHYXc/lVK/91vXQVe3RlqB0bgwWo7iF//h7AGV4lUx4osvV5suzLUolFqXHFpY1ErgALpGoLFyFn
peTuF69qscFKH+fWw3iDsYhIClx4dwj2WW4SNk/bXgxD696PT1MxbxAxgnxVOKJw4QbbwYDkMx+s
QENAczHSAJ3frKC7uyO5HNrLGaxsTOmti6gb1fA34cuxGNI9h39ZkMK+MA6CHL8vrDw9BLRPT8qd
k9gwH0RbR8dlRge0rPzNP74m6TNR7tJ/QcDTQKdSWZi/UDO04H6E93ZbV3GA4igMi7Rs5csy7UmM
HBFjqaW2rw7I2yTJb9CSA+GmCS+jT5AhNc/yNLG0jKQhM3TsUE5fxhFXwZEqhMzmT44uciI/jL1X
mRFdPFwylUqkvy3UzdIM7WFRvEPkGw4xKH6ha4/sF4PqNBiShA7RD9KSzwo+kpjFSi+naAlan+qX
EDp7GBb847dTmlW7ZNG3Dd4tJtNcnHmz+xz/qKRAQ57xhJBQyTb4bv5PrH0B0rY3XXt+m4W9ZyGU
9+6X4LdCnCiuGB6uG76ehgGjDvlrMmPSL0r4ZE9OSjJNvW2txO4UAPiNcJMm/uolrEGghWdSHrEL
bdVEsrznvvOGY+Bsee6V5VQuUUcB/OWLAHhpsDTCjt15efK+d8d6b3KgdmPB7AKWubklVNQ9tDQl
9fA/99IVfEMFvvT8tDn2Ht2KRyZsgcX0TXVGYCgjeyWkfEBaR3Ijm2aNs45xMPUawM8hf8nltCil
icwPgvYDiA4o/kGfkYabPAe/Dy3nuAtPuJYro+bfFJeqYZjSFBLh9wve7gxi50zrN50iUuPBN8Dy
cC0x/LLA3uSYuX8EZJGvvOjnf4aOQdNI29lqmgo0R1+5wVP6EalKxiMWBcKsVnH6T+EEy9jndOzQ
p0wMrRvZvSBFW8c2A9qkekQcyLOtW4Pd/vAmzzYr5pMie+32WQNovflkwihpy7dri/WhjkQ77H7N
kTlq/A2GYY5ZXHQDJFUEiNPLhdg6epx7vV4d8255j3DpRWW0Wx6i8bTZV3qjvQiyJLgUGQw8oxCE
Qm3KWiqqH0jCjT4Q/iMpS9DUhWSuAFpNpJpx0gEQRQx16UqD4FcrfXszPpYgwukQZCg1zCtTrNry
MMy7Kbl/lxrc5zKvmsZe2D3R38b83sGL+iX601knQP/ebNz2t82PWXM2o8o0e18Znpr9ifemtY3W
GFYeTAvoXQPWEagyXozTQHKXE39FZ2cU+tf8n47XqZXWvrbRcXlEe4ZB1BGnYLGZxevMe2zHjuIa
2lgy0uLGuzQIyet18wHzFOAVpaWm5dx/WP3wBvw67hmiOWEbAdZMcCKGHgcudO8XTYhT9oLgMK/V
Dm/Rboh2UwH2B1iXI5zzbb3eR6Wb/0k8AyS79HxhcA10x2pUyAwKoHhKQXdgUgX5b0TVsyEEEbLY
0jyak+pDoRi3Gpii5Elfzma/4RAEJnXAxJQgW1vq1b+HZqKWZIO3tiZNd7ZeleY23xKRhI9FNzBH
D2RsCuwU/mKmlKmGiWBvYYVlTInNNaDtiQZ9kwILdfFCLvz425n273sYvHr282pqcamUJNaSSn8V
wZlXE6tVDHulKV8qZK5/uOHwyO0h3jlzj+Yx/MpGX/UB2zr+xGEl0IAqben5UFx08KyEpikk9n7Q
a3NhAHhujVD6qYWgIgi6ygWLY6BH4bnx0V6T6CpwYc9+S7m2KinLJ9pFgahVYsdRO4XX4Jf03hRf
6Di8kT67+kXTLfTE+4Aee6BU8dpW++CZiV13Av5iDzLt0EScq3M+a9VSLxbD71CmDu2p3cTkCdni
P/rQTJyb7oG7QzvWemJoHGFu8DLp+8H45IJdJnsSAMGjnNQkfTF7OG9lQWphcT9ooq4jIArC4abh
HCq8hWXV12qJbtXti3Zh60lhCzfb8HXjpxZgASp3XFN4xWQsQHPeRo1UTT1lUVIGNuIWzwPLSPcZ
FLubSMd/L1a4RbuQd3Nfafc2KUIshDJ+i3PQd2s6Nva5eo5tXrv85lAz8WCcm0seLapvr3q184mb
Wd1YDBAgUF3hWXQ54JIS2NHiOV4NQbgTSW4WvFv+unznJthuNZdAfzSCkgfJfyesH2kb0SyYkYSd
+DIzUxHWDuMA/NDH5dQsR+P4YRJzE14lP/uw3cE0HW4oIAHrftd4ulOVhYBHQNN7yX4+oVYJvjyU
ukDIP71gRe4i9KVcqrmgonRALsKuiBCyU0E8oEdMPaocaFKb0qShMsfird0sSVp1OOhgGg8ealjt
zyIGoeedatZ/aLWK3CZsxGjlN/162Dd+7C0qstVLCK5+NADoFzcyR69Um4hfLAARZuWI0YKy+Gqq
YCJCFLKCOTwh+FWjOZO0qZ+eeildoHRJ/XpA8p5+xRfSk0VYqe6SXY6uXpzBgzauWMO87064CSIJ
a1pjb03RNvMEaJWo8sjXeHJaL/IZzDiVgF2eib7I6F5gOLpuMRXS8DcxQElbFBlPq33sdFnZIsOm
QHcMeqfKznoaH4BFh3BX0p/y206oI06ltZ/YzO67iBOUejut1XeLt7dYOQrKVdYliUDf0kffdmHS
SS27stJ5CULtivPT3CKmeE2pQKGE7N4R3GivZev9dtB7LPFFxXo7xvyllMlwf4DktLchxf1yO29d
fhGYviuOXyxT9bgPZwWDlcCtABRdISK1YV6ydjW5arC+vTr18rQ8rOoNzSQfkttQpyvisjOo0vye
ZWlUBgdYXIUETXMmdKw3yvXFPcaYbigLFOYV0nzvOmd5ij1lYdJsCvIK6jgomxbHY04qbnquc/4B
pO3kqSYT8SQEkkG6nehEExoIhsEWDDju7d1nCzndCeY1F6bkbH0sidcEA0lYBJP/Js/IBlZ+AYiN
0mzbFwG44d3rO72V1eyQbcw2Igk8iqiKFOwCzt6SWbq0t6xRsOzUUHNp/ZJ88JbDez2XFHYZDbMR
+yZtWxAbio7837EELcBeE8pGtVcMa3xQRS3jm1iSuqoJ3Q+n+bgvqdWZn2YlpyV9DOwfB5o+5K45
WRog0W8qRzjxO+EtZRTmmBkczgIgHrNCA1mb6C/aeJGlWFJgDOfNIH8MT48gMLxjupGwe1I//fa0
l0gOHGjzYcpa13NHahQw/vM//OF31c+2AJ9hSRO9oFrcnIa0cOqi+PiQEJ1FIZtv4ZpJyk4hDY4S
o7PGdmi5+lrdogMOrLbyIX2B4aDBbfRPgiWxizK/NOPESOd7MOi/chj+eRQyoDRXFQa41gKdsHSf
wK4dk3zstgN1mwIvK58pwuJSWjHq8wNA7wRhnF6xhp+/6ff0jnAez0NQsLB6/Q73sEj9k1ct/gpp
JOMfd08KdrqBThvsEdPYHN81Ak+yWze/fFNP/T2kLyAKAKcXCgnjgX9WRPg3PQkkvHvHISyCX1gP
T0Z3bSGwrbztSnWFlrnwEkJLfZg7e+dpiAC5K9gFT4b0R+M80XswOM9qku+VeLgb9UaoFkvJ5IUy
3Fc45gNk3Y/P0h+5QNhJoDgOPHScSLkNUHytEwDjtdugo3LW3xthdyTyAHzOBJNTZJJ/tpJ49INn
lkeSjWIhD1nK3yAqQUeyPHgHlwQbWfxCqdEDSvsOeIbMJSARDWFKmray05t2AOF6gAX7JDvc4LsA
uFQy7R1L/bntBoikmyY1a8cRNT3n701YB3SvRAUYi++PKje1NSIutE7WK6ceccj98CDG5BvShMRA
RU8M7ocuwTWB/vQ4vdyS90+xZpwCI3IMDL2teMJv3UrlTIlpOLZ9LYNxOPnxoUhuqGGfAJWKPwAo
BBY/wfs+kUI4V+BMc/apGpnaFdlWb3jD+pco1yTFGuygKGCArmTbJG64duIGwLXrDtz+R4ZsEZ5l
uEKgizBkMkU4RN62Dy+YzSn9ZLqHTbu/m0LOsnHeceuA7cj7cEVXMDAU/wg1Egw/dDByh4Ftd2P2
yQkjWHmxxrfwa5nqIiLV8k79qrzHf25L34ek2VVhSUiQTTVVNGrTimJYI7XU5eKYLQzO+uUpDXjw
675Xi06MfdQQ7WI4RpbsQAA8Js+EqIVnYoR4t68ZrgKSp92JfeDAXKRFACZrxSl6wd7HuAKyj900
UO+zhWLkNzqRTf8wOq57biIj2ivGLTP9bfaeks6BoZCk7KLnUUKjR8S86dK/eh0HCxMwam780cAM
Szl5YNQVc7PwfKVOK2F1M98XKGrzLIJ2GYX3u9au/20pLM1De1hUms6u7IO0ppU0GXudNORWM5ba
P5cr4P7Pgpg4Cp+dJQ1HFdBRlvYpzpEd+grALpJzqVqtdG+mM/PUA4QvfrtMTUM1GQ9CVJyvjSXi
xYlaN/qM4aWuqI9XgbRoyDUZFvXRc8vx+5tLF4I16GvruvY3caSPIbtxOau4w3NMpQ/YrnwDvBLM
6O47Dm5elbX5KiJmmRId+SAYGbz7A153UccQbA7+bXPGct3Yqz78IF9W0ZFByiI4gyf4Sxc5mo+N
Lny0fwWxsm7w9DrfwQbMgZPoVEN0YKuqaZ4LMjxnJpJQN+0S7INjxm+r6H7l5YgicDYebS6KZril
2gUPmIyrC9XQAuo35+RXf4WWO6l+q7SAuZ78LZDWZ651BJH8C+/KJYO3FGwwMYKOPfOUkA0E4q0B
/SV+Kr3Hm9CfzqhiYj504jDZH2RvrxJY+QHCYcL0haThuhQ+CHKvorCjHHrlevp/7r0+v45AOl0G
aadeuEu2j/F6EwM3WeC5ZFb5dl1sX9YuQ81xuKWazu7g4RPt+h68LL7NosgsFKbBREv+uqQq7qj/
uLsML5xqZ1c3l1eghtNU6VGBaTALALr1fXo0RZRn+fD6VybgiYqufzKMpTDJJRQC+iLZRRhAjLYo
UFVPA57sIKrlNEMKzhneaCsvWLVfMMHLeWRCuw3uueDnpXwPyHEVt34isdO/h47AdnnUrCuVRlG6
Iihh/I0if+QXSAYuPn5Qsy73RFdq3GRa8nMtoFf+JQNfLGCTsf6Kz4mxGo6D8QvdkZj5w7bwwR/V
xEL5IriD/Ogs3A4guLvQhStjw0zvZrzKs+cpNEKso7fDwprILlGnjjYCr31fJ595uy8GqBuKr38p
6HOXiCHblG+XOk/9vgaPUOPidnWygFrkhNTN1Z8qu8WV2xkiiKv6KPV7FjQiMoGkaLNUY6WRygDc
UsOcmiPTgtQXYPtmjZQj1dP8BqGyqSViuA+Z4HHdQ+DH6p6InCzN94qZ2HFL09uHVW2zQaf7PItU
jn01UO79PJKSFs5A/CqDU6SBYC+bSo1efOClCf91KMbRtYVgGdSSYWx1U0FrW9U9ynW1KlAjBO7S
doBFINFKbh0F5keYB5/w20kvS8FNkba8GVI4BRmAWWxIXpzf8ZLbgIOKsBWuK6scVTUZPx557ZMB
j8C1mjqbzHYdsYpzW4gjbd8HzQd344Vr6Z72/+kSNsoPwE3gtAXGD79DNas8dkq11JS9EeXTpNOb
LJwoKOxvMWQqgzGCfnDnO5ejso+rnidhWlIUTJV2JRI6vepmDsJ0xflCyBAKM0TkkLUaeWdQUf4Z
idhpWg41rqUzV82dwwQ+Ze90dVKXhon+EMEVZCWgNY5Voc+RYuNP7Fu/+VdYhhL3kRUmdZ6S40FY
RDFVv3hd/ECtZvmVlAJZ8ov5OPG5kn+Hm/7RLHOOdAYbGrSz6g2hpriKw1FI9BWsZ8xeu1PWgg1P
rmIJIffB5bddtnP7DNrAUFpQeskV2gwjyyn/KTBHIPvub3Y/MfoexI0NJ62MAGHkaYEdUYpkjqRI
SiuWnoxU+W2N7yKIGKSTdMd7I4regAweu5o7e64L6Kvuh09pn2xRldsJ/95n3Z5SEyl8JO1KNsY8
KuJFdr8Lj9m1U9GQvxJCeILmC2NkSEFNMvWhTgkpiJDw/ThHHnecKo+DZY8Ezn8plCHuPADU/cBm
1oGO0RTAbmd/hs8AyU6ZtNNK8DH3GGKdtuIrTZW6xcH/QkNrRooW35XiZ4z34tCQ7R9vuxV2b+Oc
XGRFw+4pFaZeAAo9H3QC1StBIHgzEvbxCcltm63lG+Zt9gGqYqXerZGJrojIUSqnFwP9l3+rcNh7
yDKWdyyFijmg/v1TA5Z+oYZCHW1vx3P2oI12W/BRd1w3WVV2mkUs0BfCO+S2MvTKx6ljjbnZtfEe
Vp0dCjMY9evBKOLVbFeQ3us/tfSd6SvaUf7j46N8WJ+yIfYK0PvptAtbnFNoolZi+90ifqUuCaff
cp7gKh8mVmzBMSzCYuzeCixQvEI0MKCYoCpMeizhnx9k7kPlaNf81FL7a0TlUJg1RvMvfM2msjws
4Fcz5Ki4mYwIg3vg301k9luqOLMn79783jwciRO8VOmh8m5mMhEHQ+Bw9Y6WKWvZvfSBHkEBYNIv
fj9Bf2cDoUcpUZLqMAAXnXBaZliJ0dD6I48Nh+5ZMkgNv3JhEIz7/oHW2GhHUhQbtUYuvGPC6WL4
u2wTJsaXj4lay1b/bHqZc4npnzlMx7vZcMhJfEMIlwjnaFodULbwQbHfiM+yPYNlE5scl9O57PK4
mwZ3Z73DwZr5nURHImxUFqtrHTOsxA6lonx6pzBEZJiCkEo+h2Dc90nxOiAb9HA4WimlGS+JxQig
rknh+XiJEQQa8Vs6LX6mFbWbwJHy6hI9avznqydiyFvD2eApTE0mGCxaIfod9BboDoGA8OWjp6IM
R6KuiqDZKTPr5fe8zTFK8orCMFDEV7x/GUtc7XNL136pN4k5jDxoc33FnvoSU02Hw4chIdLfrb7V
/lE8t94YicuWoDpllABOftt43i+sXTeJajU4j2htikn63fHY8QMgWF8zJ+ucBP4+hRFcK++cdsz2
7ApRvb9R5pUQ00mpvOtVwwAxyABY68EO9jbB1byXGVECPpHjWnDBbtXjg24vEBhuO79BbSFtU4AI
KLGMGBHVR5dJlf2rOfdMNh9792dK4RxL2QYHVTBpyeojELDSOFhDM97DOx6DjlSo1jrIC7xugJDq
BJA5AAMnz38oYu69tCJw5u55L2aBTzJ+zssePiNnGEO2yfxSDPEQRBxICBSwz+sZtBSjPwrBvL0E
6a08UPjeRO7hvHqBzkGb6OVMFuOLh4mQIK+Q89qep/hBdCbwFwAwZh1Bcc5+mWpOM/ekz21/5XeF
jn9hIRryOclx1qZwrX3OZc/vQFHPtr1i05b3P6tXeJm+xff0+KtKSDwSeL4eMwwlyOhILtnNNNqf
LzdIVvKyBDsRGNDWt0k29JH1WTq8nf9SaE/gqGoeN0du+ASmg6ZM1q7gW5d2w1WwYqPTgo4PtYUF
OQH1JN0DUp6S38tVPQkFNEuyxM2LEPAaYZ51eLmFGJjYC84x8HpKRaogRdgJt4ul8IBMpT6i6rTI
36inPEaHnIKlhetaKQpF5Bji3x/jeiWBgy+KO/EpRb0ASG+p8kBnUKHQBu8M/Kxt2RzKqymPNkeY
I4gt30jDVJbtXKJZRP4iMEbZwNf+RUCexCwb3HzKcxvOaTKZPcIypX37kFPXcbAe5LLIcpDm5tB6
c7P530a+xcenLonIWuyCHABVxyFWObOdYJHSv1fvM5momC6uO4JuD5VL+oBDGDEyBBFGx2haNMMi
NXocYcv1dyoYJfQSjcLenO974EfzJ8ZlUL+jkWVIhy9Kx3SGpxKx04dv4SvgkbEABX0cmQR39YQT
QB4ShgBYKsxtbDWrbct0iyVS4eWah8YawKBOG/ucl2ncEuozMS8l5DwyNmbSHRps80d3DqDbnNWg
xh5QlHHyLh3mSEof/Bn+VDr+nfMZggCjLoh5TY+eG5JNIM6jsqV2iwmnl8W/xMW2EvUOVPfMfSeh
brvs5b/IPhkkWCcW62VQMdPc/VPILY18gAXDq37PKLN5Pgywqnh2g0FYc5DIEA1+I5IPBlQxIKMF
8ztXteESqJWxx00LTyXuieM/5uvHsagruUX2P8NQ+4tV5zxaNb/2DIO6TOMDDRKrb9dO0+EdkRXl
V9clRoq/N0fyq2GCIHO2dIwPaP89VbwPlRGh85JmPvcRRM6IAKUBslDiH6XI3CYyzqYalQGBcaJ7
pFq/9CYPFCVeaUdsghQn7lV4DV3bIiroMFZTiw67zbkuC0OM5poCWVlMlP+mcVQN/2tVvW/H0gLg
e9dsrqgUXKLy6TMVf9EyO75nni2PpfYODT2gQH01PJVaKTUTD9HJamaiwwdJTsckjVt12P0Bs59j
PSlK1Zbz4KI9BoZsamtTKmwBpsyFH9MMXyIGdRTrnb6JgX7q96/8Qf/0A6RY2VA+niDJKJMWQbA8
U4TvKc6gSyz/xnQiGOiMe7GtCH2gT4PxmixA2ORE3rgwfTYvNiIYDAj2SPGjl8F9wVLWa4eFieGM
RfSsbA7KA2OAklKa/dt9SjNQqrxaIEeWY+DBnqxrb+06SVbhiRg7mTjwB9kZlcmoQndbODGdqdGP
/n4Az8iQQdaVKUKye17f4aShnLMzUDd5FOUooUBcJqGdsWzjumU9MRL/k5QTarEmSgWoBqFn92Nm
QHIiXFf83hbEcM6gL8pwFeGcAMNEz1QMrcoL3QvOcRb3ulvfqSiDZQQsfjzwhGfg1kVPokM0Zj+p
gP05X64XzHGtDmZoi/C5Sy6RADGYk9FaDui4ZvNFhI87VaAbPS38acholqzfBMh5VPP8AjDAISPL
MRxFsdQZTXpYyyZpnF4LGdrl0akKTCzToIhyhKExoq6gf/LFCtpNQeCK14wf71hB9iw3aT9hoXc7
oVmleI7zd0AIS2sZn/h474kUFXAygNhyP8h7A3KRQ07vyX8XdkfkO7vktd5RYSVSXbvjCIb3K0DB
D8FaKYPbyuYfD9YKTl59TLb7f/ca7zpfz9Je3AuHJZykf3JOKaHKkKgJKzFWkNctK/n6bFE2yvEJ
/LMvjNTugzZa1yBCnXafr2sMe08MVqatCwCm0KB5anAFlL+5yqW8BNwLVYK4v12fNwLZJblU1ZSu
8J+ltzjfWOqUqZEtWvl1Z2iCOPv26fZWTxw4mTcu8gVU439SZr/9Gor81dxy5aqgIs6wiE3dCJIA
YaPt9vCN85sO/24t9DT3kaSTDQlnT4NOfJQFZDi6vyh+BzKmhcDrbonXte1Y/5EQm1/xaSQyLtBR
giHUUVIVYVLQTonE3HILG27h7SipNLLnWJEuRzbUoRzuURkTU+JEUqBM1/TFrCKn32StNp6c7U+b
tM3q2G73FbMtTovpxgwlS8mg0dT7piOPUy65mnJNNpvpPuo2SfvDTYm36neRttjlfzcdEa57+AQ2
0G8PyByG+wHOwLckjL26ybFQYSnm/uSvNSmA7yTNaT154jnoT7hRypu63kl4c6Y0lMt5CRz3Boln
XC2Tw5+4Sm26CBUzyDS/qsYmAJrZRwPhVHTgVy4LHeeUtGnkhuGU7w/CYh8FmCjpgccebQ1Sxoy7
o3V5KeLf4nJO6j3REoG/WFsSdoUaiR77mTsELZzk35lE/tbPgyiU0fcX2jbqgRVoidhFI6UfKBE4
2/Gn1E5bdH58nIVkqMeWjyd7uWzb3EVWiz975gXRpXofxXev+YZO7EkW/e7/qqzYA9nsTBCsB3jb
I1RZ21bnbO4052470U+3yO0OTKEkbyg0BXNNDcu+NZRtKIHC2zbzCNniJp6CKDGCTvN5l/m+3MEq
nLtgJC8Fy56L2VyIQ5wQi+yiyEGWYQmt/8agVjbZygGl8QeCg8xnA1hWHq6AnNZuF9expxEifYPM
ekElJHIjd0BLtlPzBpVA/z/m6hu0sjeigK/A2wEuaj6feteHBQfZ578syY3a5/nldfLKy/vJVuBS
dDXwDfnatI/v7YWgk2VFKqXcMVWVERSYdlqL9bexvk8WddZ6/8CUymzCoiD+LUfhFqgQTw6yAPhY
GoknN+3MnrGCGkBAv9BD2a3STY+hJGrmfHSrGj+0G/H0s9jAU4GIjz8i8DLbNr0u53hnQ76iUC0c
CUAH7m3XmL/FBGQrtgyBPS4fjA054/ZhXAOqQ5i1ibD/92a/7y8rq/BWJkbNJtziF3mrD/+Bysp8
XsH+reCLfMv9Vd/O4L3bmSQS+q0NHMbWZChqBlZWGxMnann01c2DoOu6rDtY1CFoPaXYmY+jJ2IQ
tr+NeqGEJhR5sT8UPWXF4/hGGItW/TEOE9HvYO3lJPXIT5V7kQmBxqFk4+ykLDTpcdr74bGL3ini
Oir4c1OqP85Oe3LKnrGXKscquJiy1m1ZDEOOYRnK8KkxriOQkzICdjYp125Rx1k9MAlNhCOIPady
XiAj+SwDp1WuEHstp70mbtSN1469BQBOnEzfhYbKkRCY0oPBamr/XdazIg19eWDjaW2jmI20MQQN
oO6vZEN0I842g2re07ZQd7gFs6YpKGA3qad4bxue/pvYwfQZpWXW0XtiWaDsXoUUKje6T3xafC6k
oVchb7sbs8U+PVCI2QSlDbU+TIytYI0G34yoDmCKVB74OuUvPLbh3XytE7eC/sSff8woPxg88zA+
0MzvNEWDkSO3UanI6p5eu1x0S8Dse1uZz9+NjqMsf04qp6Z3Wo0QnCQfbIttrk9V9qu65/JttZ11
Td7cuXL7ZNK9OWG5ITRGEmZbgnsMviqEFaUHY5IEVJDiDcHcRpMdbdiSN+L58/Q2sUH3FyxYtssi
lZVaRVpSLRfMkrJdgKD3EQJ1pxrQlljESlVaeOhFHUrDB12JrN8WVQtSVHG/YFiu/sr/PlqLNPKT
sHtCLKP95SiOkbqVue8hK4bN2n6V2OlGoPygeu57Yar4/3RnZOGG2CJQF0JwhxOjii/5F15owgmJ
vyPtcKkic3eXuczqBMHUqFmRHJ4a1AnHaA4FMM3BprhO/+JorgFuxV0DkLqu7DOwIdXie8j1jA/6
bmap/R7PONTJ2nO2x1eRy3Ep73of0cnsdYTbogFS2f25DZVxta6vxOSi/Gy6BFzp2dLT0HV2txi2
NsHma43zPJDzrNtkCuFocHIhj+rFJtJeLu5xe8IcNy+g39RM6HNo6fMLjQhzZTgAC7k07F4+lYGT
zBe9skv9Xj5BMl0pQj/wVAqgP4kCPtW9T4eDfl7OVzHNwCoIFAC7QguIAEzyyYWhQr3NTTvsu8An
H85JRU/nIuw3eeKXQNCfKfZJ91r3LoWk53c6HZhxM2FtmWch8BaJDAaKg1QvxDef1T4626mw77dW
Cu2+dglE4P0eu4AKnNDXQ2QPokUUAuYrndR5heVY37KRgODnc/04NZ2ywy+yhGr/CIUBA2waepGE
AALEnzQ/Ca92L6iEDjjxHSbRctmzXdlhyVQWSkg+zc1ot6FOxI/BDzpdxYtRUKn9NAss4eVXCkfP
ngVdtg8+b8msRkN/vKvTPrxn4XJWkeI6LqJa5yG9RaXgFKkIYMQnv/lO123vkVk/u6xIoNvHLu+l
LPyvPf5WOyYpCkJOmUXoKNet9C1Yj0lPZGD0bSTaPaX7VzcEqgqpNOiTN7VuuRkEo67Bz32TATte
F58LUMFyHW0L8GPwZaPkHnR3vL8yideJk9DMBtYhgKL/5SmTgtT8uPWM8x8z5qrFHusF/5MrKC1d
AulF6tBB5aJiHvOq3xsIi550z4nhtN/iL7DLHsvGUH5e6Ba4Bqk1imckcNz26CMRryQeIIPehSFb
kMmx/zL44WZ5q/t9MvSXB1LYgrkWxkMgJEb5z5BkPhEhpaixWvOlsHbGFsx6yWEIwn4qV3HsPFxT
kNi1NImCH1RB9qZNcxgWN6ezBLb8EYHVWfc8IA2JguVp1LwrIn/H2U1WCK0hzizj0HXgBXOdl02H
+bUX0qLNSnHnBODw1OMMWgVGm1U5xilAS8H0EEy0QKFnoYjsXu/netXzWFNZ+U90ldWR3HCQBwtl
xjmO5HcHU3WCELiFQ4A+tMXoTG+aMyq/UPae/yk0NAoOEuG4mS8G6bK9x687Mhbd8A2GaWz0J9Pq
Yd+qNGik+WqlF2OtCzTUy89EY4Af/lrXbKYJkaLhmOlkRIoyxafjH/v306TZ/GRjyqeoiX6nccSY
wOAxa4Ulc9G1w/LUuGV+8Qo1lgu+sAk6//tGQZ9sjEvYFKxtswHmkSSbCqIyPW7B6Pu0RRnqB97d
OMr8syRt3Ht1W/DugQ4U9SS7dlVKcVRjOBb2VRLFKIGLOc8at49VpQaGPiD6sqkgSK0JgbWF698K
PAUP1EzqvdkZBcXqVJXLLaNn68k7A2C3UHZyust2C2Cv79+ucBNPE24mXwS4hLlshHDtVlNg7HQP
0rhrLQkbmjEma5+5rp/QUH9rvGz9MWst63LdESo1Kz8NjhAibsuLkjxw3X9KyyEatgiLyKLWcJbo
RqmlviCFCVvztGv3dj3axrcZF4se6uVGCGo7XJz5hjqc7sj/1kl+ta8CkkQdJ05tA7g9HYmJrQWK
9BGataFnXzMCuZpTuOGnbPALNQ66dC79gN26nQfeA18GGBg7CYcjQfMX4emK1EXNoPAkVACVaSOv
kTTxfAgFAcpKMdiahBQbr/iuuD0rnQfP6uhY4PsbASuKEWxZh9BcvYIx7ffVzpt4dFgLIHS4Ab2+
fvgZSYGlNhI9ZAbpHU18lcyoRYT3wixpjpKSxnRE0rhgq/bNJr/jL92xD74wxAIKuvJnXQUR52rv
2xvyRTthJgiAx6YoD8jlxjWCoRujkawZQj1v0xrmwjlOX0Iav39Orrg36gks774TJftadby5QVxg
tUzSWbD+zMhwRlcPb5SaUtan1/cetoDkT7fs0WUv9D2P/zQmxOjIl+C0n2TGjV5PSi6YGiCq6YYC
4jF4i1+hBwjvuTmRP9ICAQF1kxkadRF4mTWSgC8WQBxTn9oduAVIp/qtPM8QxOoQYOesL1bYHwgI
62Sh18Mzl+ga0AipvCJHvTlrJNyxkEWbyXuVC6SU5wB2pEy4yUbL+4Ch/byAbyu+GPf8Z4xXwAs+
S2F+Qtmv1Rwx9sGyUCXiIKPGhYxYtkoCTXmAA9fS1SPbk6CH5fLl2HkODG/9EdTQnhHfB//6G3Tq
oGVwoi/LupwXtRU102+2nmr1cxlsTaf5fJvYy/H1HnMTauGmKmOFNegE2NVZ2qZn+CL7oeUOPwTP
f6Wqx/oJB39sxPk4GLh9sFPcnPSOTfWXLgKmpLof4vELj7oDBOqOAHXiEZvWe8mCqnwTFNjUcWUS
2IBDmcjJHlfh+lI9NRqUEUt+8gCKMax77eWNgeY+BN0JsVIf3Mk3Shb4VyuAoXS7klUZSg1AASOR
4AOgSsbcNRHt/FRMCE4A+punscWX8lZ/uZxO8ZN+f0t+vCKZnfwKIYPS2DWmRAlmvN9aQuRApfcn
OPecDZvI9f0h6qFLB2s6WQUcWuI22fv1JuhZPSTeZOnsFsZlZBuNIIjIc9ksJnFzcQE1E1AtY9bo
EHzPvXbTlqsEZ2zCvqhEUufFegk1G6zp2tPVj9DvoS1As1LGcIR6cq762xKomoDhHwpAEC03JhYT
QetX4hHn6p3lUm0KhWq0CRZY1ZTOvReHvfh7mFZhhXYTzNi/R1QmsiCL8JxMoMA6VMchX3dQOd1i
hJEbWmuWQ3l+22x01WnFgfJLz/5ThOL/EKFbEfwEtDbBRSqFHuD7O/+KHX3sDNLJaUM8TFNxHqpV
LGE5wMn4iRl70WSsPrpPvuq0Wpl8bkX5KEW+5YDy8loljqlgo3vlGxdWZF4ph/tV740LnFu19JL1
aJAl8brqqpGqlpaxhV4O+mwTNXJBhk2AUjzVAN6Wu8pe4WTfI7hNhOPk+8Fjt5AnSXq/xKgduaRH
i/zpYBtqm/iPNFCs+ls0N8rVjkzZ34ni7meRNIoaeWfxWUgCKG6e2VOFZPUvq2LefwxobPj0b+AV
QHVmprT/3G/bO1Hxy1s185VcBKh8TPzfTzKAqGmczPeyP9IQ7irmFW/qUmK1FoG/ODCrjQBntuLG
dZ1V3wGUs4pSJHCsOZjsf5SkPja96w83qjjLeaFs1gvrLEPKf7OMhLNaNLhfhwoAeRuqSbY4KdpL
xqUlbCKO1kd6Z9yhwUPDKHla3y29kQd3rO2ONx0G8GiwDmqnH6OlmjBwMFOx+S5T/O3TmbEhPCDr
CKYNkm/9dCc6Ag9oMpqkMsUyUzYbbwBicp/3Ky5ur4Tuau6fta13lpTM7UO9i11Smtcxz2Sc523v
2BXxfEu1xdZRgGw4IqTrMh5dE/kxX+pfmuuUd0B/xru0eWCy0zXPld1XpFjkODx8DMXf6l9kGt9t
OGROC7wmFqVk9FSbI18J8j+s6A1vxwvDfCzikbC1UHv8E0iWj7asgHZhgFS3/StTAb1OJcZOfrPM
rf1K8RjRdJO+bdZ+uyBu5xIk0sE0WiAohHRVxb/SWEe+bwM5AVNh+JeFPkSVGjNucgRzBm0DHOgC
ViQPV9X/rBDEupymNsyDI44t/4WoV3kHZ1SXwbTgqXJGcHb+j7M8Jisjtm16K6VKjrV4f+d+j5FY
eDaJwNfUsgnI2iiCslu5zdGN1XMWpCMN0Nfcbb+MPgqoxs1MwzvHa487b50BheB5uqz3YbKYm0zb
i70J8PpMLLcoTQ0SF6rUPdGKA3gNufyWzBhj+ZqXM7pjB735YN03HPgCujE0MQz3ga/USx6cWFXQ
AjkvPDQxAEyQJEOMjEzQyRSu5kdmaXsEdBS0BcD7y0JcbvUTUnPw8oawKzLtL/kcxcD9eelbP7kP
W86ndahkE2OvRGGyNwwTn+napM9GxNoGYECvp4q0AdoMXQUb5JWtfg5GKKt2s6KcoUjdXBOnNK1i
XhaKUMG1h06EJpX68fXCt+vhK5ektkTUnsV2GF5Ao/xPCmlKQkYGQ5gXXX19LkgxsbjkjLwstTMt
RLw2WfCwFpWf6gqiyAdbKDP0CQHRRIPKuBZ03c+eisagHtWBZgsYXU7IY+mKl5yF7FwU+guUkOVR
92/IjogrpWkW9nAVfbKPOrfgTuEXcTQwlLCBoCw1hCVu4msUjATP2Gpm8FJOOfKfwtVS5dTM7HA5
nWLJtPV91QRm4RJqovbKHmfe+2FMmd0Ro7fj4GzPaKdj0Ukmr6WhTNSkPaH2s2G/bpi9+nYnRq/h
MsOBmQYVzhc6LMPUhOxTsJzhI5pn4fxFqc4I6O9kfXRv7t5tCsjlcn5q4Pii4UbvfC+LbeB9XdXl
ihPyroStut5+xyTczi6s8eh+OJ3DuTnlSPQg4VA28ZSe3iFej+xjAgOl1lIfJf9HXVq2V2gwXo2i
Klh945sTiYIk4uEIf9VEJV25DG8lCokBkV6gCcR9icV7oTRRigHLvnt2S9/xVAZtSnBnxY7cUkYJ
fMLjLhUG5CH20wPub1Z5u3/9zqM67cvCM66CLKwhCBBJtKau0w5iF65JRrZ2VeocXy7QHjblXFgO
tMOBZjCGhFXnOCMn4P6+D7hpCWsfbJkRDtPBAc+iafCvQqdUF3k8WFewkQajCNe5HldwyEib7B+F
fP845Or6730t9DunlY03pSkW98qC/GangTlDaMpGi5FZokMClciLnYegrzKKKzxp9EJ01AsJ8PFI
NZLAXDYdeOvqolBfvQHBeDW0bN+CZllCq8ttFji9aCWCoW7NM6sRtEmf9cuhszLrw9WzAt5dVIre
Lm8MdNBqOUHR8i47IWaHF8ah0j8ZOk27NFR7Akvuql1APM7GULUBK6txb/yy9/8e3nCuujx80RJ9
JB0Ivc/ZaXrcjRybKtuHvytpClLAX3NigYqwG6v+6a//GZomjAM2W9+wcHfpf+5B1ULH3SNsgOxe
Oat38IA1VliHjV7fNXZ72PyFQJKLv8kqJAktbl9Ib5QN73P95XetNbMf8iP6EFpQawHptENCbvIG
3JoPsoJv8RTP16tGIHcTl/TbxTOqxF2iOC4t0IBDfOVibOtzeQTLG4fiVPa+em47TfupC5yBvRtX
F8rGx8Rx7qMHUSWeBFKa6hJp7c+ZBLtkLD13jAGOle3YMTUGbYOgV4HaDWFwliY6bl3UOHojg2rM
qOlreMvPLfHOMLF3qSjdnA1rwA02Sh9DP5XPCoL71dejcgFPAvpx5YT1nRhhnyPuEcqiHY785Zpg
LMZFd/jf3pofQ5wh7k5Ii0cQXtYeDS/i3eEDy7EW/MOcohkETURFrPzQXZsj48nZcPSq22fRTtFF
1ByV7ab9Ein3uJqW66Xqr/n9AQDJ3CwTNqxVwbHHRcCfnpU8HgUNnziSYlvczFD0R9QYXfbqNos9
Gh6LDpKJw9XLaYOZ2i7zChgu7sL1XoBG269VusBKALeO4Mex35jf83U0jTCY8E69FqPn+IkID+v2
/60HVaIawE1IiDnS18oX7RvHzIHY4pzPKSZe0/X5sUIAySLhSsbz4ZKoqcnya+MSgls/OqLvFo9J
zYoFfzhttgC+nbhfCPkAxndNHbKXi621jpxRwreV+zRxuX+KT6JwyP3S5PHH7CpudN4fhTzcLfl/
gFgYCdY0o3gNRwyRU9Wt7TNq8fPB7ZaXhe47JJlCmaNVFAJwMww/rbAa/85CAlQiAJ75Av5TxwRG
NYEugpxrU2F5+g4KNqUWxZEdNh5oQhomzs68W8jxFoEnCoK8z4vb7QDAh3SAcJGVAiT+YrxvjMtg
NDX0kAqcYpLgZWZ10cZv4jzVeYjukQFds96rHWdiF4iOnsB9UCbrdAjaVgv+7KdfZNkCVkVEi1Hk
EF7/WXeLmeeiXhFhQMZDQMGC6QYZuVxIgMOwa28i8dd5qz6I0KpiXh4IUvhHp3pLr1GHGPdF6Uv1
6DRPfiUDnED87Wxkj0rOZvohQ0Z6Wcxu8H2XptnoakzCwX+BJ7uulDRIMoYoFki0RtOvqZeIW7PZ
WI2pl4Qcbrftrwpzdq9stggUmh0cFGN4yId3A4LzAwdIG0o3UkaOzcUJLLYSuo/fljWsck43Phv/
7f20WMVRl4QNi3PzpAY1HjyUP6vtnVfobZSSxYqT4Vtd28lfg0POluzdZRzW6MW/DcRoqcbp4yky
t31LO32X1sek5Oe0ka9HxrTGw0/TdF2ykqm5Su8ee2tS8CCvsK/NCsiqZ+M6WgAhgJP/JYdn6Alg
r1LNkZulIwcjKiFDJxolkdH9YIfdooLT0cKPPlq2S+o1SmDzkemsSvEzBPozOqF/SGWnUD2FsHYd
VuToiwOKt/AecjqcXvcIbwj2c7c1U34grcoeF3uEsESYkIQXxgur/35xPZUYSBBPlRE6T3xu0/oy
z/KUwXzX1/LvryKcfsu7ErUSQMvhFflGG7LNghpDqfk8obQC2sGJgFLYxJUnONQZsExt/vvSUswL
uvk03rB2UxgvrF6aIRswUBrmarxRZXZEF8E40qKGC87g6DM9aLPtvfHpbgd9mJsPrbi40GDIvYsb
ClLgld05CnqyeCeSPKpROsNYqJhZQzwGRxMoLPUl4zaStQ3K87LmvOWdJSe/EIUjR492yiYP4B3s
tfHkHRzHekqjFvS0H0Yxqtecq0qTZ4JEBZMoznDaxmD5W/ItD0f+uZa0D08g6jHBAvZ6zhNYv6ns
dE5RNvds3x3HOtgfrab+0k4vbAKEcY5lZWV7dXCwbv9HllmPhE01ny0JHz8xylGitXc79P679jHr
AV1UEbOfmPUAgj/qu2/I3pvWrFeX1IwW5tO0hNmgtBHVWV1cbsjGg7ThcFOGtpwCciwTfCq0vJSl
xi+oWGHXIVZW0qc45ihY1zaBTRqDx9NonySzFlcxmkoPw+CfbT/eKupOUihzv0Hg5cLgh3cro+q8
1otuRXOeDtMU7PcyxT+iyejHO0cTaYqhgowt/tA/Uv92s+2Nw3NfLLuc6MsFBOF8QjF+bacByWsj
5FYyUps5+wiQvudvsLPQZ5rSxVTOrGt5kq+7mdNNFoqaO0DVbNLN7Si430FfcvIIOCzbv0a1TY9L
MVNRq99w1GouIjJ7K4JpfSl8RuMdCgcbr4RBY4pNDQR56HNNT9oXUVOSnHd+3fOXKITJUTgxwe/j
EP1Zhv1xLET/hcqou8xMyaXa4tzoemVtk/Tmh3L9zDr6u5VcVlny5K48/Lo0s91usSr9FVEpuZOD
SyEqe9QbOnLudwteN9h1ZdtAqW/1vIXsuWsljDvYS/ojMnoKME4IxjhIcxTtnza/sTwnaQvQQQOo
JdOLllEKRmAb01WxJOr/98a8V1eHnyfqWr9/0o7JeI8JS5BynevPv0Y35F4yi6UfNTSNStPHcaMw
cBB30ahk7PZBVSOXVnXSYPeKxFobWruaxG9DbaFHonQCJN4G52K8CrrA2Oq2+YOaDnUQciNdxdnb
Fk5bDQnYPmiub7+++YiEB1AxKD0WWUSH1jtTOFZMTxbXK6ph+7rgZ/PUNw+8lDBwN5sHdhh9YGJ4
xFfwDFNOVg2MfXeLWQnBeOA3juCmpZyXpBv7cuk4lLiZS1e/AizV6+HWhmGyk3DjajsxffgvMkBj
dXLAc4RM6iTwFDX+fRlsq9sAodtTsJg2Hhkyy+ZPyh7J6vT0hZ/UN3YcYDITAD8PSbCXgnhPfKoF
hK4OnogLJxuOoPTfDVwfTh51rPgSsYJwLu3Yx1PjxUwDi3zhJja+Izzcyv1raENgkV/UCp1+Hw7i
WXoRXl6cy6mm//APvXGJGJygqvGYqB7Ebf3TVum94OdlP+lMaBtomPXyTddlKNOqeURCdsAACSsJ
wWbJVy6pYmKwy1cV6a4CzLN1bQgH5g9t4DYQZ7Al6h5I0Ltc9Gr12ou+uBS+ydTeT9AQN7eGeosM
PcFlUUqgjRq99kYmFu4hamRo8NUpT2RHAi/F/P3sMoonknZpuYSJc6MEJWJ7JW80UCTkbd4DgNmH
jNVNzgEOacg+POsydrjO+e/lTivRMfS8vy9nXpqDHToNS0ei5KO5SwWdWt9dwfat9l8xIQJhtGSc
XMKKFaDYdjGCA0sGCdJUPmvh38E8Efw03Nnx+mTNfOflztY2TyXa0ZdqIYeEyWYtN7X354dky7FB
J9XJRVE9YIRwD1oVGknQv1pfkFP8OMgn1WPmQsK/00HzPdfu+cK2fkUw92Q+dZ0lIO8yNhmpK/Yh
HYKhYzigcD//4kSkRenfhQ9RhOXXx23R5mPj5zBK2faVmcjE4XsslxHm8pCVevL6eNTe/VaLSF8S
BfM9Z3Shj4sBbD4Ie+q4V3RBUXHvYu4igIeDbLrzqU4mQy+btCeUrQYSwOPzdJ4NWrNSsEHAvacN
BFyAnd+A5/zii7EbhzJ9js/SnwhvLs4kADykF/Fx+XFaQ4UUqfWHUh3p8qnxuw6s4k7YcBAQMAQ5
vp8ebEqKo9CUVNzYkSVGEtoBjWxd6tyKlj1kyND3uylYbTr5RuKhmWZk2EUKj5CRH8V2ZfrKzee6
pgdnc8E3VXMV/51ND5SvazuLvsS+dCUaN4R6E6MnhTILS20KW8ggr2mnR45jyadm7iCMyp202UpE
pLeaznqFG0sM3XY05Zu3eSAmqlq7iuhAniPmpZjQhrdeOYKP6PrRd7XeuF9EsB+/Q2fTmCEDZRve
CCoyklldw01BTXo1v6Tdic0kycaLdie0grRzdURWwgw9nQL6JWIqb2zUj7O5dttnDpbuvqAAebbF
WYcX0vSYqVuk4f/emAvMH/9jGXfgyw8Ht8tDbHPpdQzErxcc4RRY7L3LAbyipEeOCHPY/UFdZ8KI
0PTVOsxxiSLDfhgGLS2tcXiFO3COhX1IV6RRIxXoS/ovQZoaHURGJLUXORGEN5m64MoA7Os8Iec0
OvsDO5nkFrfZNxgdU/iio2PCLclD+2V3uS+V+U6mpb/DnnZmfMOSJAjpng2JlmNGUOccaqyqQ5q4
RTkRBCJe1aeU+3vYYgTRf2urfFzDei2d8SrvUdkfy9qX6VRzRQ8e6a8F6xjPSaxE46EML9WRPdYw
3aXfUkKpRV1Zy9I8MZJtEJChMORlC+qSYfbLKeBviqnCM7az0pDebN3ZZ8Dv+jLYfD1MuEgbwDqX
/FSnz8mbwKAVm7nCVwltiFar4rWg0pYIXD4rJ2VU11p3MIY7807pUIYXNIf6bX7dqp8mMHty05Qv
SVFc6M8NgUkDFytPL/Gr7DXcJEMKyz9RhsTECpjQFnVmtCyjzouvtPcm0/petdWWczI5qI+r3Btl
0fPYI2jufYFc0BN/jZO4n+0E8ZmoXgIBhHliSi2HWBddoOIPnA6hOkLrIKJtX0DYCjsT2625nZ9u
Oimc1/Il9HDORPl4G4BB0BA/8iQ89HoFgpV3XT47+Y22R6Rz9P3aWRqPAtBchvb4hmreqx5lq7ut
nbWyjBuxg03ZF8TDi+TXy0Aep1LHAM8G9pL0dw5ji353FAZ5GBXTjLMuuKgqP6NgTchOIEO4z4ef
q3izwNaGp2rWS3pgbiQ1E6W75FME5TJJQ345uSyXXQi+23a1syaPDgQN7nBhez/moCtFw5vDttZM
Bp6u7A/sgtnbeELYCYEM4F05QLf8Y1E+8PgAAZArw+VQq/nhyA5LMYj+k5f3o5hspkniAVauBVWs
2KYqhf2Yn/TzsM5wB8KuR4hJiFdt6/1trnbAMP45c8v72uaxqQeeMr4VY44zj4QBu9g+TgNJK4u8
GdajaPKhbMGhV6R9WUSj4q1abInfiSP5FX8rMzxcYl6moDBBRNAD8b/v1kVMApZ3NjxG2kyhfQp2
Ey9Lq0u5mfC+CY7c9WXiYxChxvTvKBuaxtEjxLR/J2vbkWxXGgtt4xQQldV1ts8dkXqgs31x0IXc
vxFiqhXDxkbXR4JJG6KBm2iVo/bKOJ1bcGjqxfQInJ4AgfvYQdrEYT5XfsaKf6fTFYaXLBlqh+nW
nuHYq2XQ3GbA/j8lxArPT0AoPeGNSXY42UdAU8OSKdiOVSfln2gAxGvrsc4jvfwEzIqu0myflR8z
n8+tT9zp9w8mrjr48XZ6MEfWB4D/RIpOltccm9O74j2oHyX5e2aEN6l2u8nld6xJ5j9l2bBpbODY
uPGZqlAsmFv0ogHZwSx9t4IF0kIrpGhsAMhBA++aybzCqmjXahmr/VAsWD8nREtEW+k47aH61BZE
GOTe8Nd/neNNX+OhdsAKz4wcH76P+vbMFlwHilk/z4VEHtUjxMEOKEGy+XRJ8s+imyMxsRVOfFbP
Szzz1tHUzoGmMDtFAWY06O4Aex63bgnfZiQ79ptpQFL8Lc9wrPH7taBtovOpQA20m/x9ns0y7IqY
5xnJ0/VLPq8xIV3PFBQl/jiVeGsoexwLhmn9YnAjONclechLp92rVcDccKgAaL1VzYU8R+ow8vhP
6uZnyofkZAormK3hY2pq4GaOCDQ0EVJskErdfAelMo3xXm6Cf++oBLasplv+dR9nid9281koQfc8
mZ5XXo5scY8pTUg4ABwTckpMG7vlUz5k7h/Sa7Bj1D2nJUN4BpIe+N9AeIQFJ5Qp5pN1CNT0tU4u
pchJ41okMfpnlCvR9I4Od4KsgQN884mPPCntFq+Le4pseYKwuVAQR7bLlFA1sGeGL16WABeRJNUp
zehVcVT+xHXYs0L3t01Ruz+RxpIDvZyA8wyT8ktYjTOzYI0tqyoeCA8R4en27kWaZGc8K/xJ00xq
MIAu7VdOf2PgVm8oE6ntA8fS052F+6yWUP2GWYYq+EOwxOcKPQPDJu8/7WC6SAvaVj0Ja1JY6dgt
FZmiwzXyZ7wR0kmdjx52J1KkmkiOxyNF8hQGUg+PKQbE+X4HmvI+z+BIhr7e5QvPCs/AzOXmbZfp
8EkU5UjLi2wPeVs1qog3BxZNpdyXsSu7rn876eFuOQwINNT2dCbuybZvIsZoT2hcz5pbr4iCgJsm
TWD8qjaKR/O/zOTwQ+g2uPf5nwTFmzhIoYzjmQWCCFJ3mQV1MbCZDs0//iCyA10JLLLto8O0rRP5
7fBoRRLUkig0v4mYOfO+diUtU36kvSrrA1v1mLt/pWl0xTj3iGUX7iVIAnM7Pbag4sRvoCyLu7UL
XSh4yREMdZ9tBRrcSR31YS+8WQi9yjgERmz3nuhjMzXvh0x9wyRpjYGVJkTqE4SuoURgwDlZH+u6
zvK2VsTR1IywOgV+EFWCOGAKT1WduH+ZBdOa2/NqUsC67J8LJjnOW9o4ZhCfMUxBQKg6UwNibYFd
SgbmSgeNt5KkS45jiQR3XS2Wn6tcRccI60J/56k69Jr6tX8KX27iek/p1kBVuW0Ajb0JTQaCE/mT
AqRUrGyvtvNGvEhwm3vMsjDQABXPU3MY3myQNvjqb+KR4zcf8gybpS2/r3ipIANLLG6fDS8WQ3ZB
9Cj/xZc3gtx1NL91qhidK7sWuT35yPhlS+/RiWGYRAuNVk+I5Y7ofEzmEBjDYWB6FHJEZ69Z28yP
mawXSi8c6hkiiJXENCcA9mJZEB77YYk0xSFkLZY7kvEqVRd5+/sF7XETEXwF0wW/9QNa0FWUJl8R
lvYRQ2F+C1uJWivdAUC9sMa5+yWN+ZRGE1Lm5k/+GA3uqwdQVK+cgpwJLwdVUYvjTRhF7fvxW6VD
p5IBdERby+KsnH7Tr7+EiDNC2xqumodf1QgYJvEXmX1cAhOQJklzym48sqvrakfqjJhbpdEX0Ks6
sqB9GSM789zWPztV6WKMVobLpJX7Xw2siVDmENVpAKdiAB0uZ1kNbcPtjs2U/weSXdUgXCJuWqpf
zjN73uZgN5aXD53PcGh1HwFGkrrlK3HbQg5a7ZJEYzBnfBQOwWYVwbbjpElgU0CjfBMpXC7/3TN9
WGz8NOXPoafcnQ+dEO0FprfnH6PeFfR5x2COJ0i3DglvTSjLJeQ9t5KbAmJvcpy/d2uYvK/3AYGa
+unkdftkE8noWJZYDmgngr0IDZOH0odDUKEZcZ/mjwwGrljIIvQBppu8KBYtoJLLw7MlPPSg6TJy
dK63Fj3DWcCFl24Gkqgs7UgHqzH+wsG7DvbxrpwiAyLdD0SjDw3aLHGf5ohb5cvTnaTV7kmxpObu
fwblZv0Aw31PT+XgtxoR0/u9K8HgsOKEMsvC4XT9fGExCW+VIwYFju83VDiKPCMkCb1RlnhTkjHl
NTalY/fzp/5BSK718tCmrYiJSgfguTRXU5B+Y6fPUgTF78Rvz393EyIkldnWHdjD+GjBm44bRb0a
kWYpAJw1RYY6HX4TaWg2/kZIMRmmk+y3MeCVANfw7x0s36ALqIPKSFlSQ1VrRF9hSV00J3a9eh7j
z6mlDXp+oxPunY25UdfplOo+MncLx/QCLicc3I6iqNpaog6vdnrLmHirTkfVhzQkhdsBwcSDZUBS
Rg+5kTD5DiF/dfsFvRz9PzsbbB6l3Sgx8ZLgvGxRh9KTzF6o8I7FjAFSaR8qCfctc/QYPp3VRgCW
RC3rXEL5dQY6azkh8vniZ75JHKoAoE24ul298Whbjk5T8p+lVWyyLACrdJfHYSAYvReuX/hBfaqV
KWSFiWqN8upjd+AE2mwkKeJzhW5t07/ijKdf1cdZ7nLZvUxBivy2RXyfsQa9Otyx5MxUXxqecjm0
KIuaVNJGthd7V5qPi0ymiJ3GQlTygLPgxbUoPssq2OBUPttjFnlYBJYopVZSFDAbs0tP0j+vIFrb
bCKkhRA2y9ZkAStCcWH8/wCb37IQxDtOYUTflxZSgr6Oy/lLMlEl/AsnOAYFlGfwtg0Asg6gioRo
PLdcmjlNkPeXGXItXguNlSUnXgisIA80MHLN/NHuSS+yCqRYm8u8P1xlfO2OQUh1RowTZ3Ze1XWK
3dt7WQLM3uI2Oguk9+v60mGlBOb3mykaQ4Toec05XJYwfYWT0bLEcPIIhc0uEwVmcG/g+ke+jOI1
68Bztm44hNPfU9FClXj6+Ej5SV6r9H/birZ+eKAfjqcPOTiJ2KPOLyFaNY7upnoeSrccNN6It5Ym
MBLjOp9EYzYBuS4EAXb0Rp7Fbp8tcXvq9aHNqXxSvZ5eeQG5FAWU5Iw6a8WgUMDyjzPelzXXgz61
0PoSH55K4RcZEzFZoLO80lVKyu/KpILe6ywL8DWHEh2g9KMn9Q66ibvh0I55eAigbN8i/dY0osjM
vwueAm449/FDbFmkKYhdG/StEwakS+mZ7u3b55phvUBP87HWVw7bsvWF4urkcNlJPZ+uE4nRFGU5
1ahBFvoYaJytA1OcrMW8r2XEJezgvvF2H26AQL5tRwCLfvt19UDESNeZP9gKFadCQdYlC7+Hr5py
mrVDLAF2RKPHTwZPx29rjqyP9GHTJyIBogeFyaCb+E9XfW1rpvKgDbrLO+YgkryLspt5bcneYIr9
2FrzPjkrcZUHxnoroj15mB0s42fNt4JU+QtysmM6AOGXwOgRG6eVStLa0ApSwnFViuNzRg4axA0O
2cfkJY5x/Nv2h+y2SUZ70NGvMuF0H/7lvToQJN4uMG+wfOIUEOOkqE5w0ogRBjDPE5g/LvC2WqFi
kil9KZLTaMOn7bl+1KHIV9poZfu+twch5HB4P97A0berB4X1GuytKTjKMcQk6mOQVfomCTDJ86FW
LcCnyiWi5821qhzcbUTfzxkp3GzwVDokCLR3xVw8vB9lPMG7YOgJcJnZSntfkVomTl3lbr3i+5Sb
bNg5THY7nYkq+PnNH1NdoTdr8+6lTM3BO7uMQsQ1jRDF/Krm3fYyZqDPA0M9ykX0bNKtc//UHzkI
3d/Toc16UoSL6J1YGI2EHy89Ei84hcqKj1erGGtec1s0dlGDGIwmAgK8QPzDHOjYwnIrWJWE/ZEt
IKm1OKiSs8sXwVZGUGzOqSYw1RSYQv2CWFmVScW/A44ZK1W7kXkKsKeaOekf+W+yeWd/5+LbcwcO
5ITAhJiXJkphUYE1vx2E2gt8kDcENffkJOz39N/JXeq096uh+ta+2E21febqCHFq7/6jAvcfILPK
ZV6b7zVZ3izj+k6mxC6f2mYcwCdG7by83jdtJEZ3bUNlopBSPSbgQBopc/cPVanssT7goX8ZLJyB
YhiEuhKN/Oo4+Es5wMi3y6ibRkILmZ5/pUHnR45QmNnwRbkPzOJbUpF7UY06P42Td5/WXG00hlD8
6AadaKTnq6mPTzpZEbDDx85hmY1oaaSxIQDQWHAA4zKTNYNrey1jY7P3PPiz7LKtEgeldT07GWzd
2vpBb6HPzd1ZY1rwAHdvzBjy2zQYSOpXZyiSPGTOeW7vjNNRN4hMyf1q+eJVKCfelCJJXL6gq8cw
ESKqpbpJ7mz1vnPndx5HU3q2lfkw+f9/o0LDhImYKefyHGM/wqG+nN4Sm+9IeXMS8feiA+AyMVAX
2bDbkRi39DwEAGdVFfrIWk4sO8CFbCj409BQCrw55KAtKgvibPRrPoDqNaTtbQR4472VvQlNVPL6
e6faagBRI2/Xv+1QMsl/5ygiyjpcoy04Qq9vcdStecYGxZvi8mAd4Fiz4vt2MRtSswL9T9/N64R7
QvuU2gip4gNwpzVYdNTPiIan9g5L2YgfN4yv4oN64Y3rcqeb4vm//NNF6AtGJh2z8ieV8TeBFlIf
9mfwgYD3lzWJZUsQmsSqGFornA1SieuF26LSWdkbL8tOZ/Vpye3fYQCYrHp2NK2JZrTJWrKXaTqj
4jVYmXpvGkrI94fphQ2eGqJ9cuaKx5vG497YCTov+1mF8z4YwdKZgoCz8pfMjleweyp/6hNuw4za
QZ1dmPUqRLaMOCkqzCBAT2A5MNRpJoi6RSGa8Wruo8V9dgEVhJ4Chwp7AbIbSgcF7qX/dJlv1ToB
B/KFKkxU1DRwoaoVJ/DWFW21bmXuXTFost+RKuFpsKnwKDqe9X+K0xFzE2InFvVbLPZN1FVwLCDQ
+LAsHhd3OuJWRT4Wud3YNIBGDwtqt+UCNN9sVH2sIniQj2qyg7raQbBroonPjSwUfLC9+m2hdC64
NKnxcvdbloLYJxpDldbHA/S8Gf2ZWOGJe+E1mUMRXbca9yiIuBBBxsspXXW7M5LLLuk0kuSX8F5B
CDtEHPXJv5OsBfSujHnmdOJxxwYAFI3oa2bWk8KTRra/l8SRV1VL4iSKkNXQPPzq4bvsBH9z+7zH
3qlFHmkHHdQRLgf0wqbclACEpIpwd2Mh/zSFm1wTko19/QOnwJKDG1HkjrSKCV+/B1xA9/zGWalW
aOkb9dTudgWGUnT7u9HZfOIg3NZ6xLbGTLxWbzS9c4GL8ppq+u6ZaA8QInY6DIefNzWDz8A01L5z
OCUpnye3e1cZOm2cB77YB+B3slPH/KbE1c753XiHwETfby0XdE35UWE80CuvH/6BV9VGtrnw4hzr
Nly+ynAR74TYJadD4Ob6G9jOQLHomAcS130SSSMLWY8xrczgrfnDrMjuJIMS9c2Qp0/dW6H5D9zD
99Ic1SfIH91bLACtvsApEnXtzo5A+7uaO2ZcsnVlq31d5oK3oZC59itd6Cx2fwhKKRktmunvk4V6
AQ5TrbcIDZh91+Q3K3xHglnw/ay9YcykVd6MPcN+OsZCSrTothEh1tLH3oyBReOWSorWPeqfOpKC
v2PGMN/uV/M7wyTJeMiXagzU9pIOAR65fJg3MAi3z3CBPbUpfXVhXzw9Nl9ms/GBO+7w+83/kfvw
3t5OfVo90xo5a6BmRXSBDjGWPlFROTIcxPfz583BasRxMnLovOQC/bnzzvDDYzh81ydrC6oDvt9F
RJRS0t8bQd043me+j7+CbYhYIKKTXNFxaSfjAzZekfRbXbTk2e5o/ybooD/PGt9SpaDO8Eyzr2cQ
oXfshh7dFt3FmBVklB4fhxi4/khr12L2w0OOij/kvlB4IUAibf4nlZmRSRafNCkIZVULUdJgayKF
oY76xq40eTYaIv7aljyekPTwGXjBUiZBVIuHpd9bEAdyUUIziIRnexAzv8SE+NvdVISLrBAY7mFu
b4uwPG4SB0nHr+X333NRYCVs+X1sB+g9yW1gdFsJhMogCQB88gjoaTHGfTUUfrzg3a67p4SCOhND
cyCiOHibdnahe3qjaic6N47oEASP7Swbd7YsLAbDlTCguVX2mIl1Hni4KsHgmDTWhFp/v4FZl8im
yMpCdLYWQuNveJtrWSBVwxKIbAo8DDLOtY36+SyfD35eSRJ+mMPR08EMZs+vKzelspYIhp+dspCh
fAPWsH0OBHvY/ByjnkFnhWWTcKuq+H0BOD+efYrTrZGV9QI5QhT/rA4Iz/BzV0+1JbvcIiddWS9z
VPMR/fI6NsXeYpQmiGJWFYfMQ4qj2YvvY6fzFPKhzb1T+j9liNlIL5k0Ub7SX6gxunRyxrtDQgvJ
QTqfV8n6jA4Xc1ck/H3rRnIMGhPfKf39ngEb/Pp0L47nBSwWb2A/tL0urt3sZnEJRbWDPvL5umKG
Z9CdkWSOeBpljO7ymQLL+NbYtCZoLq9Rx/vL7siNB7KlGg6rhp9Aj3CVi5GCfCFA7jZnVRtYc2h/
o31xrhvy0YmzCd8XHpKEjUBBGzgZY9CkvWzRvGDMB6lH7nerCqT8RnyLH7LvFyHdS7yYRL9wdF9I
OkQLB73ZtaoGJl6MfwPBrq0hgFgcK87u6qU20qfOq3SO+jRKFg98ss2YEf2kbeC5UR3vSOrGbg7m
KWwUWNzu703+XY7REO3BN2JWz5iAWUFFx+VAlWIUOvT0K+5la0igAgJezSHfE9uOgh7d8ynN+K+y
mfFWwpG6ciJd67GIuygysZrkMraEHz9hJKXiUR+Fw8/3Y4muXfDQ5OiinkOXJw2YIVEB9q3Ty7o4
UohwoFenTd3TN3PQ6gd9KVDr/peL+sKcZ+78s0ybDZ9uC1DNtVWrpMUMbG6dP1sgXtU6Y6drsxcU
2cKePYzHAdSrNup35IEmWodsFUnw+vKDg2wy7ENyq0q4+11klPZSRxe36XMLdBFz/UziWDVeW//R
g+MKSyI47x+/JC8VRBUje02DGb1hTB4onwx2QQjZhulBRc59JTYTC6ZxnL2TvZIrBjOYqNT/XLUP
xVrndoFdlLGvmrzDqZNPnk1SYQ8NIlm+n7xXkp88Rhzv61WqV/Fbn6hqc5BQ1pmAx6Tzw1BTF3G7
nwo/owimQasE3YierEhsYsQAo4jb0nlddCxwgfZEjXTbJV7vYSzVWfkopP/0qPg3tcfz7pztYzY7
1S0MVgbx2Itke4SrCffNXAAToLkWKrSAPa4vzQtSIb+B76L8fZ/z0j8lz00EhVU0rhcGaf80ZuWT
D+P4jPBACSJJXdViC8Opo8ViL+KOTv+mY6BXuZj8Y4/7qPdDBMrT/mehzAgfYdNUD92gzbTcebTw
An0XM4Ra7Y1++oRq1B7E0mrWx1fUyLd4OkGPGTVtEn2dr1QIjZt5wXPwDYxYOk4HNEoCZMkElzdn
7qn43z8c6hEBdcfQQUfrACejjMsBJO/KOMqOeY/oPzTqgKV3+6qsy8j0Bzn4KWM1CCcefkhKss2T
1hl0BUBm3cUWXoQ8aaRAwLPhBtmyg3qqcXgvjI+SVtspdbmKz6xIihXUiXpDmeq4DhrkORb3X5CZ
sc99R5vUhlOCojrrrU/ZmtwmVcxKsXDSkYYTyGLah4AFZS1NtLVK3HZgX45ghyHQOo76IhxIv/jm
leGCc6pKyqfPOlg2S0w3CWiaiVqWHHSAkWMzzbOlXKyh38hEkqqW5fiNE2HeUWMW+oP4EeMZqmy/
YysWo4sPUY4f5ceaqeJxhTymbbslPOAA6YisjgMB4mdlDB972u7nRnzgiOngn+nbYdpojmK6H6N3
KOBA/nu4ZH87k/KsR6MPe5YqS3xsyj3KsNGslA6Mzx5t0oEW8g9UndyRvKh0OaRzurxPw5QBeRCU
/SQt7p4eKiFiUneZt0g6Gzo0rqmH0bXtcDFJXact8KvVdX6m9G0ttdEWBz4gEkmLWIfLPIUrFD87
yhEmCxVD3t4ZvVajde6iTuSuQqNRPhKytjgju69x6vWXJliNclYAMeT95h45U6iNQtE20GyZ6xs7
6sfunstHuFnbiN5oqk2WLa3EB/oct6V632D4zSDRVnnpJYgit2tMANBVIwlfDZbLKn8tFrf5+7cR
58/GhQM57Lo+IWjD+8+IrgwqTRwQvtz6ghYsG9nNEuXlZ7kYwf/xi7BqC/xK+AhZMY+RrdWjQ8/t
Ab+E8E1TR3Ns4cCBM4LVB4PRpA4dtZLnla2h/kEmWmaAFiqp5TosD1zdw0OEqaz/kpdW/+El9YMX
Ye47W6DKk43DLMLup3yPa6EHe14p8FEZGy/BWehIOlPlZ6yd6GWnp0JeQBiqXfLwUWr1F+Z9w6JF
rt9kwpci0FqivzOipvVtKAifZJMbxLskUNsCsRFFKSEhL8roK5fvpYJ52teitCMlbwBuYZ5dyJOp
z+luQpu7SwShf87anhlWzBHT0qjym84a5RF+AyUh/wHmxgzf9iaoXLxQZjcjfIbJMsl+u/HMap/A
0+kK+JrgmnhrU1unk3R56N/M7kyF7yE4F/nOTytdeVwehH/YEpN+dGoSlkK6J/G7B0V2B8m5kwYW
+DFaFreLD16ShMyaxbpjhyQcLRpNKQk2lKA++GtrOe2b5+gl0s/MgE0ezfy3PBGYVXWrCOgQTgDO
45qP0Qy0wS7ReWqeG1g3MI7AQbkR3SqqOngNCQPhFA4v3CZxjwB1FU0xs9YLIZEsW7NlFrKbMuRZ
X++H3KobIctbRrAj2Naif00yAXKQvQdesk/YS3bazFCM5B45PsdDRoiPmzP7Z83wpBS0HUFaG3fx
TSf2mJSdftHrTJoRo6tRKGrob1uwBydzugeaPmhy+oVGM16EjnloWGgecCjBZI99tWcBqk02tEHR
UE/Vso27tWdZt+xhWgPZU7jVVnDxWyG65UNcz/2YV77zfdOtjenK9qN8+AJMzsNWba1GuWG4tXeK
VMbrsG9OArQ1CqoCPLUdsGjOSVs8trHIvzkMEScEUPlEw498u10nw+6fBkUeAZrFXUQ23YU28Bis
c1LHVCyNwSSh5eqgQMFFX0uBHkjhQP9u61AhlcG7Uw2FYqX3IdiTynwWW6rvHPzxh2lk6IqNfL1O
CGx2Uh1Hedju2C3HiJyX7iT9LfeJD5J/0boGgeWMxqz95A39sOFreNe0eiP/rqYW3ENy9SIql9ta
dTUszaTsEfA+ZVXkfiW7bzbTzEJt/po0iZmhu4me2N/GC3xfWGhlwFdfFWe6bslJ7dsDmrjz62dU
Wx7X0NyzM8mwCqsqlBV6A1nB4sep+Te00VvDEEYj/tboYRXD4UBBx/LH3BMD/XcLr0cMJ+5ul7P0
ICU2cZA+dLb+vdXf86P+v1fOmv4HBAJ6+EI2T9rzCrLbNeEI8yIRj1q7zcsZilZxF7GUwdJOAR0I
bgbc0ju47R5I9J15w3AbknW1GfE2b38tqmwPTduVG+047BGpvpiQ4Xq9Mwx3oHq1INx4HmLa/7IV
vKDX3u214FarojucFv36vU6hJl0ALTPLt+6Rq1DJNkxwqvBbrhmCrl0NeHb+NVu2OvdtueNqLhSD
18lxUqkmTviDiLCZScfy9BiUcmOgU4T5sEHTrnpL7mLv9DFW9Iq+d/XyHplRqRwVHIHqh4otDMwK
40V0OoCHzS8TxrHzlphFyHzUMNqJLBndYxDQRZhdaNIN82LzrKB6xKO2FokUi5Jo+ugodfy3jOwa
QUp+Ih+GJ0+3XV+QD3PmNKAuyhxMDoXGCSeQVP6upw+NeO/yL6JnnbSNrn+7sZH2x4Gs0ZMgNSq4
ON8F5tHG5fHKgu3ulSdE0xpfMa/NBnN0thCMgHj7ZFFwS2FokSD12I2M3zxbp5/9N5UEUyAYRBAi
wK+UocOQtUrp39FYzfXYy9BVgCf7LqTbrrpzzT5u3qndXv3v9EhSBHCjyJyhO7NE5M7fbG0B6GYy
8UcLBPg53X74Ys2y0DBU/E6lvb4iQxG9uKFZFiD9ub1qT7h+vep4onpPqpwqm7pu7pTtV3nAytWd
1/05X9gMRwodfn7zl3ZnRDTCT3gJQ4jXJMshEf8Ea4q+57DVyalUAPaaXNshzP0DXGSjCKI75+pD
uaHrbUliuvxqWM2swqQGHHwwUoDqlWjLBGsmeM9GYY+a5H0K7d5fEcLOvzkyiV5VZFsMVMNNjpWi
5yEyo8YaY5QyyMSsWHP9umGmbiwLvjbGFzTJnLheC2kTLh/Z8pPUmwELSrnn8J1V9r7nIA2yq24t
WOjEqiqbQI1fEadzm7pRBJWUvh3w6EjxVcJ5uGvTJ/xDmzzl+C1PPkZ6U8xOI05AUJALbszvdCaq
OBC4UibOItNvexW70oYiBWqAjG3BcRiVDsYzCq4qpLTfcj3d++kSaJyP1QObAFnbStgA4GXLKoQQ
1Tj6+r4bWp3+VTMU32ho/dM1IuclvDTRTY1oV0Q8l/bwCjkzFlPw8/OP5KTafyngp7/GtfLxyWNQ
Va5XtqtK+RcL3FmUZfAbfFSrZ2ABjL/r+DPxbFUsD7EzB3KwQZ38YwSkzcCkJd3GqSr8x9NVPzrs
KzVL4OHerOq9b6Ip1x5FkiHn6Lf3lzJvMgrhZg7xnnNrZ1LZ1YCv0mZ3dPAeVtSZVvPrBtTFipp1
lGdBmkxpV633ggt+06N+UFCACcuj07jhpO39bbPgyTYYr34rLv86gNosusRsDpV9ERonYuyZVT2L
8627kjVz1M1UpCc9YMthsuOV/htTeB7zFL+tYUXOaeGMy/nD/SaBEdsOE15gJcQuPg6HvffqUa/p
i9wQL/h9Yec2a/iCMP0gBfI1IAoFrdsZyv+YYOYoemUjKNFGRHv9/FFxcWrM0c7FtpMRZkuZSrIK
aC3ffa+eMhXF7hRilk/DL/5mfCeNIRV/vRm4lvC9LjE9gslVs5NaGtDp3xd7d9VdepKKqnVfhTzj
D4j5cDP//wVr9/phT+xFU5BCXhcBWoAiDzaoxUlryj7BHjEu+ct/111kZP3W2X8VJ91AdJSrzCA8
enMs3S09v10mZjI2nrriOmFAKTM470dzGCaVAKHpuK8BG7MKykh28bEvOxTQh/LbQhbG2MmF5nol
X09JoTvaXyz7suMlnrqtaDJ07ghlsfRZGeekvtMPvR1KsIV85yFw2Ro0bJiqwYjwxDHca8/C0WfW
i4T/a/dNgeT8AQy3/ZuhBEjX06sSIEKUMYINLHt/qZzqVWyo//3GzTnrqOm3MDWPw8Dv233NvimE
hFBrcIe7fWdOd/xWDMoR7OZ+bh83sGwfKEVJKQBpF2gFvc2c4W4lH0HQY0LoPADO2YraN73Id9Oq
Br1SA1VeZqnwNLKatUbuAiyKDky1Epo/S8HIY5KIbyiQHFnf7o2QVm2ptBjJtZmvZClOuBUlsIeM
+UcLGU2t8ldYdc3krutkHoh774tdamHHGrzNUlHtVffx5u3VdhvG3ewh5vOfktG7gAOK8HbYgT+U
W5fx9IloOwxF9n/2r3UFDjkAXEVm4qvbetFnIn7O3DsIRhhcSH9zGPLc+uM+a6KHcrDxGOACNirK
51TL+fRq8tQ/wRlWMeY1wHS0FBaQvr+FM81ubRuD66gwlR60vg1PenTM/7uVELd+pG9adKFbjiXb
nJmzXROWRFFUIPPq+X5o7B2dYnL+/gYYaTeUvk0aLB978EVD6+EJcugtSEEMbPysOfE/8Yb9ronE
VVab265ykstchM0ttHNccsrBOlzEctULWGDNRr4zVgbbcOcttgrI0VcUN7TlX8NMhPkbOB4Rm722
8k6dtS5c8Lap1tVqK6njPMsvVspcNBqrqTujrk3T89/bGHqM927abhFId4P0jBobPEpsdw1y+Mm/
Xd4CA6iJtycxCaDM3jT1+Hroc+Vszdxy+00b9qFN/l2kP7uyIkMSkL7GAREMZBZrJgQqWwsaq+JO
LnLQhlj+PbD9dzB1QfmfR/HALQh2FosUrgMAykvoEwAAyr1Xs4NDVusZiRiecK2N0cYNn9uiflnH
awf7rpWTziHGpwHVVAihjESrqWx2QwbP2oujvrnRCSBGD1A5v7Wk1kzUImHPvmYSwOxvrNWDUQXv
RftSj02EUu+aUHvFiM7Ww9fvQEnbtADs2W5dje2ANh4FuOzbCOcGHJfld4fgLqi+tuUw8pgUyieM
p35VwKcC/Y5R7tEJhsZSFpsnHtkc6LrgxLUvTBbE9Xsnf4KqvO1+hWQwlNumgPL2t4L1wG09Z2bV
CsM/Oc6UaqSDZORBV08iellTptWVaXw7tGE9Ih7vFdXehiiVy5LJO3mkQ8//ITn0+ESetFva5tgx
YSfYQxcuKx1W8AKJaq00qoh90RCZt0CWqGh9/3ODlBNa9QqUX5g1m7gB9nR7Y/lyu9iuf+Y8b5Qp
OBHo3dP1qsuBCXhlY0+7diVuqoBpmqpyFJ4RrDJ692GZMykTfXcLaVlKfQPXmzgQUwmk+y5vtBB4
n9lG4yulAvBdqS8MI/dHFrgjNjltL7c2SliFhErAQ6y9PFT79PMa5cm9XsQ3hoNLQkZWOg8hHKvu
i3cChAJ49eagZMv4pEAJngNWnHQyqe6DMmY5F6J2XHOyKWPe+lGdtHeyr9a8zzLFWyuKikrBhj3x
nfE4PZ7Bp4Sih5xwd3tG7a9oE5k6llAFStDJRxcC6Gi/IoUaUZb9NQcvTgNMuXTEvQI11Df5FgNQ
ml6+kLL0i3ZKSspxQXopBHCD2wIEul1bP0JG18aTZmu09qORYX9RA48h0tBuYfCLaZRdRjvfMzUY
gchq0w0T066qoaqwbTOFWuW29loRCTjD/N9OELWOyQg1sdVg0VS75aSeVRh8ZYaM+opkgYqWRRoR
+PLmzVypn5IUDfkysmql54lcNWJcpnlLPZoy5gOfU+AAANrGvVCJgV2MjLh/OuR0kNCIvDmBd+eW
iU9lTuZrzr0T6UaUNJEJyVg/Vo3yQlwlWZtN0QfwleFo8tP+WlQicOwEqk2lZKamgN4l7iqBluYG
Jc8DpR3uMl+AYJtsLCpK492JJP7htcqtlOw+xxE4V8fbo5h4ur2rRu8XiZn0YMIzr+8s1zOON/MZ
pJlVQloa1gRO0JZNKrQ39Qd5XtuzqeujbPAlPH5T1+OYgGCdc1WmIqIlCZPxpN/tmzpmd4GAlV0+
BpjEAokvNw70dl2MjrsXxJq6QqYKDsxDrTHkrcgkKfn9PIruUf6z+iBlH9CscofpLcbCip9EXNWA
JtpH11R/hO9zfUjWEPhub6mz7RdfK3NuibvWlN885SGz3Au5lfwDKwEUlZD6ArGGlb4kZfMcrbyg
3lUHGYyxpKCzUuf0PNZHRj9AG6i89GLavr695tx+pCv1UIuKy506FLaOzAJ8oazck6G0vf0AV+uc
2fLos0CRoeaRVnH6ty+lJ8GVIXIWsVDSqbfZGu+2/v4mWkjsalKxeLJG5HT/fPf5jih7/eBruobJ
0akRawSFfV6kT11CxqoT0eppJBBvkUR7sHlLIcZCb/Z8/iBkDrH9mqisTtQ8H2m1K2HAjkArIMEX
aA35TkQ2oITckFx7WDNU6pWtNXUk/ZjoJscEsnNH6hl1o7IuE2AUe3k54f5t/xxG1BKMVSCoqtEZ
w3VhGjxvHRf4lJv3x85GRG0QZ+wQsq99TWpzIedUKFUI8MZf2+khnn0AuBg6qsq85SS8EduBxz8i
H07+gadoMWAF5zxw1vLsvs/y4jcGiJoCqKVRdh4/Cqoi8/eTIffrN0mfe1YSkXRZdtrG6676zAeN
NroqvZjYaEgohbolCVdfhGoGJ3PyUtGEuafjN8oTmaW4zTDQmC8AO8FPgCwvCmhc12FTfMgnG6V1
sr4Vw20IL+TT2WHicPWG3nkQEm8iF9wcsTyGLRbRijJBTEZFKwjh/y8n9DS9uTvBQP7EhMdnBz1k
icGfSglY3/NIgrGCrI1Fd7rJbIi++9DeoLwQgU1iYgbvCmjLGCNM2BzamJGbhez6noLC8GxwLzf4
CUCeMZJ2lGhbAhzvYELjg1D5SMd62vBXN9uc6VpDGipEGci9UeKSTMAxOmPVgFFfahcGjhex8kQw
gLRmyyjuIqu99unAKNUJRNOhhcP9pP4rXo1/v+13JCkAFZ/EACbKEkHWJBWnsx9y8EtToWV347f0
78wfLFUObhrk30eLXj5zVpynj/7py1oc1qkODUAfBEWlBuMWuUkSoBjfO7GxRwp9oNe22z3p6Vva
K+ZnNnaAvj/yD6SxNHLuQ5vz28TK1B61RKcSs2SClY6ToirAa6gpFbgZjqB0+k3wOqjOrHvAYdSE
pGELNwLT1sCB4CnNiGr1z+XcgU+vrsZ+/OFG6hqDcSLutRwM1Wt0X9BXYwL7VVnNLYf+H0IaFgiF
EQJbm7I+GzSAO107BaD76giz9ea1r3Rk4BvnG/hZfEaiJXk58OgR0XvAXwqc2nSZL5Nu2bNazLlP
NOGee3FpaG0iMrZsdu4H2jjwDhGYUREN4Gpkw5vRyBbiYih1nJGJ7F6QOjNMkvDk2nOBr4baWA/D
9uQMkemWae7yvVoEufPLg2gkRrdLRogMPd2QFQ1fhLXIK8I4TgYV/RoscqZOXoYgpbXLBj72A+d5
mXIwgQydvZxInufDD2ZXKgCvqElLv286DSynuibBvlJYtVvVvSWGf45ED+vzeIW2oRLIxJ9oFiu5
up9d0Eh49PBwQZ5+6iRc01I1rL3F86HzQEqSj9bE9OhSAwGPXFRA76VcxleAy/7d1HlnquPdGaLx
0BzfQJCuLAz7nVtbarEoSS0ibUJepcoeSsrYFwkJh4VAbld2JU4z8IX0o2NixkhIq4qmrxr6XRir
kC1bCDuT1qsq3g/JkCkw4YlTwPHdbQzic4AnBToNIEekXy0ukwuIHS1mL6QN31yq3SM0jUBXkzl8
sXGCzLKufn8chxm8Cpe3CgckaFYfnkupdC4BxHZzyklK3iP5CUvcX/pX34Vo5dxTB9bg4MC9X0vZ
up6W611HX1Mwtc5MwGPrmPODt6OMRTdP7Gw0L9c2wsB7yWm84cb83iO5+54zNvnsvVqlsjoVzZBm
4GGe+Zffd6RPW5ZdwtoJ0wKSS8Cx9Hc19ojOpjK3m3cYm82msKH6+Zw3veFiH7kxOKv4H5GWVogj
rgob/vnp4L9nFexZDxW+nrKjpDC/XgFNIjZm/f6yA6JdfCCM0CEfkoHRRDUTriLRzmNJ3nts3aqy
Osdl9tpvaTxfPp2re0wrfQrqL25GulyaimOpDIQThOIkAxJphDunPkDde7LS9j+9X2EpRf1oF/iC
cblSSuMx7a/51VWNAL+YDxh340NKCFcoT/NLzEhGUnIqKVHdtWpQGskQN0+EiLEtbCDjcZBPofok
CPpHToOtIO0AwyVOoswlS7EoVyte4RVxxAU4pMv/iae0fqHsML+4Ulgw69GfwDDZOoI+KIxb7P66
mnA+sQO9qT2yTMHxP9C/CO9e6GyLlRTXPDxMuK2ptEPBk6SgY3Ml4qqB6sBqyU/a+qGrNvKbZjTU
/ThE6bDdu3EMIKUHUiONoxmhIcxU5+97cvMMIbRW/s1LaAQTujAznJ3POJlTj3hA3qErog38fVrr
yUhBLhIS9IDGvkVpphCPtjfeeBHiutoTxT3ka07qA1+G7pUeYdb0dHWzIbj83k5Wlsx4dk4VxnL1
9BLk/byMycfOpxuH3VdgeuTbgUNPwQPLR4zB2T7UCK7v2Vxec2+aF8PfmDC56bQd4Rytkib8ELFm
9DfxEZWvsnphOY7Alq9MJyOmLyOxEKjIbFQ5nvMgWYTA99hiMCPdSJ+CYp7aqUeXq5kMWhx9vuvs
dPnStsrRA6OscBvhqM5474Tz5UH8jDY7zQwrk093PDUOv+L3R9f6nqFXlO6kULFulcwRexHUvxPn
vYVOeAZYfI/+U1luZ42B9KdAtpmgIZJAyjA6NuiB7zbWZ9zD0D8+EFi6bVGwwZXgCM/x19qToChk
uW0AX04tFHBVl/a1y7hbVcmBpVho2z9ZFxETUg+BU2CRNyaJdbQtmQai6+vMsxuB06lW7myhmVoP
FcBkksVBvpFPJFsedMOiYgIhDJCArC8q3uPa/VqP775DpNGxdLZ5abAqNF/MhufHFB8E0CfaWXKS
t+u086z8dkxeWG/iL63+9E6F562lyTjdIMAp2oOzBuFR3nmAbBX5Eb6A+PSKz891HGqOC66jOdyf
5ruDHc74hb8rLZG3+6JjvW6J3x3SmBbpncxpI1tx5rtnH4gAOCMf/Yrv1GLJEw/lzTumqqxC0Tom
5malC3zvrt3bcKnZE4KXOP/GBedAlWKrN9FzCoNcNEEp7amleYKjkX5xB9nDG0fxdyO9j4fbXrlf
LPXb7vBky6lp+hdNAB6ABErNyqsSzDI4ICsbYaggefGCh7m998UA8m2ISxfxRiDqpkgF2qjSY6c/
13zyXmcokKzm41J5ULa17M5Yku3LVgzfI/B2VPaGYi6oGgrxKKPkOBrkbewAGL8B1i+HKGhmspXT
TSouS2uL7OPSnpLd3Ydxjn5Th8ptEhzdr706wy3odeO02EwZLQWOZtkIwhNxQ09RxHyuwbebpdMv
hOcKwEGvTTWq6ylIA5Rri7e2tca7h2juCdAdMrrOTswS2iFiJYVUaTpXsjC8XldPG7f+FdCa89Tc
RR2ohCfNxDYa9z8uGTi/lth9bbPqk5LT6Mv3dudAjc26MCx/etQHSaE2XxT1qDDJsuPT/I4fZX++
d69ppHuwgw94EP3PKyIJpYJp1ylKjM1NrphU22xS2863CpqQKVJyKfjAqzwlGTX7+qnpfihtgbJb
b8ggKrvANKyMCVPZbnj+bplCQMqC5pIDk+nl0eBn0pzQfcxztcWRTVuxif7U2x5rr7t3xxFxKzI5
vpbJlDmmti/GCjSqMXCTTxTn5/kg4vEbuqyOJ4cxIAtRmrVK7lEcpUkuzvfZ7NYi2M9SMTPq1ShU
/akQ6BcUEpM+5mMWPYkLQydh0PHJ7FhfqV14SvVBxy3s+688ygb5v/Cbgif8Fgsr8Eew886HpZCe
Ak9sAbeIyFZK08bJddbPsuqDTJPWN73/aVgaAW2ZRtn8pDYoRNH2u27EaIc6h6yMKlpBPEYMBeUe
TbjoV8e5froFJV1f6L683+6tSo1HlndeXFDZcPr5f6jFqNMRICGxEAUbCr2g80tHaD47SaSn3pEP
opzF7qttQyFlx8tOEuk3G+WAV8mYvuFnic0jy3sYslxuitPEBnO0bEkBzay2riTarFc/yuBi8BCw
npVhJDlPsKPhR9W6ntbUcUDDtBg4donAaoDEOVdP8sR1CJfhmI3GiWDMjLM2WSR1ZeOF4FX/H0f0
aGnZuiJlcxRwLOeNowQQMPHrOelDBxTjtIZo/vQ9alDV/sd1og5fGX5hOb72qKgOLN3Uj9q+2vEq
aye0On3GlJa1/X/ZNCB/eG6xMfg3IpFeh/jV6MIFBAdcS/ILS0ycAjr8SivJAbzGi48RGTBA9XcB
GaLhExgHcgcg4u6CoOKVRY6QDD4S1JkBPyxsf0TU0rmMjnm+9NwPuK61/cNLas75rSs8p3t99lYe
6WsoWjuyRHtP1LNz8+N3E8F4vz+JjlU0fkzo+0eo8Rjzpmnejs9FUE9J7eCSCVXZ/MQ/yCHZax1b
TbKbYe5uxP57pAFk6OM0qHAT3Z1ycxXVOCoQkQlhL5Kam3wRWiQ5hVZ1qJkJrtHx23LoZLXKsBBz
q3jYVy9pe1Cp6Eq+VOqMMsmEjVKMh6edOnJ5gtMSj0+n4eI8hpkN68w46zuK7DpfoC4AdWXcV8TU
m2o8Nj30pz7j2APZhsW1e69ZpzKTDV98gynMrB5rEI2xyYHCebe4H81jsLDCOXO/ry+TlG6uM8py
bvvwyQJohOwyMipHNqzKfm1/rfqwUS13DmZCbm9koP4GYZkJdo9uxUgtNC8Sna5G8w6amyp+DeWp
R3TlHr0OcrW4cV854BbGSpmqe7lE7rbRwwXDBbMFbMa1fskz1Uy+7dMoZCQoKhEP6Csgxed6MBJi
CzCRP41t+gsDIT2u45AN5zbZNqMFq6ffqrshTDslMHi3Tgh5nhyGL4/Ct7SuRlfMTYUdmc5w+rtF
Cb9+Y5wFHG9Qs071IyQcIp4S1EI3AlAdDjl1bozk4gSmgF2RYIubw4lMQ2UdjrMXvbXgNwFb7SUW
D3iItaIXvPTifhAXBkIT8RqRXQW8uAUzmCzJzmevuXBhlwuulw0ygBO0jz5u9dJ8ATi9y7ZZ9rcr
IX6XTy8feEXUn9bJG1cEb2d/mWuYOHMdpbqMKucWX6FhcYI/iA563MYZHlUf+R2DPTyy86oZtthv
+ZWpM7RtfgKWGD2aAgmPRmX3igYFPRv28iPUcFNoZqCa/A5ajuipdcPqad5PTzX+aaU8ZMadbrWm
u6GpCCkrwbc874Mzie4ky/s5od7ynpQNUqIilYqJUiUMECHysbSsqh+ofQwYrbGM+u586x7IkJVn
fde6THEdQGuhioJesv6+RnWgjd0fVhn0T2hEO4r1lM/aTqB1cLeoc2t3hiNa3nExdSSIWb1BKfAE
sj9ZxUtGY28c5Brv65lP9d7/+036KCmgRpFWd2azGwBHri1K/j6sakcFegXH+ucSlDReItLxXDGB
SU8Hp3epEJlo5YwVm3EHri0rfAfzZK6tfUw7tG9zn9HJUZAKT0quERzxY6PaOvjHarkPl85VboP8
OK43ZX+vm9L4Fqhgu/qxrdT3IwtfvFI/1pRm4jkIkHAgnzBloPS0rJYc1fDqbvWfRgibfYB26qye
Mw0XMpB7+M7ifjppQ0/bhQ3l5SjygvcVt/wtIA2+ktdLIcmFdZUdKpQNEuARqZTCdagX42YelCQM
8OIXD/jTRRrpZ8qewttbyM1QwXfkAUGjqiDYcMlIHKqX0kJ1rac3mq8Gi98ttOv5z2qxtrxfTrIi
aIPw1V6/Ss9gg1pw/52KEJNvZkL9UxTszwxR5GIqSDdXhExiRXYBGQncJzu2R5vJhlPi83zDRnKB
APHlsf6gwzsE/xrVurLDY/dTeQfIGAeZPUVi6hoO9y17cgZa5Vm1aacpdgb5Vi5Z0GtrG1bbf+tj
5sIbHQQyl6rx81yK76EIfPElA5yjTM2TWq5ZP7nEUr58dWZm6COgwHHEhJvZFAQyiCa3TBrtdJIm
Xz86A4wYVUKTorcZexj75/cov756YQifMExvjr0pCG08KCgiB5V4+6ikDMIhrueotLV36ZuBwFgd
cwXFGajWUwaKLMnkOuTJoGSiI/ChCuj+J7W80PugvLvxD0HWC983D5rL4RwAeSAv/hjys5sEEqOV
yjVPwXO8pBWzNPsdXHKkFMeoFqL6NtDp+qa+qFrKitwJsBpwi9CoGutqqFxho4lhV7Jm8XM/Plls
2MM5/ugSMANAAmoYPYaY4gJ1uirHpxHdHQ7w7y0jvLTd7WrMNRxFFnDmI7Pi4EL+oWNyAMSDUrcR
D4YolnXuvFL6NftPmo/64lw/DAPMt34+JwNIDHK5xv5Ej0RJKCrd0Th+T+KfM5hG4yQ5DapnbmH6
PnRrxM8IZ+xgzpGZRnbuQcCXAIZnhGunzt28Z3LiS94O5y09bgXbZA8DYPEED0ayk+WXpM1+ixx3
qhdMZBO5KuT0QabdMAxIiKYQ7GdnKKqBs9rD5ImOU2lH5S/3zzgmAso7KygKflwuxeZtEucY2u2N
zufkyuvZMCbaL6VJaO75TT4TsBedjTPbqImnQlm0KOKJ4U5GpU650w0EW4B3Nyk7LNW6ZuHRRKje
+mOCOW9CCm1VbHoJlYntXvmGj1EJ/8SuV4Pslq2rgylzEuNDHPX6OfUk8ROXVubzLQpZC9ogWSgu
NVyuxOI1Kog2pyQht+yFGkreOu+aBZS1tuQvmNMQfxg6PMwBu32FLpo56U59V3gRJ331PTLT8lEx
GQtTW2auwKNNH1Zim3ET5R6Q60XaMoFxxcR4sWcSrTAd6n5vDnbCuCh146Kgi7SPDOIsLcFp/1M9
5V7MaINFVhuUckkZhERDHYbiVFCf9BMBQL019Y2fmz0/0RiPZRgibI/OH2rqtgrlJGpwEXGFXwZz
I8eEg0WcvpKLHBQGwvyhNByKBKVIoOOg+nnVybmIkB7aSA+tXoxgy6QXr19gFM8m4jJsVAIRKU8p
Zc2iz3I0kK6y6/SZ41d9SywAfe7dxsvYGIKeRjrJr/4JjiX3Iw262QSsOAvaGzWIHMsu2s6gfdf3
ZRQIhU4A52lt34hUnt0x7rT2/9TKpisoYWMZqoT20keALvM5nVszAIJaM4ZPaqhyBX70jOhfkCJN
QKS6PJKbrxFNH+QqqB5VZ+eBFsjfTHIAw05UOh7vjXyxQ9lYpq79/z6UqKX3EMEb0q/sYF9Hlb7e
X5Pe13p8Qq0slSZF2Jl7ViadyOpMiuddmcantSXfLry8eaLzcwqmOdTmuqQgO2CjB8+4QzHJiOSi
mwLewLKhkoksrnACUSy+QpYQOtCm47NX4NKtURw1H5wEaNwAiBUu+6ax55KP8JtrMLMOIyVXwxCZ
j8POQVuErTwBRcfTFk3OM7W8/Ks7EfqBkYoCZ5G+b/ywLo41+h6O+xOIuHU1E8u/cRzejCrU+X+p
0Wt6/9Ggx0EK5EDsepMiRmrrKcThrTDBlfvgShuopvi0o0gkExWMtZIJEXCtOQLpezs3nyBfW917
w1rzfuYpmIvoJlbKSXhhZwXjyw9CjlL8eoZdMWhIfYXMmlYpogYNG8wGLvSsqm3N2QAYzdZ+1S74
w+FUTVf+Y/gFr5lhj8JsmJTERDpcxZL80wt/Es2JnIM8iD2LvyDHLaOaRWmCnVJtKgjKpejSI8Tf
mzIN6GN65PORawxNqH9ubeF2gqqWN6IAtlVlP++Kif/dYzYP9g9YaCKy3knJxzTDNDqmgbFv3AEF
tm5aZ/efUuLh+KYe7BOKvLIwIervQKwW7Q6nLZPrHXx79lJ9IV6EYKcJ/KTDB/iH6CBaS2wuX6wX
vVRti26aA3HbZAExtpBL+20giEseWOIPOEOiSzpywCvzm4fMH7UhoZ735uqq1GN+oxcs/9BopXDS
gHPJY0NII2qkOr6QJZHz0+by+agXJqNQQfQWNt7woYahtGtxovE6ozNpBMltaRAlXthJZAyXSCi6
SwcTlc0Z9zZEuiZ0IcfNhBd14FKvmw/K7RYlKBqXxL28yTYb0ydaOSX4V666VFQv62NA1Ps2iMy/
qj9Ntg+7GFwq3Isit+ENfWcStH8Dr1BHV2NPJOfP/d6FRcu94aXPvcKLkj0LiUovAJ3/m58FTigJ
tL8wSf2u0A37AtPr1KQpx342ubAjEmfkdAGh4XZnuz2NQe5j9XruR0/afOibat6T7mHhXuV7YRS4
iKDr4g8UPbINQ/1NM9G8RG1tcc91MyOI6RKtIxikW78pAa5yZ0wnUWbnlKbKgIkYSS/QJZy/EwlU
wCpNPyr0oaKpfAtdLyCfmIGuTkhYYqKpOUVQ/m4a0MF/pM21dJvOAUjkFl0Br0jJgx7KwqqbmBo2
1pYOX9n9J5bKfv+bc+MZ1vwREiUMaDw5FI0WO/eef1sH8VnGeIkYoNJ/AT8WqAJ1Ysh/BR7fmqyQ
jykSQQTiX06iK31tbE9UNkCs3iCTL3zTWCUateoqTkrkmm6KqsabsRWqk/qRdur5S3/A2X4WGTfB
nlVQKn4IaS0rwNlcOVbV223++nktu34S9XB7HYYtuGWSPXMa9/z21o+XXC06/WsYwfJARXWfRxeb
pZW8U7akkAEblNEiwMpPHyxGJmWWBBcBLfFP6XwuV93P17hlMWIAcMJ5lwlQMIR3ts+8OvrkXQqI
gO71XYDWIY0qbZUoh6GHvCfonm266WIgtbJ78/Hkd2p6EA9BsBpTSgxBXR1uVK4bbNGgi6/trDOX
zCx9I6nv5XXtEPt0lUeReG2LJcKwT60qoHETcj9jadpZC/arGVtiHGMW6EsLb5wj8m/g+m1HMXP1
fK78tItDYCpD+VfQD8I+r3iaVYhKGCH3t3opMRKw2iSeOdMrefJ9d6FQbiIz0HXeskRhpH7xDhSG
ZnWwtqPO/VkRYlbmaCcpKfbwT+v3WcwkxCgh7tBl5jYVxeOjoU8iMNGEaMXuwR3TIZkzEaY1B8ru
wabQ4zIdL8qY/DHwKMT1VeP4ViU9sBLMOY2rIzaOtldWeRlbRSoUpNZC3rebbT113kWHIg2KdkX/
7D3i6lKBC8O/Tc/fDO+utyzc8lznlLFfuXwKL9P8QUM3zhfYO+s9saL57t+SKzGD04usGGXvsuzu
lbC4pvr2ZCl507ztFE3xHugNQY7TGqeYlmW9Vxdmqpg/mzAgA0xzJz/T9nptMr2kc8U8i1In7/MC
mTBjO6sTXFWe8HZQllQUB1DFQ0yesGsW/MjVGzgayb8Lu8hFy3rurFNBayekDL24mIfUicnNi5+m
gDStswj1Ss6adYXvhWC5gpqdFDP+LrgHGdhmQfY+V3baAyzVXwTLCp3XpyK+Q1HeAApUonZL79wS
6vxFkjr8n97MFONv5HIC8t67Wa0CTr5sKEgol/Q1GOmwA1Earb2+jCM2Q3NsXneDPaCHuiufVM/u
Udj/i4AXj6veimDZjX3SLSdZDuBT/sGlsV377Y1FGJrJFQo+Aq0wSz2DC/xG9z2ZbFrhEAdIOf6R
bidrqlw5obiBvs3PjO+L4NJgNUJ6ZR5X4SJRWrWjsk//GoEfpg0s97A17Sa0VZEWQZlWRHeMRMDL
U6dGob41ctlHu4Mip5LPOulvFBLO+41InF3rKLHf8/xNk5oxIElQiWKIkVG99oD1TWO1nHef700e
q2oy2kYjH2kLqH5sC1qdoEor5OI4TyF42ibqEqkn8K9VvI0okhCC6J0kCXq4RKsirjrji5vJk81n
SZerarG9/FU0P94fKZh6fmwwECT3HN1FXKIGS08gOw72TOp39BKX8Gj/xZMvIL+CgdzmodNFCRh/
+wuBNqUKaj7v52EgTRHOhpXIqblQlDMT+tLtzQzZkuxol3a7upe3FF3HO8WVHvLpB3wquN/dosyI
6uJUL/FVgO4P9uqAXG7KqwcDFulHjoSgqSNnja+4jAABLMHFDP0CtHQdcweca99mssd9DtgBXe+2
EtIiYuUtV0fuD2Y6zWxgpsYW94hSUwWeOp4p0c4Zx2SI+q50DGNcvYGZRc/jpoeKWWH70u6Tk2lJ
0qteYzZmSnrW7cWkscQZrwDFkvnM4+xaUxvXYbwLb0MUx5GDRQj7enuCFYoiaYKRkkyYtiDxwJ5H
SJXynmOs7bh0NfcNTcbC9Ik2bRChsYbOaoMRirycNwnkbFXLYboske+5hVoXgohSSkI+B8vWhJuT
7F8WxwcWJVA/4ha1VrZTFTX+dxklSFpf0JMhgAME9hoohaSkxxBiS12cG+XWde1LIABQ2N31vNMi
nHzVQBvd7W7aD/bN1cY5T/kefik6UfpGTtN7BDTttBup4PqYwg7M5hn/8Gzy3Ft/J569y1s7ZB8E
Khe0ju0uPfd6PwMr7U5+Nguvh7hhnXl5kU3NgEHuR7WdY9uTaCpjXLy/LlIQ+GCC22UZ0/hFog5J
tmrmeJdLqsPY3/b0Sey5FOi1zLmeBFrrVnLOP/FEc4PSd10U2qMSTd/iKBgYQHOestHWBTkatLu2
txnKLisQICUu3JhLjMd0aISgeb6TGQFUDRxTCjTmFFBoRP5iIHOU8H0dgp0zVnomJjSRMIMShCSg
n1ynDXu4ygzxKeqWdeH1ZsGS9o8KCTDUaw1rX9ObLOHvcBZlh+ph1LSnQlLbQXpwVjLdiqF24OaT
AoyR7EQLnqRnFjPEk/NEgDaW+aDGL1dcYdvMupSi5CCUczkzb4evbRNE8jQC5BX4SiX1m2taiHyL
Vl/jv8i5riFDMVmNnti3yo90Af8NjvD566ZyWFSFAeBqLAPaOGWCESwHaXdVJlEvhmG8azk0CGbW
fPWUW5BdE+7HrKQ0Ks2D/w7HG+kkNx46NmFK+aqHG0S9PUjiKL1I/Bsi+U5dBDzNeUVudijOZZ8K
MbtgufaSvS8TZvakDx0GLTehFjlXgT0xIUPlvZIXAX85kRFLPmJx2ftYq/fDKUEr8o9ZEF39oVKD
yO1/k7y4ywa9YVTQEChVKODsM+k2CmL4kyGvehiUpGLXBaf+tGp/oRjtJtfnEoKrIh6MDTGbEpbx
ZUSO+3yiKamZNZnOOTSjlp0/vzyHILa8hP5s7zLT8I96WJI7M0C0dWB+4Gqk8olrFTl51+2JzCI0
qhGQtSJM/JH8EDmEAD5FiuG+WFyO2BfQQTywIBEeOzhT77iv9Ps33kLHbSH77FLs0fgtL/pYN1Ni
m9xj3J40fBacFID5D8J9s0I2ZYYHdv27RpZq5qCnZThWxGlz3y4Pv2dHPmWIFx5rsDbG+9SC1bRe
Csu/iGn9cZlmBBxpv9ZkdtmRgPZJO06M7SX9JjaVbzgWkq4hsAFFe+LQbsOGTCDWH1gN5yvaJwYg
T2Vza4XFYlCAcMWIr3+4cnG82eyO+CqTK/U364ZY2jb7NxnA6Al4xANDYgSfxgoZPuBiBpAxHPZu
EvwYeXVrle+jkQ+Cm3kwIGgDqKcTBeosnfw/bjEB2uH/SPx6s/aZDwT77ZY/kYRzqoM+i/4/CKaJ
emrZLvHmr8/FolAHqDIx3FqJSUc7YfFSaty5vX6Vx2gD+py73hYG0Vcjurv9EhhJNPJhD0srowTM
RtpWIrvz0kdZoJv6wL+1dzBnAOF+FU4N4CSO7EMu47OYcX31sDGUOi6/evf2sWj3WAjmetB4LIsS
dYiv8wFr9zusXhq8rP/1qK9MU7uMgNj8wBUcCHWF6pv6rmeP8JspOb603GHexzQW/eKMKq0j+Gd2
qttfQF6WFpPShANGFXNfwW4Jm6JXALXclM+D9M2rrOFJq7ndv0iwrD+s1xYSEOisepKt+BrclklL
dLfoxYRnjTX/VtkzKRb1HvEcNFGuoTFSnwX1e+unv03yICcS+WQ2TBYQbgSU4rz5ePnN32C/Mp7J
dIciQJAieK2kdGT3lnDuLV/XtVkx6giSKlo3YVRSjtMCmx0cBSvG9GEOMfsj2LCqqbVLm6/Q/+rz
FXX4R0bhJ0291m7/znug7cngBW58ZVbAL+nvrGjiCR4XJsdCAAMFsclLmDIN9cMd9LoVQilfqf4q
IdIj/3pvkZfoe6seg+Hsw5bBYP3I11wjHGf1PIHm3vojhhpjgH72JsLF1KF2bYG8byY6Y8tYa4S4
3qgSVLMg5FcpS4xmJO80w/chbonBfPAmjKCEZroWvD1TTcGQYTfZoyRM6l2eAaYQK7brePtsXwtq
63uXob1VlUb+l28SVmoFvE+uZ0dRZOf0viKywhSrHPlBTooQOWUsv9VMhSGTnHGQnzrn9EXnpLe7
uhfBX6XNtP2/I/moC0t4JHPSI6YC7/jOO82dOvttCupOzM3gSm5PsY3QuHtdsDuWTZrHiXzpnc9L
gkw2cBICw4f/0CRoZJ1XzFdDypktt3wZxZd7lijIMEY8CepRni2bkyldmsxsLplhPQri5/9KnoO9
ecwJn9sM/1LUM7XonsbMm3OYB1YPAVyKfugmyMsuuUD6I3y0J/Yk0lgo2bk30J9nnWXTcl7y4zjt
I9MOCHK7sm+IVdU5F91R/EkpcHugyFJ6329P8OQ+YZR/JnkgBr0YYHHEaXVbcUOSdXPzRvblS/gU
ouvap4/yDMrJJWPYFQ5KDYMdpTJze6RFI3oaI4absSdxt7g+v1FtJ6sh1HNjHGc5gOPXhxM4rjEi
E0ZU0rRBx6Bl20ndSIzPRJwLTj92znfqwl2/2mDH5K6YWTacilLOCUxv/KA/yvFHZNEIUpX9ZrEk
6/UmHWZLErZB1olRPkKtT3RK4KOtN00xYSnrUswN+YsLQ0In3aNPBM5E/ZMH8Y7Y7q3Z7Ec4m18t
uRoLg3kJHlUamY8mheZdfMNik+3Y7Ywas0a/nSxCEWICnrj5r2F+pU2nZ5labnzPUfnmtJH/2kWg
FX811kgVsmQKqJ9mf6uvXkM5bt6H7Nu9aybnNwk3Onzxc4f6LqnSab/9WhuUlIcx4KgMJHkxQS4E
8l2F4M7eb9Ocw7DBSJ6s/x20LXaa/Li5vVJYGUtqkM0j/3swNaoQr0TEBR4ifZz5PJne5VKhAeGd
TFf74Wt6OepaLEU6q/C/N3QfamcTUyBVvSmsBxtrBC2sgkhFBbfOYdlNCMEgptPIJp1lOYGX+2BO
JJt68ee1Z8gTlTtfow+ws120MD2uwNrG1kBHBmiGqoNWCpgL+j6R5u+o0pJNVxGmSA+1mqhZ5/if
4pktNPVB1BaBcFlPVNqIg3BWdMgXdNXFLTDDNuufD7xvXJyIklWqIkSiIVHFHsSICkqGCnL6D5LK
XckSsEmQVLCozYtCgCdMAM8jXZyU4Nrn9JGdNA40mTNm4kNi1+WAvcS8DLpxzCUIO/vq8/0aY3Rg
aqU0YrDMnANnKKq0Rx8dW1AQ3WXZE8xLHG3FBi+q+2W9ItBN7CzZIGxsYArINROBaWmmCKw7HXfq
xMd3J58byRWx4OS2ULEjU5pjHkx8bz8LjZFuZxFIyCmofNVirD9faAKGd08ka5GVzlxL1uKg5jlj
gvQol4v+aZ26tCs2PRxyEpzrG0PAF3ru26ZRjOoqn1UCzNeVPKRLe4di2XEDGoL2eNRCxB5IUCBf
rCufwLTbZFSkD7eb/HqIxbTV4Q5lD+4WJx/AE24WmGeXduY0zX4EYWy/050UKafvfdPPJ7/rvEaS
VpLhg0l6MSQW+HGxng1FtUCcN3nukwpzObbi/D/QFk7cm2Nf2O3r8hxWS/GXRYCuIEOu9BvMQbi1
KGK24ZfxPGLcCEOUqSm2OKmwFq5Oticd53eKynNK3X426AR0PQSSVd54VIt1LiulAkvAidGQ/ji+
f8SgEKCXtSI05+GqpKoaagHZV6XhML+jIxau2E4Q5ot8K1fvEkE5m6goCcyGWNisMjtG0Zhsin6t
dikYJYAawHrZDu51bw3fgR844VNI5fdxVmKUVbt+pSsRa9kf2qa/14tfEyq7VBsG496dWLomeFDc
LNVbmMJ4cq2N7VJyqrxELVhHjQzoI/z/yVTDWGSL52U9Q7LiXpqe4vPzh714q4c+VDpEMr/Vo2/e
P+drGHBxjBkge/AGxLstmWyIIumszaaUOD2lPusr3j8RJMeS+hdzWzoNOyTvScLyBfU7tNFFpwlN
na1urQfDnJucrGVeYm6Xt3Y49EU6+zxHsrFT9lq0cLvXDf+t2v/ZucWTcwOq8OIBJHNHkfpwQNoV
vx1tAVkfpm7FURm5Gji6n9/1lAmg9xk7rbwbTShVfjR8EVvKNm7v7wMj7WxNjwe43ju5pb8A43j/
SuOybQqKIzuhedZKaEMfcuLke8wsMS3Q4GyoQQFqWshh7J68nax+VpqOghm8gqcnSaJ20W/8uv6I
u/u8rEXX64LynUUDxAmknBBOD4fao9nQpmLUsBQwCAYp3OeD6rUNbWnICb7yuCs/PA+2NAm9pkKk
btwSy43hIspInhySs60asEh6SvuV7/AOgHItPJ/FAv9/l9TaPf09z0FRG+R3Jy4sPalQcJtPdcQ6
9gpDI4uBvHkqc3b5tMx6oC7MA3zkrouw+IJ6QgtqlS4tIb0yU7j8aIGgZPOnTJoBIv4Q/7p5eNjW
8WxhEMuNSa+bERAF/nDF97N4pp1quP3weDWEtjfkv6GVsV483yzxB5IackNT5TXpGdTIJTaPaG9b
2vUIKmI6yAGiD6JNYxmQc2lwEWCIoL2ALeOSR4x7+wF8KgV+YeYbAo2s7LEjQ2vcTi6HwhAktGka
edhERaPbNvAewlzkJrqn0taYt3YieAzJA/xMjaTJ+Me35EZ1zWNBqMX8nL+dQULIAt90lPiEKNgo
waG9zZeXIaEuYR5XTFjAqGnGn79LY4fdR/N/1wRCrnUZJ1XaSFQj254LMuUUidLEH8q1uoslSe8M
i0hm4DUa64L+JddFl/t5FcICU3Vl7K94/PXa0xRBm4Vi4UepABscewR0s94dZSb4deycuj3Jhign
xl9X93vzOyJqxTgVsyWCa88Ux6LOX80TnCkXo4q6Muiiy5xmbx+F5oPivDhyCFZhIIEHsRJ3Q/33
Gh9zsOboRKCsTwUHo6BfgUnBRfyUsmkIWNBbeDy9yyi0nbvQ1HgWrza6Pq92NaFvhGKzqzOyEyJT
e3I2QG9fVJstgxgQsl4Z1LpGLlglzwcHF3W0gOzjmu8FJRaF66YLwQ14dqz1d2JCLYNHDazf/umJ
bpm+M7vMqDfkP6V6F3SHpZRgw52W0qBiZ/qsJ7aux7IdCbL1gkrkE+nFblQ/b1dRYOH5+YsSidyM
R46LotRCSFejGIZKWxDAKXU87S7YIaKAYqV1l4BJ0BPAbiH9vWt/+CMIpzw65qq2Qr6X6NQwOR8q
XGmDa8rI79pns0oVfnRJOQi2FpQovRcqUOIqdaRQ2J3djZ7J+7fS68mEIs7Xt2QIYAnACS4oUhtw
xli6ue7Cnazokee3lteJcN2TQfT1sagZnZUnK79qyLxuGJdCoJxxxnYRWpDt6YrGMSk4u7DtRRBH
7uipsODburxNPqrvg4ZAPSYwdicRwis9ig+PYVw/AGnkPa16/zhJBAttQ+e6yIVSKlsivAcxG9er
ovnJ/zR4S3VXbc//DhJC/iJUwVdnAPAlUPOmANU2/AQT4i18JGJZyyG9kXMKXLvpQmxH8pogH+x+
lNCZjfGvBr7tBOKn046ruhZXx4zGEf0ACJ/eOdNT+k68bK7coaXdaVzuyTw6tJCVovxGTuM9bQ1x
KcBymH/DHJ+zjJa1QpzzmZ8hby085UjqhnMAjpLUe/gcJdaCYMuJU17mM8e3c22JU59LuO178Ajn
9paR6nKjvQG08OrEOWj/25Nr7Bd4MMMGItSm4PZ6Z9L+6DEru3hW+nz3xabr3ADt3prME3d1B4Dm
xUx4jVs1vb12xhU0ZLmMHdQ616XyPJCIzFuspsxveJ4h9shlgT5zQuyAHub5XrZUN6KLqTt0pNwm
45j2aQ6jgUL9pD8qm8qAaoJAMkFXE4KobJsc50haiwbxWGSvCdnGCwDbLLREgEULVmCAZ/QdmJL3
UrfCjvSV7Oq8tEjT1xPnVHiutUDlSK7F1WOepxRwwgsyirYoVDwwOg8oNe7MLIez9vwrrNbU74ML
l9d1TQ7m3u9XVZ+0ZKQW4K8jtHD11T6mG5q/f+dCPUFUaf70Pl/dgXoumuXbKCH6DVWDtq96PdiN
aYl6euC9oCg1j+1Oqvxd/LuQaysZutMbvAsmAcOXIlemyqN4arB9knJqAvJAEPdqA1PZ3KEUDBEF
eLtYT/OgXY0JD+t2ttDTRpLOEzvNQD+zrk3tAxFe4rRn+cDZ6ig4uSXhO9EwsgNKEC1fec+217WB
josMKAAxSXbkqTcv/HkaEP3XtBr53iA46An/Rba5ohHKJH/EXOoSbFjzRv/Al2qvwOyIDWVG1yev
I16WFn1WPQZzb1fy7I7jYOte4zZMVVmuC7GFcyM4tw3mXp2CNkg6Q3tgGfiPL6JveLgaV2mh0hyN
VPGV+yeUOh46B+6SzMBGfHJ8zEmspBMFz3T+ClgOlIZt5GqbgbluTw75u9kvvCB/mu3JrF40+Izj
c190mL2rtOadjwpd+R0nWXUGR3DT4IDVv8aNQXI06OPieNdfFXtoHBfeF4Ds6TOnCj/S9uzPhHS6
5vH/URC+VYAJGbHEEEcFprppW2tLIwYbtbJLgMUgUXcTvZUZfZVZ8KfUEsJCOgVlCmxxLiu+00as
pzxnSJAAp2oTnP3WRa4Va8ugyUnLoEhNBaI5dwvPHFJyqGKtaO5IJZgjHs+7lj+8Cq902MEn6iqv
p+muenxgQGDnT4JGiwpquYtq+eQ6JIJb5gDFXTn3qg4l9PhKw9ghWB25+9zYPj8g710MUX0yjzFM
4odrl05LNSZXTVYM2h1OpJBcWEUS6xyPh6ONqctbt40pGcbz/5WRZYHC7iEAzZ29Dj2K9uFh8bTO
9fVQAcQoBxZ5eDtpyRqwgrArM6vQ/OR8RzmtIQRsI8peRR9Iw5MkkDchU235OdvDnScYG9tnVv51
1gcIIAdM0IP73l9kbpffqxsurxxcxGspMgp08JoXZ9M04Prb4KeudOi1MAYuNZ2l5rF+InrygYh/
FjLjzOEc3Y7Cu/nwbN7xL5X4M0umH2UEeOKNfI+OuHs/NTVUzm95gv5uhr7cProzalmTmz3SOPhk
dMmlTngLds4S42CyMS82k9BDTOsOyZGvEPFwsLTiEuxFA159TfW/zYf7mt08+cIOr0IQGEe9Xw+5
Q6wjwbJ0LVp8Uoom5Xr4ECZgNlQMv709MKbUclSHYkWHEohQd0x6zoWgps33qL5jio3npuUV1hFn
Mn40+5MRYpCJNvZEHbLDMtVTzgHzd92MykGc6t9efrdWwDEEEWA69smFrdiQzJp45zUGEWWBdgQe
mAxt7USrjd3hA2kgkZKfw0W94vwxKdm/p5IWfuk1ZlPSpgW9yN7+8qZGTezKbk+C6pEmrl2hbW98
EZVE722EYyfCK4kb6qXEOrzTkUsC0dPwnr/alAX23rOAJAgvfY8d8U1FdCIIo6f7yEZdha/LYByF
KFA4ub7wD9uF2hW6Dx8xvZrQJl8M0W3QiaN6m0GLa16tgkqV9vRLgUFHIlCSJyavAU+HWWVdEVsi
7uNQYiDXMq2HMq1IkQj4LRAlehZo4HUROOAYU6sfpdlGjgb908mAaOZKAa9xSpXTGPYiVNzQC7/X
Z4OtHGRM3g9O+fI/DR4iWh0Hy/fhNXihOv9StXPhfOHIfxW0Coo0KVdXKvH05OVYdyzWQOEPQpTu
vKCJ+DyCByP7zehNqjksVqWd2yWfd3ACcJLG+llAgczIYrpOWhZQYKPGudFQGxUFwcareZCyUlVc
g34t3HQjwnJYu//B426RrTVop1JixBc60EajqVI1pTLvc1kdU90PkqGPXnWlLJSBSAWafYLJXYiY
ZGPghnMTQjoiMhaqlpbtImo7XuOHqU5xFp7QmH/Baa5EAIENG66b71Ibakbg3+QHVFy9UBxjkSfc
40T32/S0/O4vNXnwgii0+DgmzIEKyZGjq1c2b+BkpWAYa/tSLXyVO83J2ZKfgfj871Ujq0wPiil4
rMo2trIVSoY8D1g+laFCFl/xLyUPiWFKekIA9BH/lSfZGE8gKuagU4mbwBEJB/iVBBQl4ld/zAye
oS6E8Svr8X7RZc4zF79rIdBhnVRjDXKn+z1Hp3L4Uz7eZqB3gf1ley1iSv/apW2FEhpWJe/hQ+Ka
UJPgza2ngv+3M8siIT3qbgr68IatoBhc5HcD29Z8zTksCiF/sYbYmFcramI9c/vzLYqnYzJX/krE
xMowGarNBwey5L4innvxgZYeqdNVIKD+7kqiprtxZ/INYXpxfQ2nYgSM3o5s2umrlr/FqFKKQzD3
vADn+s/xC0nH2A+l+AEyryQK0eA5S+mhouvr8ce+f+vDefKPVS7Vblc4bY5EqbTVcar4RkscDKqg
7T0V4XzBNPSeN4Pd8O4UZT5idWzebeXy7jv3DlAOSl+OsFvvPNv+sWItxQovJ/qIc/uZHztAzcJH
a18PqSs6IivwGJJyXFVJ3lUvOz97phh8/Scwpuxhl8lUm1LsLo+jgaxv4sP0oxZ/YrUD4VxpqkAC
rzArqPIwdarms/KyiBDJBkDCRPq8cS4Gbhsz7q9XhvyhHblny5Qnz/i0xtjLXLRRmIQKqoPeoJGz
Xe4X1yvKUcdICThxjBuXaFDFb+1l5/OLss+GYyTH9uiT+7vOP0LqCCIYFiS1hFeZlOVCREPYI+Gp
+kgd/onTW6fD1WGBZM/qwMCxPJCmP7dB09b1IInzCezgkpQXZAGjcy5YoNqpWkHOium6W53kTyGd
Sa+TrXDsB/xAcdqA7Pb4/qWkiV6Pq8cdR3KKxla6GNGY+4qYN9na/pjKobClwB6nAUmPO0dWNC+d
3c49Lu91QExoOOOhwyHX6xOj1cNcSo3SLFkGGDI1SzVMb/QLvdm8DgFtAlrI2PP92AZCiylepav1
CTylkExxbhWsH50+9YZTV6nomNJ5gQm3/ZW4BcEMEIMRMc1YIAz8F5Bf5NvUAzyTSklBy0Rj+K8o
UAjjyamSp9mP5CaDL/Qtm+4nsbKB1hMSUSu33idVGj2AXCmKdoIGnNbE3TuqmyJd9fVQ9nVgNkV4
PWQtKA4dq/5rEL95TofgPQTp1cVPKCZOcbnRs7CyknP7/P8L6JSLJq6nqw9kQw8QYoezHALNPJWr
5C22x2yPibiag3iUU0cfb7z3lRCBfTDWsv233O9Y9zQKIwvfH/SmISo81uPLuEOWc6rs+snPbPS5
06SKDlDN1I3d4JtrODt71pn72mXa2S9CuF2AOSGYvZGGD3u4rZFKGbGfmRYeAhA2DsBi2gCODS9p
J2/+NXE0bhj6wNSROZXtdmTKD3Ofb5Sb2OQ5wsKC0An+lvopAcebXQwVfppSl/LWpCCXzwfL+V5B
GYSW+iU5X+tyJSAjtGSScsYVZ1m5o4OF9YPpGGWz5kDdtKSbaT1qDAXzX9xDYiD9zeqsDlocW+G4
+DEuA8+lWIPFPgOxpZm3FS4vBlHaDDc6N8GRNjuLB0YkpxSJ6qyrjz2A2ve9FOrs8eUc6nmPSXaU
GzfXqq4Tp+owAtiH05Hr55RtO8VE/LEysJmeGtNwZDwHURz9rPSec5aZjUgoZ/UjpgDsVaFhHZ+N
DjW65tmT53dgmkexl2A6rj/ANgL0zs5h13+lSeRc0utzNnWZNX+Tc99QYuLVV/B1u10inCGbTjo2
TmEHa4HBsbWMo/PN8X/mUZwHpq/jhIaWyCmhLFc8nUM7xEjcexTijzu5pZpR+pxkctM79VwxbZ3u
XhCCsx9szkDuvUxW1J736eLGN9DwhgJrU8eB6o4p22fJ42Rcu1NRN4GH8JQvhB7EancdepPRk4gu
ALmUG2Sm52ajzuCJsz3RAwbBdagg7JlQ95D1Y2MAsWyBRSiB8ICYQYGMAhuo2X07RgtkcFY6rc1F
gEUDZD46eV4ymWCsseriUiYPdNb7q44WHx9Q8TJA46VV06zbI3Kv45NP6gD5vOipX4VyDC1zSEi1
XwRFwvQfl9kNUMGBvKDBJbjUK8B+tx0M93OSedtclfjkK2qgS3aq/yGbWXU2xBC1Tn7KOzN7EUY9
rUfpS+mN9PzT6tCCLkBFmPgLA+/U3zNXdampwmPO7/biMWQNn1SJAeLDSZRC0IzK9LMZPfXnIfeg
1N0Vek+Hh+hkzVzpEo+xW/g5DYD6Ojkfi13o584t7/JdSvinXwd9mDDJ4EvDxCcJP0cWKzAaQFK/
2OR/X5Ct+sBYxwN+IdAAHPsJ8AC+6uIzeOLJGhR4H8ZsNbCOYRR1UKibtrNkklNXRrI6DqyB2co/
m/KE32YhWiLQpvMAeHBx7wDZZ3v65I5Rq4ikLIDar8YaxpYZ3es6DGmccWCgt5dkukrWnrjghCVX
vM3C87BGH5D69mkXSCR8v7IIsZaAIBUN9iMJMsoVXsHeuPVRhkGdb+yob/Yg2P15R3g9qDYEXxXD
fkip64pI2lt+nvX3wd6K8xLpWrJj8ap1qy6OC7l4XTtbwDTtg7iqK9k9cgrIU3Ok495WFMn+qHcg
0dRGG9IMen2kiAyB8xDJO3ZTtzfS2KFQuLB+SFNJtyI6r3vssb9OsZA63M7dNQ169vVZERWDstGa
uxAvyb1uu+QHYaRZmPBL/cKFF2dLAf68yWucmvvjQmhB3wjE+GnH95alvyp/w0aASrGMrPfji2Pu
SXUs144YduQNm358PHUa47l5xUF7gICYgo4+BVop2CxDx45M3SQY8qR8LclpapTRYuEeu+quFHR9
NanvXPRW5LAnFSTWHXGP+/mzfl9/02ah6J+Sd8e6WVedxA/yYTMvs0C+jcMAoIaroJ3YA7rT/TP5
ipJc6U2x+kVdoj9a1i7LJPv6h7KYAD1lJVi5PmS8hd7sGnkvhaO3ZIt5NWdefJVR2EHure3nu84m
aDePqslt1fzyxBkgY40B0V+XPR0ente35cqXJDDmsTzN5RW3kyTjIdVKWILu0jV/XVCfvdmoOnhS
IcI0EfbSgCMygY8SHWTJNC5w0duuord0y8RbbpDh6mHaBR7q+1GmkCfL8s6CgCNy6JkVj4JqvZwt
LDYbMcMteBCBKeOfv1JnxgU+66nIyC68TP2lB975pghC09OSXSkBQcWs7uSQmCpk0hJ67Znf9eJN
WuAThiljUVDWRYsgjXGVzU/+urA9FDrjqhCMg4NC3RI2l/x0sypk/dR3ElFPJLt3Wk81nEmFOfUy
kIgFCVtKT6hDjWKGUcVZ3Rc1c+V6O1AUkJY6YG2EjThCWS+0Bpw+ecTVvq4N8jzLB/EAAaQR9r4r
g9mzzS9ye+bUGwgGZiKlVIPn1bAS+NIPdaDX+iy69bK+01kUBQdeFpyJN3DcEmZ7nn+k/6NN0P1D
AYAbr2DHWpnTQEGG82ROo6WNQ9bGnpYADeLjE1fcq5dbN0klfQ+iEYDr5hui20lDKxx5e0ei4Bqn
YBvYdTP0kgae/YnR55TN9hfpMknZgEbsfCX+6qiT6k+wqoAZEq91GkPsD6mHgIUULrjCvF4FQ2n8
4tRJnCHiogHXGMhLGI2SQ/YF3oNnR/14TBtc3T+sRfzOpNGag8DvErErpMeL4IEskRX5bdZYDeI2
A/HrFnTTAlwjQbqhC+9J+nmFMMIql5JxhZwOsJ93wvTOLqKP5Nvp6pBjJQ5BiwjHkwoK8EXvWuPd
QJM3GqIyPb65ydpf/GgKBl1v6eJFjmenoM8e2aBxbRuTp0YTuNceF0oJX8ha59zLsuVWDYNmGgyP
q5gnOsHgLS10uz6Ot4KHUA/tMfgDXD5pmD60UcShUvlyb6lqgtS0ucr60dH3CFpq/ALwwrQKZGiw
aMqroPhSMysx3fTrNfhMoWjIOmZtC0AhaYFXY7D//c9w0N83nlo5yRgQU5Sgb/ks5cYWBWCxGQmq
wmXIfS82fbC1SiC0m9U1rVT9miXLyh4FJCYOvLhZTXlKKJGSboHPOCOM8f+V9D9SUdBzj6SoGML8
FPO0ZBVQxQsSdxpOTaREO0u7r01iKOkvF8zjvn9mhLYDlSi2/fEaGERHi6PM5mv/SfWYiitug+uy
ijpFYFp45xZS1jFKpHYTfNpQEXPl08/oEwAmvxWnweXS2I/V1mlDRqwvQXON/kyH46w9SNLfHuhw
FbKUn4tG/92lH/LUc2mnjQXvaCH5PiNx0cWySse5tqvE4cZEJ/RiEfebBCHjtRn5Go8ZYXAK5oYR
a8/N443WXtO/m7AJeCHppAAX97luHL+yh7cqjlqNaaPgdJkgupEs9xGzoFTz5rDY0fhJBNrpiY0e
GZgjnqazYO218w+f9/ha+R5rGHdbdulJU+df7Ztx9lKCUEdo8eXsCqdI8bqveqxms2vv1sIBgDv8
NJNz6BFOrIL3WpzqlDZ4oLjsJJ0mCRA7/Y6/RM+o6QVrBfOezlFLI7Eak/bZinozd5Iy0vhyGlhl
x3MJwjrld313GzzOQaKTYnURdZcR98LcnuKeAAFOb2sj4wzqjrSJFpCf9QE7ld7K8uOf+VeFdbAU
0jtB8UFTyVghDHfY8zIzKYEroXplVexaN+h7Y0s8YbYGykE27cZUQ7DUbYQbJ2OriQe+37qynvkL
Pd4nNP6tMR5X0PAjhZQao9jV7eVod4wm9BrTNhX9LKqX9xnTQLw0/aFKzOLGlsbKpMQAiAq+v03G
iCHFIVYHSMLZzLaAqqfMtA+Xl6FDsk+epQpdxf9F5qFWE+lsxhG6Gg88+R5sw3uTV5eSMxRIWnRx
bQJiK7M+tGcMbMUWoUacMU6RFL2PjKEJ6ZxaQRJzoFT6y3tLe3zNKImDJOh6Mwm7vJamDuN4NS7h
/qjhtdN9pNVfmtjwNkoI9a4+2ChFVQWcbgxaBpjxkNvYeo50iE0QwouGIxPFKnIA871K0qnnShgF
FzlkjAHfsidzaBrS+8pQ+zlhgsW29u5tEtnaRI9ADBSihbjnprAVKe9IYXeXCyt3u+7vt2tXsuOH
RJ5vzoqoYCoBpHvyq3bpQ/sRJ/aCNn064m8/42jvN/9CIbLu4MjtkNVOtQbOUFgQB2B8fr0x5k5S
m4xTjkN+HKS2eYO2mj6EURcBKJDPdgAYhV0BMvwZRy3yeFtfCOR0gh02yOXeBkViV8H5j7eqN3C1
qbrO1PkWVO1HYugaTAxQuHm2uS+t8559+A3ai26hnAKP6jBKpCd/bveXPFrakwuLg3M/Hs0reuLz
/S17YpB0TjOrhqrFPRz7yRzcjQk9CmcW+TWuSdZo/dN1XriYmMqzG21USRsCcVmu2RNChvdlG9rc
EP7EybiTVUzb6VPSyeDhzGwm7VXgnZuXxWQmUP765odUuSRiNbbJaviubiEQclMSEFJmpCvfy6gD
fPjOaolNaH4+sJbw/V6p1wXvQfUkwevG4Uk39Jw3zWrlIIltrBx62zFjBg/wK2qBawB9J+7FkXJo
4xLVhjb3trdpUPVO0gHUNDtpLWCo03KaX6v6MB4mJVNHH0GWgfMuP+E/spUEcZGDi5CTjcHWomcR
UCcWbdrkG7D/jIBvGvIL3OLkhLMZV0mWTrHuUiEgsSew2DtDT3Jr/6PZiRd3eICE2A5E6DvCY5th
0Y7TveStgFHXCldSzca9cyRRVkWzO1C5c5yPrYHmajMhn10NQSvQ6Icz1m3KvkziTqMA+vRqXg7S
3HGpv32gRUiR7XCrFT8SGr2sMA9s6aY6LPyZQU7BtdwDPTv/7Ev1J1cIbvFiVtbkZeO7OHkFAsAv
yRbAl/VWhKhW+tUju2O6+pc7XQ9WI8sxeMLHUnSPDILlg0l5K1CmtpiFiFDmsTHjmG6LAfxBMDpk
J4mW+tPFYYYN6LSkPCZaWl7OqwWXsv9M/nckXnkmZMVJQq19sM7LQDtxUUBvTyedkeeOKQwtlo0o
haNubRjT9v0SKt06smUCu8yKTJvwar3YPNpHmbFDx3QTv2SpM30cBjq2v19547w//xlz1nkQ/agC
IEFTy58Cl3Wm1LMMlrzt+i9SVCyJXb+VHFC0Sc+X+onK5l3XdDnk08dBAIJAqPyv31Okkc9iOFTJ
rD2KTbcDABAxon3llAlWedT3B+oi4Z3IO2AS3/WCSV8l0M78G0kkfspQDPdDT0SJqwGRsy95onmC
o8zEHguaJDEgFVq1ve3dgDhBZUqboM07P/QIpM8IQ6XmKyBc42AcAjP9908xOPw60lWCLi0PcD6r
fIAmMbpzxquyv+P2DBrcSHPy9j+GxuzG4mBDSJSDHqVz2gHl11XN8vubNyGlPO2x5mLIBljIeF74
bpTlD9znrBYqBarvWcT5EnqbwOar8nNr0l1230Joo4OCT5H9v73d6RXpfvrXo2fQx9j3RA4E0l4F
aiY0YuR0ITlJXfyvreNq9sln7OndS97HIW+lQ2Ry4mGW0jB3x+xKYv3tTrt7L7NDcOddxWTsbheb
W3wMdqeMZCYgllAe+hvWDQxGaQ+8ennykSkbMG3KquRZkgpBrTmKCso15yi6DGi6DcNNY2BOK6yM
Wp3FuZlv7rojQq9ulg6NoryCriimQvojCdgMRPVI0m6T8ssS+Lzp4xURdljl8QAfncOzG2K2uVuc
Qp+RNmWZNfeiKiu3QdwdOOliQDPLZnOZi7mtl2p9IhU3hoK96rzLzcSpCeA2FRDUaLnkGw4UXmvg
h4sJz/oSGXDdE918eQGzx3TLXh+C9FSFGm92mcxVRSd30cSmRRdMnDvb5Qixea9vZgaW0IKVXWHB
hYbPBKGy6za3G4mV9eCYMxolMs6thYM+kC6QV88LJToH15owsNhTaT8xYwe31smGmI+/It/PxQfO
2gku0e8yMNUAWZR/ewJv2PxMcF44kcVfa3jCU0IotBeFvG2RRUzgkTXMMt0NFG0cVHFaFczEc1+2
fjp1rDyyzbNUUZ5HduH1LFC2xn67zKmM45cIALU3QVGC9Bn7KIMWov8pu0kuf8zDsi9D3cPzjywR
rv97Kmgb8IEfgLp+6sL8rMOKR8cJc8ad6yiYKgHlvPZjEWOCts73gz4KPEY7jo82edIwSbrM+D7a
YTHIt/9BZaxPuO21u+xT1glqRfqglXHhseNb+UKLiw7G4HwL/6cvYs06zXfKNb3gtTY1qhsptq2b
mPxyWBbmy4jCp5xehAJNuoyIFZ+/SXgVgOManfaVrYBTnDVBzuzzxz9Vc1duYnnOrs7iOZaOXe1U
0NdgqWRzirIqBH2aQd84V3IdW7i/OgULBrqaezwWpZrUF4K+IfVwEBEEfiWPtTPCj9Kn3pnF2Fgz
DkJzpyVyMb1s9OPjRqZnCKQ81hWHXwVYGAspuDABVmXorVj4QQ46Tiu8qbeUynUCNVbDKGmM9DIE
p3rMVc51HDlOeW6qp/hZuxMQgXE8wdVAhKt22iHJzcabg2zKxMWqXr06B+dktSo57iqn4wQ5iP1Q
yFo5238sB4b9uEy13MuIyy1bp7+7GvNevt+OSJjgh3TCiV3GpVFqLabGe77gYQW+tSHurs6gmDTS
eJ5iWDhTSSHmlthRhQUAVAD0RFXPUY7d/cTtr1RJvyXLHB6mYjA6pmy4bNzi4BbaE5qusS2TFOHK
U7upCCpVbU701SJIR7bxDEA03rYRSImxyHrckaUOlzQ/XI+/3qV3zWX5FJde7ilutl3BmQKzCJ0v
UC70A29/7hHF6nH4N1+dyMCOSqMrrIajs0kvb1/9IFtG51JMPpE/KEJlGxbrZ1b/UOCJyuvVO1Iy
x49SjZtN08d4CVzPol+2koMDGwueSwJx/q4l+z3quheGzkRK9RgGkXmanpqYF/3JvZkMBEwZ2FVB
iEW3C2Fqv5XHOxs39aeJhV8hHOK4YCC3Rcyw7FcIK8qpWQUjw7Kk29ampwTvBpTTrhKyAqFntqMh
smprLwWoxsTB5KAuLyF9W6t3GW/GYZalf8WbAHeklnEQWdyOkOuS2byt/XaPhjPcD486BLES+IcM
ZdDDvI5dW8erwY06Vs9AFmtUs7PHtnQQMUsGgwXLGuNZy+iX+wlXbh7kLy4dSTGgWcpHwdyZ64Iy
KlfI7XMYwz5sNbw/kjXJxhD+xl7x4C/IPkjrz5EzXiNNzqhXc4OIrVMoon9PPx0Yc5e3RsKFh8fl
5aMLMKPskHcatRfDHfq5qM0jpbnXfkGzBO8azWumzVp+QXxrPVwAbMEs8475X+8eHiYsBqCDmSwF
c9W8HhxRwMGcHSlVa7m5pJ1LuIzCmzVzYTqMbW63duY6HIbfc06Wd/9zhMq3smUqGD8Xair3g2dz
jgLpvGSrd9fiNUcsZXbNlPml1IstWd4ZQi/DUka07Bxa80Y9LdvlL98NliVuIq6OBdspLrgInOmL
Ia+ZgyLjpvW9k0QyjK1iW76ayIo39UeVLkeZFh7CZrpg/qi7qPxzNotsiZs7ZYId2Df2nEMCt1Um
TfwW3lHhhKSyp7qUD+IcguH/3d6BZCAx48oGUGmpM17aTFzaqs1kK8qLraTNVfqcUJ/Zw0CY9WnE
ftOHakclwoGpEZhyCFRWaG//VqckoneRaXgwOc3c63ZDZHQfSOdi5zzhAj/sOWvJc/j1qLzP7eoE
hzMjOqLIP/O1lxVweLgUHXdVAPxpTsPVOUoN+9MOI/V9uLE53PBXmGXs2jnqejiJg73BkeEasGgd
Ll+dXM1WSrVZONY4uA2G9/WEfNd2VrR9ejhoixLVUpmuu3rKewA+J+3nuqe2oN6xCm0sFHraGHkD
7fHClFd4M51//zBc4ket304JLnZa/wR6ENr7hOr1CitvcwoCUMqe1gGMiyNx8oQjNFn3RqgGqUV5
ejVNQbU1KCxvfGmJ80b3pt736M9MDADFE3sXHID+T4jVjt2aZtJjSNlKt/OchI94CjfTIPf9Hqe4
uCKTjS2k4326Xj3LYtXTBOxRwVozeS9GoyVyFHwsO24si73VqSfX1MlArpDlGhKwJ+l5BR5nWVwR
Lgr2P6OBcyaH+Qte18YktaWibWJVOTmCR9ujhdLwmwdcBAhPB/ToNIo5Z8hXfyicMb02B7VvC2Ne
cvEyTbj4Zx1gJ4jtwXcB+9WVkC30diTP7TMFwlyuyCe6bWcjaQMmCU8kiKcCPYJ2DVCTcmD+30QY
AsfufjRxyw6aG8qje0OX+mWAVJWdAuby0Xh1fDI9gPRqGJdDDMJSnywIPzuy0jVNsR2YPXAOyNhD
GTpwcgdwjaXfQ7I2Ii6JHxsuyuwl3Ey9MKoqL2Wy6aEDMO2IgLw3ql3+u5XetaMnOQYMHUtYAGjm
ogRF4fxodhZvECcnUnusaTw+FPzvHLrMtwDgxRGXEON7qBTIWDlLjJaj5KUGB+Za+4h3DQLsSMiy
UBR57TntW7U932mAEO43qOqVlBJ7vufLdGcKMyEsxZWucjOjjGrQa+xZt9JUovQ+uDT++uieodGZ
cvag5EXnhjLQdWaCR0NSuZeyztng5PqYCxFPDk8MO4PJDlVbxj1O7m9togvBNtogYvYdqPk0TEmS
CxtgBP/TWOoy224aTtgoULz9VHRACZ2FDc26qfl8EfQF+xo+RceINrMINGL4eJhD2FbLAVEXJW09
kfV8T8S3kmLo05/AqxovmY/OiMTGl65z4buYC+q1+KY1hAXWcjoXLaMDfJCtN1CMKWihDps9gzQc
wO00gvYIDJHNme3+rlDrK35BWH/jDQcvqfifqZUzzUprVT9Zs+LVhFyILmgLfRDVB0niYcmwzl1i
M++sdEeGLMQBex2Z/WV/2+8qTFy1kUxMSLqzrmY3eVNBDAiDqYbpFmczdTNetUbQBCZ5WeoiF+SA
lvHBklxRnikBaD8oN7pMPbI22KvtM4Uru0jURj1x50fjtUvqaOL7M+kJ0eo/f0woeYCIfIzOGG6D
sRMkDU6tm3MA0Vt92SARHd/d0XIZGLFzJ88tK1is+2qvfej+y1BxZ86aA0K4PDFn71JCh0Dn73y4
N2eWDY7BWtSU5Of0x6isJcSkSuVjbNG9INtxVKrLxQQS4Hx0wuS2caBORaS7MEm2W7hD8kpiKC6B
xIn1KDWOqiIw6Nnz/AD9OFdiJfSO6aaWBOeYT8veJnpSFIda5YXPPnDcvIncK03V1piL3UB05Dh3
LvQBfJTGZbLMq64eFEZ6kU4V0KzTAgneBsoUKafvDxzK0nTOLj6FQKeb6taw0sZyFA2XkVhaoYZx
zy8uPe24TxMIZ4DozFARsgnqiZ/T2zAQllxmmEGn4Q5wzKFS9taUuZu/eEvApZsIuKCOLIoQ/9l5
jMpWfsIlqlhvim/090xfa725PZImWO7uwcOd2lVOpOrPV67F6JDfGXOyq2ysZvUw0CTW35dNuO1J
iqyXFi6x2A1Q1sxSu4GQC1RTWJqSUz8uRBtVH5/x/vyVUEsvk7HQd2M2yF8FEvP9YD5NpuXgRbPz
yO3/+dinD7P2b4ANrHJqrWp8nZvV1lpMGyzF6t6wvLiV6V4zL9+1LEEN+tEsHoya4M3E6k2NnbeK
nBrW9Qwd2wPeCmJORPJfZV3nmoQ+KADmu5zDhXAwBlXexW/700ItfZhDR5fS8j4ZXbYwDvnjt/hD
txdWOu5CD5ItFiW7bvDuybFUcMYTw6KHW3kNO5LLC3qwMj4VF9Jgg+Hh3b6+Yg/emoeLKd8VJ+ag
FGIPnsFQFRPz0mcO7opyQY7czPmf3zXQs1mYTaOsv5Mo3M+oP2ugbgbaSp5s3j/YVDWofmU6SFDa
ko43Ey0bo2Hb/zXBTv1qfgdq5/TufGEFacFL05YRk8ShkV9SCTc2cmqqneOR6Wy7K/Tpl6H72PBO
Llv/LrK3IBT4zBSjbZNtnsAsnJ/9qZZynBJl9m/VSewPtE28DmupR8wDQ9ZCtOA2IeIHlDQotpcW
c0j4x5iLw/kZocdk7VID1l5/GwMM4OFCdlixP7NqWyW+tmY7YB+akKcFpETWnXafOdd7+E6f9UNp
GapRW4FdlT79FLs1+VcpHGH8g5FBGTbPce2o6ecdq0MTthAkysCkpLOR+1OqB4CNBX3JJWNR7VTx
TwCGJGA/pRuy/gQWxTq/Rh3SNspGFBVbz0kMxSy/GOT6FNaVfmrd0AMMLd8OFMmHcGwRZ6CmwRFY
M4Ucl41djTAUf2pAWq3UaMihWw7vugNA5qLJgQ5gYq9mVuFlpKKdG92C9VNF/SI0eMsq4djusiAE
nQnzwYe6lfwafU32kr+ppF+tEKkztW2KXdUnhD0cNrAjkhlqxemTwpChR6TsaESi8qxJpOwcXkfZ
rofVCtuLp05atEmCPREZ1jQlqrtLJXxPAAORrLRHMpH+XQh2Txyc/2SsZx1PytcvN48LWGmUX+w0
wJ8cpj9HhaH7pSi4npP0m+4/DRobbhrLM5idcnG49cVIMndmN6YfJR9Y/N3iVHxTcxM6Qf0Eb8LI
YjAKamKkm3ovbpzNDzE5/6FKkzEfTWMa7bOUDtcD0+XOZsoi5rA5lhOdYxR6Hhn0DqJCczuKfUub
iAp2dXCNVx6WG2iiVCcjTjx3jYLqgUEELVUcLOMNEiDyd99KQm+WqIRvp9Dt2s58kYXLT6q3RuQ+
dVhZv01IdY+TldUoRH8C0psSwCWiZr35KPYQRKdrxiCvuHECiQ0qvz8grm+L9iX+Sjw8KA4CnpIY
NNdD8UlLe/FnKt0jlTZGD/vq7RWVXAfJiT8IjYOsdfqg4bBcgpd7eohbRi8nxx9lfxpgjp1qDpFm
N2pG8yucYt0eeaIZRI4ndOb+USIBogt76CxGq21jziVCYgZdM5t5ZQbH/rbK2i13lW0x4Nr9ETlU
onYluIoqAcZ+CgQaPWS/3mHQt2IjUdnaPoCd+gG5ofuoYMeOlJXlZuBZ1QKSUkuDScRgAhoVnWXK
VMt8oPLGiEOhgx+m6zUkJkdFIqZ27iOjebxsQuLfOEny8f/OyAr+i/oxg/oh+kI6rXxE/079ArIN
KUN01cQpBIDwsGFm551WFHiIH9h18EXk2ERXmJoXSVIxrQ9yOQk2Ov0Txlc69NomNHGF+p/1lp3i
QDrex9KZfcR7Jk2urUS6lopzYy/Uz6blXzVWLJiXzWc0VJkYmuyvQBExnqrWARsXQSaFMcyiU8wC
ox6M7D2noByw+EtBBS0+oIlH6FVDDMnR5sJuYzDMeaIM+aak+oug0yq22YME6LCMEJtr5M59ECkI
R2QgBvZPOB+OUCFSq4YZFNt+LL/dk+I1bzgOhtntBZDP7ooYqkPjCHKPEQfmTt+e/f+SpzIUf795
ZDp6gHlQ8kJHPmgdsiGakcnUpgp3jI0n2iweylS2V9ZTIc811G/Gb/3WgNlSL31+YREpqFJzQtOr
9cPzrMWpfv/EeM+dcP6HrjkGb8hKUeWq8CkXxpDjPJEG6mWIgiAsMEyMZlI5EOC25LJ9KRBN803+
96shVmI8Gf/QhpCBI7asr77kMJP/Z8qNxctHhAmeCkKRfhu9/XY9JhhNdA63rZ14TNqN9fBgJy0v
7LThn8YgXn0SS387mJh+1AJ8YlKeWfa1t8EAhg269jqyBHQn6G+T5mo8u/EI5o8WkyG6FIQlek1m
RuUDEe9zjKKltVvqcbAbvWIrMpjsoJ4kDs3jEvFhQAU8uq9KJMKoohK+Ut6v1PgsntLSEG4m+Tcj
/tbN5sEsSskwsCGIi4BkOjlnQn4EuyUqmohVS3NW6mDVFVirHPXeBCqkROmFfg/PwSRCKVTsYYVo
FzHSrOmf3Nzr3vnyzw/Ytb0P07J0TpDMxIr5V9vN2alidw0+chJtrKU29HtJvPtnwgh60YYDn7Hz
CIJ3+uyiMxr2DhBcFgnEe7xlsfuBATJy+xPHepZtZFpOlhiGfGbO9I+uDMZaASExTrCp1Owsa2GE
2lnR0gmXvyQoBE+z4zAitLh8dA8+gouHVTz2aZ/yQh/cEUAxCv6GbKTJwvKCOoFl7MeMlLrvx+Hi
ghJQPuB+wajwB9yHRZ9v5nWXBZFGBhQWThazzQ9SS558vQXn/t83teLKijmkhmJzRRkFDVTGr4BO
gbyixGAR2shMUJoPl2VUHV2m/G42iw2TQ63ZaCNl8ZbsuAheJhSvX0XCAtGgNnjWXv2pd91R3acE
NX2waoRImXv8xq3SLvlb9/+3R0c9XcVgWph8sF1gf2YCRzf+VVldroVJPlc1a39UFk4OqC/IL/qH
/Y0hOJcym138K9mBcYWbBeyW6o3/5JldYTYP5ZPU/vmam8oCzwOcYtbI+KxMsNnnICox6uP42RxO
e34mJ0/idjIR3tNnm8SR+Ju+7dn29VHo4BOAF1cL3OrDK+bT0Veiud3bNigshk0jy9UH19kDH665
938poZJl+31VsBID7bUKb35afBPdTonTxODTB7KHUt53jt8F7QUd//+nzDQFCxHsfqYX3hUQ/ypg
i8nhvi8P39OSEdboNS/qlACVBnydRIhyIM7Gr+H/wfzn7x8+FURldq9VgFLvSc9gnmxhX7loL3Kb
K5/G735W5tbxqRriU5mWQjolhQUxiUZ/OHNYoiKASmnyqsVAFms4fWMUqP5BU8VjbmoA56W7do/A
oB4fQxamleM8Sv8xXWuyXHz+IWmJqCtpPWQNcCdTHRdZegsB91RHLgH025Fabgei4aKrw5IajRMn
kVhNlQCVroSeMuxpuoP9obryQIaF3eDuLIrqfMvdsqSEZTWJfPT5aoH6Etxna+vIs+Nu5jUVAr1M
q1rK49D3OFTTGWjgXEpH+kgUrjVBkih6WlVWeefWg8sZ2Q2tzPiBQhR1idQsPnh5cidy+4iVp5s6
ldrndemvs5UXYCPckiPA3yn3KzCHubAtNwvA+5C26MRALYY2b+98vQrS5qXHimfN21zw8HhG1sOV
jMj5SRKAdY8H4YjxyusSa9qsa5ojb+PeWzcDYxrM4/Rr5ApMuB8AVLOWSf3t28bpxBTu7sehNJgM
h3F7F9rpAvQqF3dJomxjnJb0INbhYxsYOt7UJ5ddzK9XuIS02A7J1fSGA2pr7/cMZkb0xXwkeBe7
6S1N2fTcuMzsdwzZ0nyWM1oYOOwR05scTUMF6aU/poFRQba+4m435J1lgPFGe5P/w53aPjP4Fm+r
M+EuLWFhBt1jJGSuoEaodetWYXdSESS8yQJbfugotMEaPQFaMB6cR9uf2cDKebTBddlZtBBYVuUz
XeNRo7fWgeBvKRjLcZieJwCsef9iAVSE4M/LodnUwfcoe3uumDaEeG63zZ6yTX9j5eEW0gyvrjlT
ppGVST+GIVi+U9DK8n87sFtEK6muuZNcXxtCntFUl+oUNxSJDxbvU3eNjO+h1RHyR9pw9BpBZGAS
RiRN2xuA/ilSMFuKP/SjarpmhgUOtGcp38ms3NgVSpDRSSOlNvMejj8IBsmS574sfFuf0PH7OSJ6
4R+oP+DjdohB7RUMZS5LoKJiVrzSEGSW4bWJKHs+aOQsyaUNJoLxNInzmOqt5TaGjEmx3jxIH/cE
l8ipxj30VWckS9AZK78nz8gIB2OS/ughoqqkOkGe463BzMF4wXkAUz6u3ug1b4bQhVUe0mRnz4ei
g+zAgxVmhM0zQVkDXyE1aB2hAtVu5qDgmmFGIQxtAxog5neWgVFHN5HTLtHOv0BIzxQE0ra2WLhb
bQTy3YDxqC8uLoqBEb1GH9xLH4xWySyF8xx+i99LV2i4VyDwNB9KDy6dO5xlnSBk8OblNQECmEK9
PZWqdJGVEaZDLF3AbDlltSPOb3A4I8XnEPx2I+HBEDtO/2QOeHP45FnByqIVGyP2m2lWcmtD8jsT
H/4GIuMdMnNOB7dO0/oFQWh+/Ur+ms8xB0TI5x0k0YQKTE8dweanhrpjpMhgOlVqifYPUc5ej6Jt
xjklB2vomA/tgR0VbwlygIzEgomaVhySBKp2/7wLfOhKINFMqJnd1UUOVbTJp/AFhMtTU4EACZ1Z
ihBDoWFFFRFF3cKrMHEO5rGpDTsajlj4y8lvKsSJKqt5DJvhRbnGSR5MKzljXsUtRQ2S7IdTgGDc
tcxyJt5Ih7itY1rkO4SxC84xOOuyN/XKPrBxuqN2g9Npdekv6vzNn4+1AScoKaAeG2fGd6R+UzG3
CNwuSDZjPFxYYDcnSWujhHtVVuRwQ9OhlNywcWLGXZOGRhB0Ymj7Zmd3G2Jxk0gRyp9fNiUBomGd
k5hf73BBeoOKP1pI7JN5n0HFR+9mAvwCZQAd0XSWP96wgl0vTNlmCnsrTkZfdclLprf0D4PE9mh9
urnizoq5QBkdm1iusfvMgzKZsI94cUjKk75OpGoz0A/c/VkaFnSZ7RKSKZ5zgS67oVPh9IoIgSyv
JW6BEns0GsycovjIEev/LMuJtee1Rz1CpjTrI72AvZhY3BBdGJYnxqaRAc7Vt1aJeCmNAUtZHe5U
vVxlx27qTFORjAJIJurBuuiOLFvZ2doigAtaHPyjNIpjxvbi/HmH/CJca1pE55NI2k6ZozlYv5bV
za4sSYcp/fXSuF1DcVej5Dd45X6Y4+hTUYB9YUhCVtE58tnckmsvh5EufZay3osYlf5aNEAjFKDh
u8BZeg6jtMh0Onmq4qzVb1g+/Z5Gqt5H05QiYyse89tXF2oj9jmuZ1ut+pbdaInd+12Y1rT97S+3
hgWOZxXwAP4zV/BtkRqVEbfBbF0vPKXeqAlrqv7U9lFNbnfFUph9211DGWfwXrurGvFnGKh6e1Tx
sYX+A0ABuvkbYKCavJkIRNhSMgzLhzwY6bIe41/QIDISscpbIWmPxHSaQaNDBItbGdqqYOCRlLuo
MvEeoQ1I9jk2Z7YHhlnqqylMYKvdwoxudQJDfATN94ybp0x0GkDDso+NfcbBURJHsxP7PYPIcvns
FVMlr0cOy8T9a7AOCfpe+GH1WtUElV4WXtg3fIwZdg1DS3yKeOpUAz/rzTMUvkTILaC0Dof1pwey
WzpPcZa+/60Ndx3Mee+5rK02ouSl5DoJ709y74Px7CpsvMqDrfDZWLa5BMe6F4flipwvkIeNMePs
dYlt648yOG2RWyiMhY48PnZqkkPRETSvGU8HiCTkC4aImSAlLhu6NF/ze5rD5hsPbkPMgA+04k3m
XIuE12ZK4SryWkk+Fjr6CFHtI1dLg/Tw6/2vIDBUUhSESfGaOEXr/wOY14ZKYcN3UEIo485eohVE
EkGH8hlO57vhqs49QmTWIgisnve4GcQkbTWtk7qTDwI/OycCBum9FdSNM315sRKfyOrILciKPi2w
TIqx+F+8x89mo8PYLqSclS/1u+ZeFWoT0go5wP5FRNJTzfRz95HCM3kKehDYrdVc/rY7xarqLpxD
HRKsbw4Q4oWf5/WrXP6DU54pWvCOVq6lxqYbahvcQyM94S3ZIcJ3R4A/VewDz/1OPlMMU/qsnt+j
2gMHSI6bxc1EJ1V5h22SFx8bA1lOW8gvCUSD5NRb9tz99GeUsQRe7Pn5xXV6YCyCz8xD8gI4QvKX
KzLCUTpFiHKTxbsuOJKyapaDY5bmgK/o+YNkLeiJPqU89H1Y3KDXE8Qss8dIh7fp4dTFtZ4bEi5f
rGO3A2t9RbgnLPjCYequbsuBR5TM9Q4Br/MPu3kDPs3O9Zf2HXRNSWqACboxkJBvfGxUVpuHGoag
AkIH818iSpg0FXiAWxLHRsRDR0Jc+Y8lJ+NFySkYyJXJI4CzEhf0So+Psnx2M6Mf7S9qmD/5KMRD
ENs+4jm3SGH5r2fiiPDgOeCDzR5/YhXk57sd04S0YYOk8qO7NzQlOxRGRb0oS7xhlAhv1L7tJL76
gXUV6ATW5pr/FSpSWcnNfEOarkKnK6hNh7qRtrdHo2YrM1RoMFjDaev6kwCb4f6+QnPuFfcmO914
oVVaZYpqvso0Jt4A5w6zOCWiP3p3IdRf2ALuZGniNX9oBYMyMVmmEJUZnH8NvqqCAIoXe51FWokq
AwEehdWB7V8TFE6AeksLUcC6xaa1KrDzItIPtrbIbvhSNLGOZvQHrCH65byzzE1S8IS5zi3lD8yH
vkoKzsbNG7LtDjZe26lsZ7yhYZcixRsb4z5wR9HunKRUEPpJ+8Yoy/Pu1+HM5XTaCswE7Q+OJi7G
zktyjGAeliZPXJkKazb0wsxttxmoDHFuktC0i/sFcFQowaErLHiRxE/I2Ds8Qh0fC1c/efcAtMKp
ATKc9YbOkexAKxGmSWUz6jxavVJfnB4bEojLZwH3P/2i2/9Ln12SHskDcsIo3WjhOPOn/EX2Q1Zx
rCkuN1865sXW9E6JL/ZsCSm9hTdAAXSCvLjeGD2XHh9EJ12vfovUj5gaM5ijvU8/bQ53FA0rYvTt
zIxhD05R9RLWW+MJQ5xOlGnIsY1HrHtbUW/XD0kFN+4piw0kyt+B7VMbJ5Dou7hrTMVWuyKacgUH
mttUTWAvWNXw7kKBZ8U5m9Hsg7bpWz/G93Inj7Jzaweamgf3jD/7FjIfgGiY3pr5P2idvIHBYVHR
mHYciy5VSoPeB+HjxoLXrLoN5sxpnIguFkZYX+FRal9hLGaBR7TIo4WlI9ffnN7Fkc9zXsYI/3dL
cc9YxNpHq81mtbFjFRbn9VL2LGsU3UlsxDfX+ZFNGQP1rnhrvIgZGucsxkvUNxh02McDTEzalD2H
ccu15RVk/yb9XuF5V3QrkFOhgb+HKc0aKikCL0evgP1T2TXo6HSCwR3YKWxsEtwzw5ci23D68rNU
6TheRGr7jTked7YtmxL3j+ld9eebD76puj1vTD66k7e1SL3TnQet76lGrE/2KJaw2TZZSW4P9P6L
/Ri+D+OF/s03VEUehZHNtX5cJgCNtUXfA1Ieb3UX9BZGJiChXBPeJWhPSjvsmYIzmfrJOMLy5r9C
7WR5CW9UP1DfKGGASe/2wnGwbUyABMVq9OkWA2nQP7V8hqKzPi211LXJy5GV7wWblaJxI/o1CF0a
KU0hyHVQ/1lW55B2+4JVeYv2KwJvlRJP5oW4jN7g2MXzTp7/olATBWjytJJISSJupvlRwjzuiGAN
qse7FHOHXA86GH3iz9tCYw1gYfkm4emFghKfD//7jVppmqzmVVGpzZGObEEdqvbX7XjjfdohMbUY
fht6ZogkXe5UcyUik4Wv+ySXyI1UDNzlP+AKqLzYoZw3VS8LBfHbg638iObxxybNIrO983lvu7cg
NdJkVcC+OrLRfRNpO1Sacm0TkxbUCPtfA3jtZn2uoMRkAFqniTT2bw2y6/uNpfS6+VQUt7IcKDOp
5ZwzfTioslEYjEgwf+3V6/jI4AzRzTxLtTK8ZYuMSaymfoAy4ClgVcS21QME5THFnWnBYjUFE87J
J4GDxXtGSWn1Uv8xkciSEDL3qsIzcpa84EXESSPqbvi9dUz7EKaaenlW31Q+utHvkHLsbu1iQQlA
+xOX0pHDgVlm1e4GEZ86Qp4cP7sK0heX3MamQqNuX8rD09lBXl53o2vvkk7t9pcmyfE404FFG7KZ
N4/77FPPyKbe+Wc+LE2X7AOdaULm8dBNXovpW3LnR7S6hUf30jfw6CHmvinrraDobgmzANYTug7p
E2wbeN1Ntqjo54glk3KQf9+s82Ijtgrdgazdu59WU2NTaMxtkf9psSackNztO5jxpsmBgk53W+p4
0Ea2W5aG+cQgpiz+zp7euAEEmLtpGMAloxdXn4s1Xa034d7x+2rnhRZyieTpAreRUwZGgEhzpNxv
h1pojS+b3spbJ5FRqkJtymzkKtKceD7EOdExp6Zv2wPd3ylSvq06ZiUP3gDrSu4g6HHPRavhx+A5
Hb0Ic+8mjLnLxqv8ly8FFHlLtQQJj0W32SucYIxeqi8bqBpFtBs778oHMl38XZT95dNmR7bZL68O
J+xUk4Zmysz7/vOuDiR44ZCqSIueEJhPY5QC8aEJo2ixRMHTCnHRDYZ4E27xJJfc9fLPZIneMtv5
cZaDctYFiNWe2J3EJJj7tmlbKdc6naoNaJxEbxigAh0tLEr7CtMF02CRk3T3Dj5O1YNlTnmEEDv1
ZBoBVehdNNqVkqlxSFc13MU4DMHRdv4hMIAwc5aGvj+VI6CSURsoZwGj+BEjuK7CONwfzki0mg9a
XVBUv0BAOSUghGdvAlyWyAF8DoKVN+dyLzB7eBg4Y7J92JrtkpptGbwbmz7RVaUkUAg9vRZPGlh2
6qiJQeHZ/X6U5Tkmye92Q398oh6sLJ4a3P2Ri4xvyPXAC2fJUO+Pb/gwxYvt9UllBCzj4/nvOpuK
g8NeNhi2ggTpYYlGI/8IXLX8BpwtPUberQj97unF3qP/r+7Q1O/WFxd4jSm3mrmBiLz61fECChyI
aecnVRzr5Q7NG3+14KYPZJne+2ZpOm2ydobvfzEb55vgGJsFo5jsT8KqoC/4T0yBRF0/vsaH0OEm
ZozTDbr7OGWHbWls8q0G0owZzqZXpiId4pr7XewfOth6X2+s+JkWHDuC+Z+tgTTIcezKU+l4EHGH
nbls3e5SuQireg34McUbZ4F2bOl3OHfiLAlc8N2UZ86wijWqgAht76/ao0HaApmdM/khBkVUTtEg
/MP2v634fYLrRqxgrLdik15VMASgPfNLsISuljhdOe4kR2EoPjp+lQcwHvqZtzSKg2Ha+SqAqNxK
ul4GKtrcaYSmv+Q33kTEtDlM//xglGeYFDF+/eLc1+gwHI4Drwn9ZmtpZSSaNTzjwz+1V3uztjUg
BXyDYTsJzrGJKcqj325yKjjin/qWKkkbQ3rXO6k911VGaMI+vQxNubFPgYOby8f44ntNKOKD+VQX
pxAzHpywi+MLwRN0EVljZqBNiNKV8e+U/1IYEnwbjbqIFKX7wQbmBnZuoehxtk3uFgQKpqq8s2cp
G/oabrePSjkA4kg0s3fsG/MfrBpa5auZs9sfmhDmj75/JzYfN9mhEGby7jiDdngoandM3qoHJkwA
ieKOErjgpkjwjbwLYpE7MbM2IlnOG7F1AozGo3q6i2M/lndnb631p86TLBPIScOajLG/89uNIa7z
0KmJosqtzL/IW1hGyZVpH3i0R5s7hbFSMQavgl4tDAha9eUivkMTCaVOYo1cgroRhHRUttBYJkX7
PUKfzB9s7f27urRnZFJ8wBtGdCgQr85A+wYvnrojiVbae3ICs5jV63FyVSVxEl6P2p87Qg6cFGXW
RHJSNXmxYVt2ZK6RiBr1ccAY+9CgoiWGdQUTa5OruhsCcsEV/bf0qBnw0NbdjAOIsEMAXheYiaEA
wZcZknZl9AVQh5rQwJrkn87mO64z4gA4jA4o6XoEb7c0VkHUXC7wdLzBwQK7sUPEL+Ss5SKTyog5
I4uyYAO6uguhMPhNJsYZxpnB+37y0ohS+j7WzDYdIeXlqLWsKrBBY88BiVqMqe+3WJujzwVC7Qcw
xKMzydE8wmgWcbBaKvoAaJdYGPVIZOEciu8nfaUm1fwwisjXMa6GbXbXJSEp8qgo7FbeOper2IS2
S/sISuue5LAqSpC1MNEH6K/QFcnVuLNi6+ueoGJDitQxZ27BM8kw+vpD65NkjLsWLnhmkp2MRvWH
StqT+A+AIlqV1GdpfuPlksoyhzHfjWXAd1mYB73rpcm+u55NhtDuMVXjoFGa0ne75PAyYkvW4uUV
Gxg1vIxQTim7VcoAncO4LFI46fMyKHVIEiUKXUIeZWhR0jNw3XQ4MbMbsGIZq/vgnyH2jpuvWVQG
W8mHLZZjdg80GwWqkzYZI3pMlyqRHH2w/tefXmiC1R48rkueMwkr/s/44nIkuWNYzq2T4KwyuGwO
iuGR3gPoKWi6xlHqGgUdn1sQ+HEJjj9Vog/Jn1ayUfz4q1p8u53lDyhAqIUpoMw/6QG+n2F5FMqy
763P3p8JUfoLgh5iylzPYP5kWb02B+JRNRkgGEd/tSNmk8SiTChvpJdD+WzH7mtn5SMS+VEro1Ik
ChoR9VI8dZR3IdsOZqPHTbuBJ2pQlo/4PlQp1EfXAEFH2kPgjDFV2KnTnfHIb+TvBfQpyvmI3Nce
F5hLZB6Fmfork1dVRqmm/rlLjid+lR/TPA6+XGzA/5THM5uVKDaO7lz3jM742vWycn+rTNhIAJx/
MsMchVurKRh+12TWopO99j0B7RwA8vOcSMq3knOAklROaiJq2PQNP31CMYCwwd86+ODy73FGPgVI
lKXjXYxEf8rFPRPpAGKmR/SXJ+iO4GmtcE2nJKds3bwpK1Uh0VbtxeX/pMKs/Ur9OGl5lNGs5/cs
Vbbyf3q2nfaC4gi8+Jx+mzC+xVmt7B8MEn5Dlfol3i/m7E4NnUwW4gyV5Eq5QXYnQ7eAF+zOj+DG
xvlQN40QL6ZEBRnBI7Eip8tU5pMIsYFeGTaugssKwhxIwDDJfCab5lGAcwzU9AuOrujnozyo7cbS
SpTcH+Z9HzI2jtMSYivONJU3ZLvzemIP/Nyo49FtnwiVUrkmqwjNVgqdTxX1fBnGTS6/rKmgJJ+A
0CKmcpHrCQwWsx0cNgfBNFSyw8KNlwvX56WkQ4t8HRzQJfW4hU4WTuYYfmx6X4B4a3KFnX3ne4Cz
xZe6jROEj5M2KCauf/5N0adl7qWeuD57cNbrTk+89t0lwDu78WL1510SbCLpYRSvQiCK6sTovACi
rizh55UlGdtAz+fDf30gdYkkiR+ftuRm/1QgFZCXka4Jo56SVW52sBZWJopV4AmIJ2sgZnKExix2
Ade3pHEp6VMvTvW6egjTB6V2e1F59qAcOaJAf9U/GLHrzaR0vepzR8mgy/FtcPDxlIWhsIDSXcD/
vqkjzQvWVkpzZutiQ+YJ9m2P5HEcl5IfjA4vYBJYUHRF95X9gvtDffY/ZS875xwpuGqxfBz8IEjI
Awv9LqlPxotVszUo/52cv8xDhiowtfAohhoYo45LigZ2wYmHgftZD6HuBrmRNPgjm4Mx2lf5A1Vx
fadcf9tX9xMgNHJiXm4vJQBoHLk+OBwKbQwAaT4VXJVurJk09dJRGn+0bR8JV+YZbyqc77ppa2oz
ziwZO63L9LXXwJSh7eV6xRqNVjPCxeI9qa1ZHhd+PVNX2zzzgyh+tcACA1bcnF+q0UNpOGoJSbR8
L2fGfB0CtEYnXv4m74lgd/PjqbQ/sEWhEEVLBXtQWmNnkzr4kUViptymk3eFSsTpe0Tl+kzoxDTm
YXLgxtUTONXP9WokM1B2RjaOuCVx9PWmkS2hsFgEyG9391Gyo6M0D/EpxGccNhk8SIVlw6qSN1Cn
2DGTIwUxeFb5UNhwo9qPY/of8BCt/MSA1bcDFuh6I3c7LNI56OIgUMQYGliHKqFolq/KJHrs4TdY
ooqAr9cdPtE56pXzWVDfhs7VFGurMQPwZU6qPn59g6ZtNjOCI8MyQUGkNMbULxd215NlK19F8u1t
g6nLxSU/f9oZ8nfnjsMzXUafF2otTUPD+p1PCe36hN4MpHFSLuToWawvTQyY4+HVKSTllVkVfaf4
aPHeB1S23QZCYm2KhI1wEPaUj/kJ6qnJHKqvNZUptjaAkyfo6gDUeN2Bd1tr9OCNwdzwLQEiGyDu
XVMm73MAs3JTDtBgSoAO9f16LMau2LFvsvAFxnlFNnIbeic6qg/raeVjSmkeb1DbiuaKuiM7QXzc
OX268fVZgPeHlM1+V2V3YQZhRv9YhdVqbwp2cF81i1iXqqrg5zWip0QcgG6ly4mQjs5xCVx9jv6l
u5du3ov80Lr4WdNHKKGCTzvPanUHlLWyr6hRk50f02iA+V120tBDhj93QRb0cio2A6OCxRfQ9M3V
G6bVH+3pW0Vd9UI4DcaV7jwVYf3PB8ds1L/WD/1pmBHtVmL5mI5QcmhlaQ+jA0J9ulVhlIepZChJ
BZeeSe6mvs4tPG1VY8zFianqzWjuMwS1fbmgs18VVi9tlAj5khvIu01N8T/MN2sAlUFlHIc3nPhs
xRYqvWDeWsUkgprfI+HpQF79/tEAIIsVQdsW/7f7u0kmMogx6lsNXM1Zughy2zdoEGJpZLnTwMqo
3ALsTGZl5eq8q6S3fqpGvHo5zpuvU/Iswo517MoLXr1Jb/ncHtPRJ764M0xjkwZMVAPS/+V1X9gK
N5iWLwxcoqzjqrXXFrtzx3uROiaKpsRzP9e+VUz/O9VETvHxPECCqeLFgQI/K0jPKqCbNdpis4rm
NRxWeA1tY7J7x185JaR1r5uSqGxxi5Mng27SXkx88s8VsPPr/c0VDLDJXXC7OM292SnpoGFdiaOO
A4KeS+TbG3WMqpRYIGdjdHOhaWM6QVp04jxlUWIx6j5oyTRMiLlfC1HGk2NQS7hWwVWO+Keub8Me
wsmsutC8yUMzlXvUilghJFmoJBbaAvJYKxY5+4qXp+jrpRmnHKsvqTJiyEv0g3GwYzqg/hi9xqqp
wYAU7wSIpcpFQpw44/FKwNnvzozOmZQ/N3nM0w4c87PySDHTGbGkDaMg7+Bob3c1k4q+RWKfKtz3
4LsiorVelfOlgKQYiZDvkBYBg5gXCOnBlcPTd5Zrut975qwGJk6y+WzCklrtCaCojdDAWjo+sAsd
I4nUJRA/7Wg1bpb+savrz/VEBOKjXAftyjCUc/s9hPbxnZkl4j/7xi0ydeMJ+ymviH3tgLCEcb3F
Au+qkkL+OrviX41xSxgJzsufy1lzzXgpX0PZ55+RA7kB55OufP4UnMgO7LCoYhlivvV/KQ+Nblmp
sk5ny2KLGaLKtsbCAPE7bZyp3RrNa/v/bYFYpeNHE16iGhLmO25h+/rWkmkmYDzsPxiHRIOhVXYW
OpZgmgACDQkRiy8Foq1Irkh556OeWmeBaoJo1oM/v0PFH3tI7mY2JeN96jPLx5ISg5GjJSoyt3kC
qyijec8N+D0FcJ68fSEfg+0cQKLKjutdTo6qQvkbzf/Tv1qB63iRh5lyKvAdFAvK5UxQCq3TosOj
TgI2am+gs+mlGZOHSu5RlOqm7V8lUAT+MfhXZfxLntOfzS1zbG4EnMWngSMSZ60fAeB+taWj5cuw
Y6BC/hb7KxoOcrzhPRJ6Hm+9tZJhTTihxRoGQaEA47GKq2W0pq5wFRnzAdxZyKgsU2p2bhRepgN+
xcK6nSiLAWdBNTB7cOHyvlaw/Tht0+r3pwhtO/U3plBrpQgIi5rpKA3euRxzum21I0anJj7I/LIQ
nQQEqtAWX4xO9wmheUbTv2uL3uUQrtWNUNE3vWsmDNmHrvuBuftXzFT0EsbdOJQeBnE5pzMIOo7s
N+4QHMA/4bmQtirULof+AQZLrSxFnrYz3Jwmr7HqgNb4X1J7U4IMorBtsRehWU+17qRH4lXsIm7U
eQMBbyesYsYrOZMutoSrrXYUBxBhdbOWXOMn5y4dAurcjVEeMnS0PfLePObJ44dybdK1Hf2XfY3u
AZYCAQowpPmNBrXuU91NGv5vnxFhigCKlC6Fpjn2J7zPtbFAN6uADGhnuJduJllHEBLPIFQcd3mQ
WHgQkfYETMdCGeusijQsYVBmesBAUZjf5v5aaDABwDQBKASRCwe97vm3bY/5STTwtDBfKJf3qlr6
5wWPuExCvn9iGbSYdbv001ovaxd7qADY+eg0qidQ/HJeYHzz5/IE6JKQvEFuHol5S8PxlcX5B4u/
XJkp6IUmTUEL0sgJsy+x75E2o9KejUzguMEUbZQBmfgJlH9JXYq8CHru6xzni1f5crF2uxvqHWmB
josHr3N2xf5nsplbnGedPXHt9gW0h7j7lNHStZJ2QNF1UaUhBIJgTyvs8iESh2g+v1/P/vEv80m0
K7ZbC1rFn9BRoX1vw4F+MU2slGb+qxsGFxZU9RL8oc25iQuDABVoyfdpa0zT7JT9R/z/KfpYfDhH
R3iXxkFGzZN+Zv4t9/1A3N2u+98afhb1TcSgNoA5iYrKG+k4m5/N0wA+oUCGotz1NdbHx01b7otM
ZUEwIn5QwjDb8uM48URoYzyxsUeOqxra3oi1Cu6f60JMvvDCqV+qyvki1e2m/NPZ2VhW4+X1EuFr
sZ0UkMyIiMwvonrrb3qL2tRxWmEddxxZWWSoayjF9lwZwDeDobyXlJXqRYcjujOauU2ATuMVPYVG
FlAgHjXr1/rKYaNCyYakXlAyuD0Q4I4SCnBP8zgVeMhg9ZC5Hu+i9C6Xf2UKrmNkI8cjxWA/5UNz
49xqqFmvJMN2oqJOLk1VElI90CXvP0c8pbiZQFxAb8NjG4f7cnctC8NwptlWd4mPIT6FM5agXXd1
28GR8FPrmyE2zpkQ37EndBppkCKyC1BOkprjgxWytFwUzIj+8FS6TQnq2vpQGkFr7Y8VDiFoQ5BX
sbAo258g+6LNaNehtH8Icco+Wk+3/Ht1fMCEIiYYZCzOgVZMhFwsSTxQCGMYJvvd7oOq1kA3+LpH
JZs8OsCyX1zlhCzkKTdTi3jpiLmAWc98oigcSMznKpDfCYG1qKJu4m97UKZ6ewlNhXXa/Ljt6hmY
MspdElE6mJyp6N72pTmDBAsL4soZrtgc54rwegLKXPEYY5hqTplczDp+WI3nV/hnKu2A93Nybg+f
ekscR/eVo6WA4UcS+7TeJyhin3/LNZedQpzIGobFpa4fWErhBKOzvUUxdAxMnriEZHryQovqfH6B
j9prcSCBiS/0XqNixNYJRpIVH49JhTkF48UUJcvlniAZ9F8vcrfpPiYHF9wMfWZEwa4OmTmLdHE7
bMMb67eh68PcyuQYijf1UocwLCntEFJW1MsdLg/zCxnYIZ9g+dEg3TnYfxn+RKuYtobgy+uDP4qk
D/BvSafAoEV8PS9hoztXsYmlo7TZfTv/5r6lLuZrjKTAmRrDd+5gTtLmcZ4RcHIWlACLXC39C06I
tnoBkDwHUsef2HtgkbVRMQpZJ7/oG+5w+FpyBzRRsnYR8q/PrOSOf7d0sFWwtPXmdFQaH9H0wiG+
zRWxsL8GR6hqHZUoYJ/9zTlI6uNJjw9+LSTrZHe+0rs2fXhnrOKccGdkFYVM5kfagyF4Vl1V+Pt9
iNf1VW53rYYvT/b3BX/IgmCW1biq+P1oaXK/SoMX+yVkE7cZps01JGTUTAdecvajCl3SxZnTo6FO
T6JlIMf6NekOCDtTdeFfVmKPAT97EqgD8IQA8UhykkmxB2txSLaBvFLZM5O5KynGVWAaf1SnNdGQ
fCGxEYv0fqK/YAepKiji9sqXr6EN4jk/4CGU3/tXrV5gOQ6UgvyvFPwnrgNyRKdJhlICXOFiRsfK
OnPYEPHuYOT60B629wwNUflk5yNJdPvkdb/5Rct8VHdL+SYUWu/aXbirzv6+Fl0zyDm2pVAgPdfo
+2lk6Cn832JwgKggz/Da7NT4IjdngC5WsX8yBusUjninLJSA4aOzhMrYHyIYd9pPV7b1T5Uqf2vj
6pK/ZSR7yTH8272zTNn4NncRbmwW5/2adc7EngetzXiPxeKcLFM8aqKPf8gxMJdL7roaS9VEJ2nu
vkYrISLfnpjyQyZG5y5SYOXpHA/bDR9xD3pJsWuUUiWQEky5V+kfIAyGlrT34jq/FvZ/nhUIX2vs
y5PlgO36cJruhMY8vCUdSSiv6DdavXPlZpij2g/pZMPP4XiTi//Qse6NfDqEgHdae4iyJBdsuDo2
PT/IxcAbRHgNOsaDQZ7PawHcG3edWYgVtPcq4sWxHDirFYsJmdaiSbUzJOHOOu7LibaomK9BRWvt
L2uAbXxj1Ezd6nIbPWZRZQilk6vq30sZAAbJLufs68G8JzxB9j11aDWPDQ1UEo2Qp36YNWApAhc1
2aQIk3IW87CVq7KNtaQVqf3lLSctexXljRhIF4A7VXQn0afRLaKmiHt8MLAipCqfs+pRoHUrgXnP
J1drTUmhZZOttDSFB8qAYzmMQzPYOJfK8bcju9J+DGCoPski4MyNVQq2Qmm4SF1pdJdM0e3cbj7T
2FbMZ/6UYz4KQ0HzVdiVmLVbx/Y0EpQ8NFUcnKdgbzyABltT870C6EvAPr4D9yIhaOL17uxu6Q6D
EYL/SuXY3kxf5GlP0MWRu7BLWug+VD43MaB7/EBJoG476G9R8LjXzdMUTWQGlEbchBohM1gljYIm
FlIpSs8xvNmt7SYjyvucdaeb7CWDLjFZghhO7a3W5Ravae3o2ecB81rKfcPI8kJzKPOEj8eToQCS
spDSg6m4SCa3pYg1DenKChG+yT4xiRsGa5yQqmzzAwXwf8mUB028CxvYa7zGjTRQ2NKp6SM6gakA
j0J1uL5UvJk4Fj8UDBrnT0Pk2O1P7Xvgb3Amao6v+3TAcXR829bxEkOin8ZmhROkXb147P1ep1zv
WINUKhoGaoWjl1PYGct0urwJ56C6Ksa9hoff3ORcvN0OzOujy4Dp1yaNkGN0cVpctUL3EreA24FG
332g4v9JzisgDlsH5ld6dhV7ntg1aD+mCvHqsua2JUmjdj2ojmZcHIVuiWjkHVgV3EcS3jI41KPM
IRPfzEGO2OOolic9wU0jS0I92ZShXhoW7d6EmiyA1T9myja0GLDmFiFO3FZOQmuWbJS0c6VlJaU7
wQ5L0bsqVeq+Cv2jtELyHqj6XHNsa24uRCxnnydLgz6u8NKw4lOfZLXwO1xc4Wk7IujjWQfbCNHs
f9AZBrdEJpfwL9WcwzQJVQMJ5HfSfSCixqdwxUSr1KfwdHjwXo+5ifubQZ1qiZzLa1ZkKyMOHkGS
TBQtgLJwbA9nrlXxCRtmnkAPagnSFsBMH+ROD2++Y6MAzFFUkMXB2KJYlB+9jbT/Zd+d+fgn0Dzy
Hr6WZm3bV+mtOy5IFdu9mrVsAmYHiwjV095I7VUm3tqGiw8D4xtIamIcakvCSAHw8lOh6vB5VVF+
Dc9/MpmrNY3H0mHe6pukdy9KqYBDIvDyBWW7SXKbp7SQbnhvp9IoLGoe09aXE7pnj53gqk9nSpgM
U+S29Ju8jLW5UCJYYG/Q/VqKzPV/5GbxOe8oXxWtp0/wDP7XoJEIJ1P+dNYZRsd+kLNquHj96kVt
YIXUey9oiGw+Xld8AWajUGUaEga5tVKjTNd7Lop242zT6PPUVp71TAjZl8U7Fk6vomVkY5sXU9A+
iT+Zpe7iAOOCYi9Rd/BXnZaTpHAJjAPwPLPlbC1VF2NpetIg/7lg29A45f+em3Pu9f+N1K0V/edP
fRWRu59J8IRjcjf7p+7rq0xoWRimIRoHAZ2ScapmQ7Mve2KdiUMm28JE6gBu1MwCAzBOHBtMXUYb
e7VB9hMz1/D3JnWizgVHzlFh0ML/ewyGaeKFAfUYEaSnk3Se797CFm606VbX00QVE+GwEc1TO7s9
yBPFHwZ9892cmRdqPuo2D0yJQzjuMaaek1sG6oxq3+/DUngfY+0YZub6OCRsGV6FQ4KbKoC+2Xz5
UH++OqWEWt0NhfNmS0cmQQRXCWw0ZpZRYKygbdQlOxCf92rEA9xUtOH+AbrxRqALCASHMLeiIChZ
LF5/9lh9czhGpXAT+56ddzGViYoT8iWIoVoYb5o/17nFEq+jqR6JKP11UOe0Qt6Innurskb+IHAM
6VTkwwtkPSUXQrUPbJgOE9Tqym8ndnrhnAETgPB8l6Rmz3qyCe29eRtcaFzYLXHKJJ/Cs+ncqq3M
ToB1zcqcIoGdgCNi6eSb19Ai4NsGZVOqkxca517uh6x9JO+p33BAhzs+YxiRLvOUrFWNceSLRbms
4BCYFr4fhA/tJo6ZMdS+xZhC5ErW3/qrKviU/9ZUOOuCM4/15QGmvdKyn3vNX5BQnUq9vmmbmAiF
DPJyQ0vJOwSc0KTkyxn0ASkt9tEEoEvnNjx9KPD4MB/40HlHGrhGLj7cFxPJc8/DoShdexIZ3x8I
vAJadF787R90sxXK9ZPRYsWNL5TakqEhnkoib435GHYLqCT2VidoepUWHOBaacQrLJgolgLpVOmt
XZuT8nWg8gGXb/nnZy3w4CIhYKH+Kpo5v/si21NQdb2g1SE+2ru3yjwRr7xP8d94QT5AhkreuRSk
C5zYOWbQdVoHlfWqXjvIyOKXb073F00M1vGIkw3kOJ1zUbT8zic9wdj8C5NblwY7ePP5ccAT7fsu
/11637AydMtEjEHzf0bmmRq9jZYDdgnNXwUvoZvfnxqT9RAT8KKHtVNo7JgZ1lnS6T9U0rlL4Edu
e0P0xittHfe7ct1cjlcKAdkjezHN6Spb5jyHjZJs2fmLdhpbXKsKkHCzI7GapW0YE2PweEZNTYGQ
2X12LU0CrhBtBP0VwMLVBhUvYv8riMT3If3Pgd6lVlXZuzafreHwKZBpRW8wcS0slErUwGCKe5cZ
AjqNDT89jeQhvjpffqtXNn7mT8IEIvmwmadMCzrYsCFMEgwOMzC7UMNKGu4x9hgnMYiGd+m2x+Q9
uiwQ7tKwn3VbXH33J5UEMNI4R9rJahyvKT0x9fLU9r0TzhuYCAnmbryN574ks8wnXz6U8fVNqFv5
wEUpehKC3VXVvTUf3VTTy8Kavx0ROaHBPvwjGStI842Jo4WAiWVTegD1Fwe9Joixh69aRlRPBVi8
XP3icRgSUh+nVLJg7qLjj1Z1xDXSyb5SE1qVp6Q24SQ/oKPyh0c7pGPFYIT2cBlT3n9l4EX5D5GQ
2pzD2qHyI9hdpKL69K4ApsjPpMDzM0TiljxYA+Lt9KiF6JYcrRfZCzP3Jqq85ytDm6/G2H5Dkeoc
STjUZaFdanlNeIpc/M+udw2tLLT6ZDhuVM2K0YwkeC+83lAwrq3guDirN9ecAkGNPAoucgacbFPG
0GYgNBuVxufYcEmsE9kLrg+eISOyU/RMRt7mJPsu52EyA7LuRyblhIR30BNf4KHyTS9nHl3ENScJ
q5SfGyivhiS55iFK4Ba7Jt2J//HWVdnU/WbPG2E9qEIBfUfPqwJ3stDyeotfkZ2lFg2I2nf5sxSC
lGyRbIKfwKZdhWrY8YVLxUF8od3C/8X8amtiwuSi5rHv7mo4fn8Tvz8keUokpdxv7iQJqgsaezRi
3Q4wUZySzqEp0vlvUUQCYWPn3JXZK+w4e4dlP6ZSbbH1kDPrePikYqT6grkDUumjZZ+P6X+wtFPE
y3ngQwuo4Pif3ognDng4Gv+Xbo+GCTbCWqKHRcfCqJuOiUcF63uYsuS64Us6eqKesz3EGNknuC44
+nQwjK6f68QE9R1uDiR2xMFQvPAyRdRfRZChPcWBJO5J/EU6kNhxDrRJiIEycpDAIzFji/7r92pW
hvt4xFnd94o34PM3xpXprfr1rEgvGt1hRVbTW46v+ZGmqofQE6GtPJ/s9xYDW99d3vdltyhVah7r
nuT2zwMKadmD9mlAMiAR1jpwV8qjDRbYEl/tEdaePfEC7iDIrfCRipmlnZVKLoMnkmI/ER1rQ6Y7
4X3TfbzSA67wKH9W8TTnxOOs7fQQgob/S7aOPQUuacSMT5lmJMu7lOw3yB4Cn8YawaUbVvfrKtYy
CYlnO4HaFrUXh7OkPPRMXvE6x//bC7Nuqct0HbrR8nBkN/XQ+X7KRd+6oHgIFtvAsQYBpXIWFi6o
zZluFBJm0Egk0lQ3rB8vdjPAe9FezkD/tQ7IO2lWUewY5X7eu7hOa8T+QPjlqtJz2fwMv59bxRxt
p+MhVjzvwhTCZc1/O55S5bkO19NmCpP0giNXQaCSkIprZvSV6jILo1ATVgMVi/V1GigiBw6uaAao
a6UTuxxkZ2rCgRiW2D0lE+eWk9MmG+7g5qmw1+6Bv0sMDbsBxCuMsUdcVu2RupHdFqA4cN8W0fdz
rYo/55tKCMuCkD9tq+Ty2zvJuG5QxsUQJbS95aETd9GwihUMjM5ab87A5gV6yvOihOl3kt2x+8sK
r0G0QgVrgHmiJjrLweNQhn2H+VWhnfDR3QkamirpoU2lCCDqPp1o3KDJMTOUGG19Mk4np8XJoTKT
drBfxGo99mFbrAub5RKDVd1IhOnBZcip7dBO5vL2qBTgrtvTw9JJYpj+zZ/3y8CO4OEDzYgkYBax
rTIHiKpRa18VL9S33oklcNf8ShfJNI4ApyrYdEwvvadBgNe+ct/Zr5rOF9YV6e/7cVI+xzBJtWZP
l5pmpsB0nl/MemBUDoKKYX2+gLU8UEGQZ26rdlks6MLpe9I89aoHb1VnhxwKVK0OsWLbpR7F4z0c
bISfFEr9Omj7zirmBg3sIbxhqHbbPyNO/PYBMpjVgR24OAG75K86vgcscAWZMbAww4RoJEwD8dFo
9jXk5j/71PchOjNDjeOKjgiBNiClbnzjxsuGfvpjdY/8mX+lrx0/tOPiwsf1Cywies/TlTHV2hmG
13O8DEhdI3iWlHvb5otBNYSnuDQkePp34+Z8gRh3sV1S7n4XyZKd5fRflLNDpgI893XwIE6rlv2I
DRYX8ElwPEqwgaUfNZlmoA+YvVNIrdGxDXL9bjw7yappzeG7fHOdori/EsI0m0f6uoRg0goKubMx
90Yy0Icj7W3uUwxohXROcp4kZ87vtRP9LyYVU+bcN8BasVI5+UP2wNV+pAPyFGkWjxghjPMoq5Us
/tYaTisuEtiiFVYPqErkCqnTXT+7QPdZ7CB8qO0DybmpUjJf/zle+1Y6rWj88l7UhFPnLdog9UuV
NioqIj2sC5+etZwar/HJGXKzux77C/rhEuOp0gKXb5Frmd6jtQD+c6cf+eziItoGOepNdFwzQyue
pdhV6mpwnL/K/aLOJFNysbp+aG/sZlkD2KbZNgVIIsY9k9GLkB+nomo1pNywlOD/iwAx77b2PYA1
94Yo93QpULbj2hJTTvysiLOXhWdL5yMMVBIwbWaSVZlT7RjbOkt69IuSvF9mTAROZnYzL1GYBBRD
QHKKivz5VEfjsFvcFIwZn/gKZax44xRfsXUKcEXgfqoinfoZvP5Dqp23S0V+7RRquRR+QPLg195h
r+j1PpyMRCfnxQgp+d80ZgFJ4rXLlqQmrmR8xcYRDhI+wpJRVzHDLOT89JFfBtbIzFN4dQl9seHm
TXz27P0CM+hBgBkpx353EgmfWorR8QMxHlWsm5iVx4t4JFMAcx/9WQ4SXRyIQTzN6TbFncjHLAA4
KvYZvtv2VotOi+xYYxxUdJj1nF+PGu/ga83ruz6a9ZAETJm+5jlDO3ZLDDNdcYOvayDM+LrwO4Yt
Hb9Qooz2NtgD129Dqne5jVaqCWn9KUkzhhIecL4eM2jE1gxFkNRdzWYh8to814rxA/yRLrOS5y8H
IW6leCMCKBiyiwlc6xRPQ5TwMjluxWkexfRq8wlZKqhAuY3+0rBx5jwib/cCif2tQWzVP9FflQ+7
HAjJAkn/xtEAES/k/7iKQ2+QmNPgbVmW15nkx7veqvUQNADB+a6Qe0iQkf2aU/BUaj4Bb8jnT4nW
MP/LRUKVrsc0DumJiYH3t0WoWanSgCr9qXOs7wR2A2ald9eJmJpVUf3UNNndJQQFEuVmfeVxeP0o
Q4wljNGkJ7vCtOHvkD0Dx6D1s1mCIm9XpXAsjmayDAsjw7vUgOcdfDiCQB+ad9fDR4kcN8zd3ezK
dH3C4nqJoJ+8PAjucguLu+sDHqrrjIGJ7IngecFvTLuuIjYlSSFJNeIQTW7EhWP4HWupTHem5+nM
7HjCupzak96b890WVLXS6vExhoAE4O+1uRawtNQ6pMBCib34PQL1VDu4wns0J0X7J4sUcboQFci/
AsvfnlLSzWDtOA1OrNH5eWImvm4DVkhSbJJ9x3I2lYjwYmotAjak66CHTk7ZDx0IPi//Q1/+0VCJ
nQHPF6nJvphaPgFLpzMn2n24dsT5FmYaXDi9Yt77LCqquZ7ZxbBsgVkZCascPpuSxMO/Ehd65b/4
872LNB1lK4rP5wRlJwloVqlS3s86Xm4E7rENoTN15RPbt7BoykvqjY92Nq2eYnAH8hHM9f7EBAm9
IxnuLDgKItVIjBf0aP4jL48aBQIfR49MCLKuSJBLbpuSUBCrvoWqpHKSSnsMoMlmaBPOyuWe8WnD
zpzoBcLwxCboaLDLmatgRbbtVb2IjuluvUTKkVaEpnLBcrEgmKgBC4QUcqgLtgQCCtLucWR1ljeh
nJzhz90EeLJ4WONX+z3bYaXFvmA5uB2kDtMTui4iX+wnmdD/dv7eKZIAtyFtOTxm/DfWq5jDwmEM
Ask5FNH+22xea5Kf8P1Fa7VMkyV1whmhdJkSurwRssdPNgdg0ZzZYpKI2eQblO5Tsro3smpPWcaX
CQ90hqDwxxkEqtH9osuF/xq5wnaTVvy/D8sXrHLvHrsG7suml/wxdbmNcaGxLoAhRms1MY5/nqXf
RfN4erbtGprmtIoHIyNbsHf/kqU+kGGx6ibaCZ3zT76eanPfuCKPr17ihzwDJ9vemRSLER1VcE/3
77JYtf0J92UMr1LP8dVaNNNgoiAQJ8iqwGST0vQx9OaF+blWAin8FPOgRBONXFXPTuiz77ifA7Hb
3zikM/1afEDUMbWAKSVqRTAjNiEUyRP4U7BompGn70xycrJrGTT5A65PILStGi/s6+aCJoGcszaZ
AiBIO5JMwPhPmDffuFQmeU6jnAzmE237w1qZrYcl+w7c1CELxbs8SFQ9b15XY7kuSkZd0TWzZhJD
KqC62J4zndusL1brMpoRPXJoDwGWX+Uj+4txkV5U8d/GZ51uBNH4RgQUw1eI0W5BUXK/pyrbyu2B
0BrUy2A/xbD5Gt46LVqd2ONJUyehkiYLftbAOHAGryMgrOrPrXsj+NCqYyjWGE5Hnv7YjYiChnxT
TAJ4C/DkGxus4Et4Fg/15FieKgyVmQ1r8Hzc3lcVtoiQrtRm62jQ4zdy/c3k4dbvn5FhCf4m+IFr
UHWbqJMedHga2TUnVLSoCQMxVNiMrNxcdFnOdD7aigxJh2wEO48Ryx5BENq2vYDpQVD6gWGZ2i0n
MA59NXa1r7LnD+pj1I2ZaUZQg9Nhu0on0zwzReg/YF5Mt9EemnJJcbxHS9wAuAhZNFoY0caMm4jV
4S2/RgILC9DNcBBtE07qnafpjQr9CaoxnPPqxI/OP+BM/0nAPtHzzYwgLgjoktwgb1Mqpkitjsoi
V6SM2wTyRBdmNOJUKPNp0Ld6FSsjhLNw64HxeUCaf6p0tdTYWqE8kOHd6NlyLwsYGXxDjR8A7eWh
swTipyRWQIEkShclR9vXO1dEABokwgC3mfC4fHOQZe8ihAwxi63wdj7GoaJVuIgwRXLyXfWJlZxq
4exPz4LcKffNK57Z5dQA6riZXCRbvvh8e+6NOY4MXotuLkVqlT4iDaguTavb54+mVc/HvEvJPyVW
NasZD1kTKQyaOcxkjRkVfsopshEBTwPDspMZbaZVWmhpUmzdU1fgOLCMdgGHKzPtUxqShRlVlyUc
7WXX9TwOI4+qWrNG4hMNv753mcCABI96pbk3IifnP6mxC4x26KMSGyUi/q6N8oxncJHuFLhoW6SH
URVEDZXr3ELi4xPfnw+61myyACaFrGQGTY6S316S7AHkkXD56dMRanbzpIfFiYpRcKcVANkgFNqb
UAcAGC9koZRnV0nPQwvWkTZ5kIbqeAB4l1XLJdaEfL2UwRuN5urLdMCQF3WzkZJDcr6LBXhFM8Wz
NnSCmy+F7ojF8ulueJ4aK7AkTNUhwQqj1n45c7J8HrgMZ6Hly1Niacq0+VGGi4MlE4bGqoh6Uz4d
eMlro8VEUeDNCygp+VJJ7QuC5DgbIuKzfe5G7bC4hV0kDXx1Xvu3FUmu6ULtljHWzB+KJC7XwCYe
+SqYRJqCx6+E4QEbKmOCrG709M/FkWZZplcHrDqmHsj8fCH/+U820UqMc88elVzCLRm0ul4YGWr7
UV0HLEMJdvB2On0UgMjpx/7TJ7alKN4pSonhFSxz3o8WZ3GNGNc2Ea8sQZXhk4EzpyAbdYIBZU9j
U/4jnglLg0K1AEnZRGYOvaHqPG/H+9ga2PM7jTEExy78tqVHPjQtmz4dzc9SCoVcLL3PLk9oG0nc
90srXR6T+WOIGyVmzyzbB2uAJ2kcHNPArGWGTVTpGuZS6c0EKsk5bzGmFxM1i6Ek+TF72FtIT6EJ
YFuwpYpo5e33vtb4CIDBahsw1c05YVvtiW+oj8bdCkc8D4VUy/X+b56W/spZktdbENFqZ9Whgosj
btjZBIzGh2sAWg8Bqv97iQNeKEr6fYwBUi+7aisXKsN3o0rkuiyBF9E2fZQ9/5kTRIW+RcyQlZW1
70ziPO0rdlipXxHzg2Yll3mWXp5sHPQ1GjzUm7XeHoTvjQm0ZPi9Zhnc2XGnBl6n9cZr/WVASlAD
8kJD4Cg3of3kqiyuvmDd7pX9DZgPYsgkfAvSoliwZF0P4ZEgXItt6GG3J8h3cvP0jpUo0auJ4ERJ
AFWS0qfnnckEMKJ34WVXbuRG1xwt7qY1BIPJHOtfzqSXD/8vWipugnzRIH4qeTgYYhi1FULcAtET
JiW0Mo2wdVETRtf5hwwdc4gCZB+/9x/5WBa3VyPg6zAUf4u4mr4CJf6xirOT68mh5GwTK4Ae52CN
IlK6BGFbGNAjou+Whdq52pBajEulb+xNweZfYRHKbzmVdf2azEi6hn9mo2xMrMr68fcYE8npvbyh
9pUtnWDxy8Zmm+LXaP6TlgJJC6RvHiLefCnl6tj4I7CB+ulfVzQdaBuWw9cHB57C5Az1WoDww8or
SGdaRkLIKV53bUrHT5NUVlE/HhviBtS5mRJsTN10o7cJKC8q0AGXgr+0RccLYoWE2BLxomKPswaQ
mbZH+YEonshshuMSkz9Kz42ca0Q5CywwSMzBnVMFa11rWMhEJtYWCovyYuduq4prL5PexlajpoHJ
Ckvy+/QE9U9HSFkna8DZWxfBXcELp1aFLDZN8hU9fTgSTcBeE/6naoFW/tFlbMXfCVIY1TfKpCLf
fouH5duf6+o2bzuu7cBKhZJf6lwrXgPVm5rREMRlNpmtxeAjljXU30S+2eXNYky7ovu/L7xZ+lhI
tBY+vcJWAHHpCWUw3wRjwLKw5E77W8MO/Ts6P4H91z9KlUULkAP/5UAnfA/JfAkLFgvKOsifEKK7
cEqOuJlgiM4jK4vwp8pG4WvK/0ePsEZcI0IDG/OsZq559ZFdZtNzgSGYv8NZjGCoucn+Yi6Nt/v4
agfzaKnwOTGbbADyDXSCLiam3JdezgYBcp6Lbugr7Dt7nX9YeRIsHY8t7vIEqZKMdNgc5sXHGTys
er12btPZbqiZTdstRsIuSpB9jOZofBeKNgklHdHzc8M/3V8MYE6xo/ox3CqOhoW2Xjn8Xr4mKM3w
zuBUxgUQRjqNgBlsJK5nLkV9E0PK9i4102atUjNRn26CK/FwfzJpoEWizV4nGAbAVRD3mSPa5rkA
X7l5ABzbFl5QAr2CBHzGD/QdOo/hfRaiumxW+nuW37UE+jFhd8mXehcVUq/eUJrJoQQsQvfptTph
63Yp9NZeecWQY1TcnKSpTpG33lbD7wunsRiHLIhIlJCZZRt8nkO4H88O+DIHnSb9cnMHvxlREOL0
tigGSIflQSceN3BX8sehy51s5+wxAViQOdpanVlDkq4Kl06SD6GwCDUUihrQq3ejkQm8WSCWeo1o
XLIdV2hBqy5hXunZwWYMOYUSvWdqUkRobG9Xkx1C0axVcKbRAHfFc6IbpMjx9gN4sB8+vNZOr4p6
5IExVQ/oO7ExLH0r6gXVa08KEEmoT6ey/q8Pm5RKSJrJQ3L0EMseiyZ6+QkCbsqC1QIHhiFr3Rtu
3rw87CvP5oPnNgYmIDkQC3EBRkE93xlhGRCQcWnfqgQdFaAcDyg+dlw+up73OVXXmcdIVj/wMhWP
Dr+V5fSMKWArWLB9GRsXkU40wVoTmuVC37L2+55BVAm2WMGuJ+H2jbtDbZ8Wu+9x6yPHkZCjk4Kz
Cm+lr+1P4meX3JcbhTxdDdSgLz7JTGAtVbN0zPJd10iDbdE2X3c8bnYrtSQL5JYIoHujjGF5pxiM
tOoxIVcO4SMhd9Us5q3K/y8N8GfCk/f6csbC8fjo++VdeYgZgS7q7Jv/r8WnvLd8JRLJzOqBsS1e
UHQ14DJkrzKz9df0zmZJqI6Xl0mz7bmnlgkV3SUS4N13fKIOT9FtoKINqyj9uLIamu+kX2IK3EvQ
I+4MKrSef8/HZerN2PyXCRGxlEW0P0PPTvSky7qhA+AO6a0oZU49vqn+TaoRImlkzFi5nEwUwCKm
3EG0+RgjBjObZCc/fS10icSIhLHvB+P29tpNAAVSqEsjyDLxnfYmoq6XYX2S1v75743GarHBwBx9
9MBkHYXkDs/l/IP8Ym1nB329QzsqLj63IuGe4fHo8zNde3OnqBZrDbAXFZlq8D0MFKQP8Ja15Hog
3+oSX9ANKMdFifTRxMtays6ezW8jJxFLquG2sly3GDjjasBhPXhWyjE3YgwLoB8FNLjoL/Vce/3Q
mqZvcxwpoYvTFaMoySsNoMf+hO5Mj7GrRaXLYc/dW7Hnpe6Z9mk1LBQ38/DFxbTyweLGjExXZ+Eu
4I4GKP8W5K65VqTcv3042kllq+c4zMmOdfo4diygaZB0Blji2kUSgI37QXYa1LeuY61PTdejrEzT
Bci+6JL99SsXz3zoyBF+yEehJVm0SQms3ilAMphRN6E/eXrXABFUfN62uZ5bKLVZIsV9jMFEuhCw
hEnT7z+naprH4/YBa5x+U1bAeCDpEAC78SdmHfDN1yY+X7TYv3eliPvDBGG06FrgBZWjTxjEKhuf
Wk7Q7XqMmkL2wa+PDQZ4PtiK1spa5MRuLG5JcBFnQUXQTwbqUqiHvW8+zQ7v8Wv8UPXxIXGR5TKH
X/isw66uJztUJlY194AoZ6GcBV7CWEvFwq1iftO+MyWGtJf1bRzfb+M0oIkm0tjPgymkPeM22rWi
1M1MzCvg4zWRlr2c3rqEk93FinLZlql/9+xIsxGZQPiCYM7GBKYuesH24akEOqle9zvSpQelMR5N
6QNaqCmMWBGy6Rlf2m0HHh9FTJghMrz30VX2aEZAko1kC1bjDOOppd8iQSal3qMHAoc3oFnDhzZr
4XtQzER89B26cbTZIHTHtRJbj8MCvsEJ1/WQkyoWx6q/bcqvHUkJ3QcWVUctArRIQs/gHPShi8Zj
GRFmM9tzgdOo1bJic+wvL/IQmP1T6noKqwZuDv5qmeHX9J8cFLSZt6xBrGnesmJ8FizPv9Mb7v+e
SYVwa1jehmsAUY2zJWQu+o7phBxCCDadrOOsnv0/pkh9j6J4oEnmxj5okit/QviuIVzz+9Je7uDo
WTD9UXe+3fqG6qDuZWik93Jx5KGSp4hfMXHmjJMrieJyYEM8t0VNC/lPHgADYA/YGDAt6c4dVUFi
M722uskxdO0KM12pjXK1EYY8mP2RIr0VWbrBfS+k1Pta3f1jO41PZ6PCO5GLAWbbYMUkxXFaZMCu
iO+HJtsAOQF1CkgBSIY3/f/Yrzr/zvKuaCxcZT3J8Zy5ttPP+3IL8XtQ8hVii2NcaxO+TrZxvb+z
mvTUdibfp79jYcQ4MJVlJfPI3YmT2nMzsXVJ8iV/Hyb3cv7E1iltStp04wBBUr0DqSU8ANDU9Nzr
FdxV1RpvVpZ5ChNITdR7iWyXkdaGW4wHtW5W+9tGhcnxHi3T/TBBGWQfOlmeoMCpXZGFkY7gfwbI
uUSIyqUqFFmu/ya1ZWaFDkXDBcfrDDN1Az0D2bGlTUwIA/2SGmliXj/tH4/epE5tb6wt77Iw1/Jk
6soCwKWt4jcf35P4jcRifvR6jYSP8phYIrz/nUNGC3LsA69cFfeHttXrQT5iQYtWwhq+V7z084EH
r+MAmTI/GyRhuS3H5KNQEd4Zj0A5kTxwMaHN+bMIfbe8LVh5ZN9GC+Cf+IlkoqebYl4E1B9xRwsH
Ad7cthDKb4tJt10jExchPCDdxqoBbzCXrdo7If5oeoWpdi6Pp8PnPfP8reRaY/Af9YSnBAQhkPuU
1jlkJYDDOdG6LojRB84ksh9PNj9ogAnVLwhhQSs9CHDlP08wvJ2lhR6JvQkWAeQDm/vvIqKuk3LU
mpZlOo5R8Naclm4LLS28D4lPfkl0vsHjlNbHK4Hse3J/uV/9DFh+z1KyIc5QO/xgWfiCC5EYMnOj
c/pV0LIM6WEeAVyVz6EKFPyizmKrbJiAQig7uFhOcvY9ZnrXx/weKutMKFaBVnPFbB6xgO4Sz7Ud
sarL2rOHUjsCZJkmFCI4cQGP8xhvcFmvtgmoDmXROoft+Ip9oVpROZe404n/mXGK5ByBMZbf6Vv+
lljx7cE09dPDmlign6Bn2gVOdYzUa2EORGi5PReiD2JR047Ic8/CHQnUjJ+8HYmsbzgkhTQ7ANZW
mish+dfctXcrzDQODBJK/CT+DeKMDn220g6EN/tuf4tGeqoRpihTQ3+gWuWodVSBmga1KxCeirpy
/zwq9IF1c60l6t8jiQLjOMigyhFXWGqaQLw6wbhnCG5Kjl7Rci//xMWnwGejECNbACIU7PqC3CX1
KvGRWZkxxv8/iygJzKBaqlEF85INGFiqg7/U2ch2Ni5I7xfA7R2gCwNv+5qbPFAr9SeyvsOumE/w
ONTOiUrGsSRSzu+6jPI1Dfd7fCqkIcX5/oNyQaQBfakAbLbz9SSwW76NP12tLHpq2qPVnHtApbZy
uu2Le8oK/qIqsHdzNFwLIA7Pohmw3EcOBXgL6+6YqOpkubASwTJypiiKznwOfLRD5wVEq0hPJnOr
nSyP1bq3hUqV2tJ3V1kO/9T7rv5X8N0LDqPtONE/NJ7SHf6pmIz7XM/MPAMtBAChSt2COngbidYu
F5OMuLpMmBbW+GHiwHjCrvo4f4JIXUzhfjPM7rS7ADdx8hx0BP0cF7QlGVHyoZupzdWMKt7Qxyvw
mzUQcl/ebStGpMhuVSm/QmhecT/Qr8l7nw6nK4EZbBCUOH/xDK7N2/h+e/A8d//5V+K4kn+iQWmz
0qJRP4gojCJFR2iPW7yFVSn0QE4dVwGTyqs+pyc812yEzKST5u8MW7a0pIbLzT/BEZ/vyY52Hxdp
eqf+yfOrtfhA5jg9siSgHA34P37AdGlpShNQH/l6egZifh1vq0Dot+47GaB0czl61KXXRAZMTyzJ
jCi8qcTrq9uO5HHx//U3j504pJzQyE68WsFGRDcUNUa47/7QPvEvw3g38pAaS+0u0HSlaArs2mkV
LkuJ3DlxtW7TKnEvshsXRcI2pEVWzQ/c7h/pzZRChmBf/RGEMDaXjhBei+cKnV0Mrrjg2attOW4u
Q5AqlWgP0Qrv7+qpfIGKVfkmS+2N78A20XzfYoOncx/mZzC0TUNR8hci/zm2UUq5bFz8I/v54bZT
Ki1g2fjRXfpIH7tqUjWOu8TldVaNt8ivGq9gyE0Hpyb2c6aQgRZxD/7THkr1b0SOWCNsEpSU19SU
6o7bJri/StipEFds2wTCK8owe6kf8HSe/Yeu5UwhwKhLfI4k5xxd2sykLJ9qPkTQDJFY+5JXKZ49
vpqZPf6uZ08zrmNpwAYEsSRMwBu8kpH7oU4fCx0w1cjH+OqfDA7tlQog5kob3XmkXzy2Cuy7glh5
8GGjvPs4YmW/KzI3lPckvLfoZIgnJRJdwoGKN0/rjEG/eC3Ka5wmW/ixMk9Dx55uGnfpS2L91HZK
x9N38LN4YvtrJakMNN2FQLxIaSwTgT+CW8LIfkiJr1KgzpE0Xwjnz+IYuBwPBdjUoK166HmY8hfX
G2pvNbLfMV9IAMXZVi5yXxGjYYvUWmojORMHmGNHuqQrZYGV/NY0N2Xn+v8PlEd45bj933Cn4OBK
uMFF/Dk28WgWY1pHV4nZ957phy6MAnRoFetyZlhwu5Z5NTmeeTyWv+IVAfRuGwVWBRajt9rYvVGp
/X55+gKv3ghYjdmq5VS1okPWEV34epGELnNwBN86fgxtusDrqQ9LThgnUYESj4a3iLok92IykS5J
H1yNK8duW8fPGUvxObtC1cdT6EOIEkylHdCel8rUvBk7dMJojlQrFZTPWs8pODlHLNuUqZyp8aYN
fmEVVh1VzHMQnR34+dIFRNu/pm1mS3JmLpco9RB9NprO+cX2G00Zg2U9diRAV3qa3hCMS/T2I+zf
j62UpZvimFm9KV2QEo/DbQrLL/baDqqkj7nZk4VfoyE7GHKC41GVMpAvyfZoMK9K3N7sadooWrXq
Bvwl/3Z32XGIxGK4YfuTqwSYVjR4zMBOkHsEW4PDNlEQ3YMBH5DjcZZDVrZnTSh+Kcl6w9lHKUO9
VlhjPahDsKnFOVyZDDG3rWBd2eGvQE0aI14A+/MNz+wdwWVOU4hspU05H8LgBoMxMuN2PYPrV8H/
GSqHTPLEf42tF4vhea0wxtP3uZXdDt3m44Ze3GElIkqnfDXpZB2Z/iS9e7jMsq2ObzmRQHkCQGmS
yNLyf3C2FK3Pxp7KkkJwdM5AWUwUhxK5+4ilPK9RgPNBNXGAYIq7h8NpmlnONfo7uhaOzxd5wNnQ
4YykCe7UverXgvwuNWLrsGKxGE2kQcP/WWP0QGqzq7DkLBy2+9VOh/GqcjxyNm30n9Qdp+nPlmgT
v1jEyOTUZoKD99cnC+xOBwT9zgk10lV9IxKDNqjQmgV8uIlTZ7C62MbZzbUPRu8XTYTypvfb+Ed5
9Cp1GLgp91NFFXBCNqlZ1UQ2SxMk7+f53/889VCamcAzZijYvf9GUlZwnyikpKZXgWdeJoDgH84G
txpMh/RpPDzWBrITxWwcbmEgYATRZzM8VNSf2n2YWnBjI6qPF40yZuM1a5712lN4617lFi6RDZTr
R7ZWt4mglt43KoViyZPA/BFlrP3crHlGbTWomP6PLfs8HgkcUAE0mb2u0G6bZYLCmtlLCRUdVt49
Jnth6aCybxu8C28RJtLBsoKRQribqh8hrWJR23m/XgFj2AdjNtWwOIeFWff1GG6ozv7aTH7P6USJ
z2ovXPyIXYpn8CZDwSZigQFOhMSIiVJGkYbNGtA5+3tQ1RX4qQkeJNaeLm5atLkQ0hUHT2l8v0hR
ky/YtRuyd4XKwr3CisNcCMsmbhSi2p7sGHR66vgzdOYJvNE3f9/IDrSl8+uCXPtqe3gBERtRp9GK
WW7Bbb9Jj5Yf8gBJz3FJtM3Rv92xtH7TzI7J3uxoBo3EixiPZmLk41WU/ry9IT21h0zkDcBi2LXA
5YHCSh5AmCA+hKbTFyQV9Oz7uA0/b2GYokCg75ZpGgRiJbuEv2zp73P0D2pd3bmbc+kRADg3YupE
05ejLe7Ph4vTBDHkkcC0DwS3xWOZfv0gMDmERPEeEjfJulPzIMyEqo+bvgq0bpM6zMYS5L+dPcyF
979iCAjHMQqd+aDMjAlAeTRVmeN2jBhTqL+QnxvAShpkOPG5X2cIlLWXBVuAsoGfB+5Z6C9UkvJb
XIiTRHmGWjPhW5I177XYjuj3kw08aGrkUVc0KAggXFapX/j+wqzjotxb69Q2bQavYOHDsj272c3p
Gj+9tPRheRyKorge+LrPNF8lphonQeEd0gzFTz0WzKCapfrsu4oZH5LMTgCB+p31oq3wPYrXSQ25
l6uIiuHg3M/yRpGFnhJu6dW2LBPLD520eyItZ52hd4KkFTisJ5+GbQJoHFJxJ6Hmzz8+Owdl2OVs
Y8UZo+pTEeIRuOv7gMtVBaE1VDccdE8uNg5MryIRxf6gi+NiXvQekuTcaFRLFRtnbGVypdk8KdZ5
5pLwB8YSQ6sMEjUoEZG82nmKHcPeLZ1tjBsqiuNbqXlbdzelS0lw/VlNhCClih8sBIlfqt4xBoFN
eJPqca0mUWsKDtX/0Qbat05KhXAuBC77YQbY2dnEYGGq08dsapT+snE/07dRKNlL8fgUKmQaSFdK
ky9RsppV3zpEKyxFKPiVf7mbBKJ0mS0AfTK63vJf88QlClcL5kOJef+4DFZiSbRjwHKajkR3qTwO
VBcanqtnLh5nCK71XNQx2IxoQ7yNDa22DjBI2wXmo8PWk4qEKTYgqnvnpj6co+4VC0JBcHgYXP9z
cj/wdiRm7djt/fdXaqTw6BdBThShYOQbEtORH+BjHfOmUy0ch4UwedHRfks7BeaQM1uDnIBN0tr2
whNFv1q1vlC4yDGMmcXmJ1+Io0d3WbfndhPhnYYCVdbDT0o++WLeSnp188sZPXbzEw9LM8VDwca/
VMnNDz18r9VKokbhoMt+z89XwNMAOfpfjvZo2O0aVqLasN4L/gijWwn7pswWZM4rhuQt1b6rH3sc
ssLKXRsrjbyhzz7vQ52xgkbbylImQTTCwpEx4+WsLIfwUq6X5AgNLzBizzMuFyLpJ0EJ+WcuVvex
h2I71xmTGvaWsrWxfFMtT1HU57C+NEbYC5UeINtIZAoC2Qo+bB+Qet5yD2tkTaHO6iDKxdD2+lkI
HSyAiISyBWQ2NIzQqRDYzO4NPJUQpN2qfEUW/YM2xLFazOvHqb1xyIllNWpvfS604cJh80XmwWdW
elOGSCNeX9w6cNAlEw31Pk4zb6WdEm/9E+FEAFWcLzWL7RK0hcsyRaXdpLZDX+4SXmwGvL8fWfE+
qKlWArKo1fYC6EQtwAUI86LO3eVAJ8fp7DbfMnHTOL1eLt02HGIEeoOOASADDawsrtb0WLBLtJDu
vGbaaYumdet+0mWXByk28yjhGOiY2BMjWSlJ12LwYhjk0kXLRt1Lv+ToQSekZ9vnNlMIcr8XKoNb
dqb1YjAWgkaZpM8jcX+qoqribTpjM7jAU/JsGTCUWDNZIApJP2H5ku9XXFSrBImaUwjhUyGinkSG
TFomJ60oBaib/NoiI7QBuGFOHoclShlVfII3rG64d0YyP6M87SC/keKKSpw/fAcarS/4otiA9AOg
E/GFQr7dMSaPZdPOA7I4fPobn7vB976I5baFa8IIegGI/S8cdJcBG7KI9DcITMzmrROwI5OvhQa1
aEB1uLgwhdh/svMpRJ/ZeSucQq+P9fxvpELmEQHvay+1Zy5i8/vDRPiB3JOH/Pf50E1ObEoXTrw5
OlPBYIdnucmRn5bPgwnUOCPe41tTIXGsn+X4152W31iJvkft+VmDKXIy3V3SPGiU6K5TGRYyongE
fDoiEZXlp/EQFjn79T4vSwELduPVAnE6XdtTdxFew7/2z0q6qlfKWNMKkTeaSUrUWdzg2jM4fYnt
bjfXrqKnKWKxUmMMIyxhET5KDRqL3MHvaQDImP7FqTvdMpIND2uhnb3GuHQULofkrd0Q+p0bmqV4
A1Kss2J+COSEBOD/N081hzJiB5oD2kb3j48y+lLAPlKebyyERiJzB8FxSWOUCG91fVvVTnrI0MwI
7WijLFOKXCwN7hwiqDUp3Sj+1s53bbGdM3bKg/Wn+Sy/Q9p4WivmrbAin+V6TLIy2ssCLDDG+ivX
nQrnB/tuC3rjGjpK9ftYcpbQpz3/RNYYuGa3IwVSHr3zpw+9Wx/zYm22QKdn7Cczz0xk8d7/co4e
tugPY7kHigoZ2BcaqzvDIdPqGGxpidRRYO8Wf/e5ZfTSieYu3uo0zjZrpkO9qO9rW4TnDxSxDlav
62YJsSjdtXovV/JTTNu/LxLBETPJeiaKuqRuk7REllxUSmpkCl4yUw3GsGI0lF76FlppR29d0A/C
K0Qs/N//bUxUhQXwaJtmtxLbilKq6ry/5QZGGMZFka5m0LN16lKl7QctrddGSuYTLBifzUhiXK9k
8bS/04C73ot+IFfW/eD9C7JxWfCnrKi9JGXL2IcLadq6IwgPm69h12P2bUBYP+vQNAF0zdDifvQD
dg5xmLzvX3wyiDd5H2u1j7YATbRU/AMxfbuegeP+Q2T6LnLGLe17tsHN/SHFB8XJ8WQJQ5D93/Zg
3aX0E1nEUs3XFT9t5Ah13sHTUQmNbwhA98Ztqxc4exGnw4zT+xr6vUamBvHHEt0PVq03NF6AGrep
GYGMeTmuGO8lDIRHR7etW96IkW4t/w7IBU5tfUxunSRcfkb7ZGiDuwMS74+fPFYxnCB+4nDvy03R
nNpboPdFG84TMdcbSIwFhBhuklX5pJjgA2fUJQ2F3exERdzxfXx3uLQGjtLaTx/l2wmz5Z4iiNx7
Ho3ySPZhsUR5kdQJGBsD5+NY6pcQnYzxOH2ypSLoxKwZO81FqmJvIdQI/GAjjeIRMiKmZNt2hYAB
+Kzr1n6tYW2yAkgt4A2aAo66FAAfMeNxq+pS01Bi+qaLdQ1XeDj663F6WqlRTiXOCT7YRwbP4CNt
CMk9dMdJBBBWQqsL8ZoFEhaXlqk6LpmO08DYxCtWb6klWm6bPbmrfcxxJq3cUQsTO63EnUlvsfnk
cDS2KsFcGu9sRbrvBrgoH7FBkDlx7FYgcbGBLMWXrA7oEgdomJ6WYPd5Py0pu5zBsut8rB9Qm5YR
ujaI244rgyHlrweNzbZm+fKIXpzORXymTxKAHqYHndFL/RbnE8hs6M9o43RPrfg8fFPUYqtRHmDm
nMmbTzhbWGkAnYIXtO/yC9nqk1r8fBRQeFP/nrg+WAgM6Kg+QPU7INJRm2fkjB4KW9A8+EjmLsHX
AMwVFkOpCXpjedzQSKZpDiQ+mgryyd25JnPFjnFdx+q4P7FZa4YQ4sspAE3vtRaZ8cum7H6d458z
M/hCeE/dnUkaX/rkftX+FYr4ncic1/cQ6BBPOCIhwDh34gUIdMJdAe/pNg4FqkPk6wQDRD2z2I/6
Kl5rykIWtWIXkTa5CJBYO7ms1e7MnFKR9B2Hn/CG+KKlkzrLVT+O3HlEpNaI4hvt1M3glHDFYeli
ZGX7pdl0uUU8szFvsL2u0sRik//I+Q+Gsl7L0Mh+Z+KYoqoZa60gBtVLDyr6QhBBhPPHF5CKqBBq
Nybb+PHS3nbM2CCBSACDh5B3m/uZDpT5lEhdCFjxn2aFHTsnpX7cGlMXJKKcLMIAGrdsW8pG6lF3
MHytHia/s/9kXxGDVL9A4H89qIwOBQNWgNfvLQjbf22RmySrzzi8sP+eDr4ac5ipDUtXKb0A2n85
WDRcXpCn4CgOSdjy/nfv4jox1InMu1WUICz8llFxXqkrxcufcFnLQFaRNFObncH1nhFut9mpVA9C
x63Z7dGkY6RImZ1ZWnCiiW2RWBDuiCPJsnGGn8KMDIlGNNNl8UX0PLGaxAiH7Xgph1ggVMFKaDx9
ei+AJq8PHrulSeTtTdt4rGKDCOgPbIx0DGK9fkimJ9oBoyZDpE1nFfHExkHUo3RU19eI1eeLFr6G
Pa8jFaV6dAWd3UdS74i1zRhCsMtwmSAfzYHWDo7MtunL0wJTFcNoQWfICgVTwR5iu5Jw1zbsIDtN
U4Usshu1x0PlTKIybC02w+ttw6FPl7vneDfhkObvksYm/1B0KFvS3A1sTMoRUc1E7oyNsjTKeWGK
QRjrQhDWYT38S99ojXcd+CNUrUklbyQ6bJ66zm8Ba/3YV/CWUMJ75nOuUZj6A48gHCTdz1htYX45
rcwSINC5nblo4z6FJgLK/IBS5lOOvVK0CITnSLvvHfGpORYrAVg4QZmDoAFRTaN+KB1wcemTTTYf
AogDsBeJVl4HYn8snYFFAxmcB6vwleyatGfG16Y4ZQsSqehBmXs8OR68LhXH+8RThFEGBSB8XcHG
udMmRkl4AwdcO5tIK9JNUsTxtZA5qR+BVGl8rgobN97biMG6EM55AkLhYri4NXMxLEQBLa7erLQv
XXsGhOsi38GFJlyaaVQY6n7aPaG0B0p0th6XEglA58Wn2Iewv1UoDK3F4KN458IrFA/BLzw9bfxm
t42VNBlEk4VtYU59ghV5WDlCsuPApxNZRE870QPb/UDXy9gciT7GaR+l5Bfobiu4oHFyc5nL9Lxt
ZTEvwGmYG5s7RcbnlPmHOBlFE1WJOYjb/d0iVIMhus9EmadNtOxI6DC7dBYWmDPiGrA1Suw5gG5S
GFswFWQI4bI6rrdPu5YUG9KWs+zUzbjr5wEvpvkaCV8YpEdXp6wbsaJ8jTGMIGW/R5JgVSrzyyrG
o/5ioSSxoeWOgVDVGt5WYl2DQqDOmz85ovQOkpbZ7dJarTU8SX3P/HGNkPmW3ZSixapUWA+1o08K
eNpI4odEa5pUL/E/8BQDbaTTwJurX6NXz7UvkZkPw+zcV9KrbhDSUFT7ghuyzgseoA4Gl/bjGNJ0
J3vOO+1+ybJXhI22YIn5s6JWpF97eZF2+R//72YDyFsG3FmzotqN+9cHd6/kJmWYN/zUbs/hrHYv
fgFCBcd+VJvDip1ilcy06yZwlOz/HMjH2dr1CI6PpQD6zSJ44wHXESPgR4ev/SiDL0ggVGl0GSe+
Tv6GsuCmhMeCysmWovg3mDuuZHF3adUXwPwHfS3tZUinNTphHRY3XcHf6J5FADU81B8/uhvF48et
47VNtWtdPsBWYLGdSEEJU3juOci2ofl23Y5j0NDpdHdx3Nl2I7JlKNIL+NpkMLj52r1SZdoUI18I
VWen1WkaU3p9aCr6xnQkiApVyvNaoDiSVL0sc06T5i9us+uEdheTjpv/mB9G/PPIQ10A6S1mY6rw
klprALXcGAtbB+IUiVeAhqx2OddRN4Kr6iZqR/m7fAiHYZPhkg8HjBnRd34rcyYNfjfz/8s/whT/
TY4nCGJX42KZsnBi7HsidkFmm1LRiIyNJRda2WmRi75h4bSlKiWkQjxSwU0vioxNCt9ss5vFXsmw
wHni2L9uOOS5w3p9QfHd3BlIUqV08XhCRWVtGW4Vprhrswj/EBSCmZ/pk6Qm+GBA7NN3ySVPwATN
nEsbVRxbFZthRA6/ac0ifLulXFQQNAt94uwbqvhr7HXOsSX6RI07vABF6CQ+ZuePfpE9r8wS/q4C
7ne/xpjVZJ7MrngZMVHyD4XUQYJybtEaO2mfQ5uMWE95pX4HWh7HPLKXIYiuQ2jH7bFyOeqVre+6
mUE8+xIMx6gdgo93lQeM6CGQ4LE+pS8uROlyLzYE3Qgs6rEbcAoi6CwGsaTMYou+KsfZ1JIgudNX
pCbGI8z+foqWtn2eMxKG0J2MgMDMAZjTzMZDnD4QHXIeevRzfw8P99Z3aUlb5RSJ0oxiMBjLguag
d+/jBRiQQ02Ic2f3/Q5J6TRp5ndUfVWBTQg4EzF211d0IuRJvugr73TGaVPhvTXNs6rumW3Y4XRb
N15AN5GzX6/Tb+nXfv40o7AnxoqQ9oNYiO0wAFoW++MVnvSvgmbyhV5l+HB6B3k1wf45DnamEM08
wJcNNAdG8iaICCZpxShNL12jXRTxwTNOga7EThBenwxJW3pCSTCNg7JlWP5IihKTf1z+ZK6azlIU
ZDS20WLLDnRo3usdf/kNDKCgDI177M2Txex4grq43fmI9VbQk25hYTklLK8wYC4dSRyqN1DlTKBH
4g1WEaXGnNqjC2o2otIKMVwDx7BfBDViKl6nYrLaWeQvdeSsb1va/fBEAP3xXjsHbMEnespfri4L
aGAfewvLq9sbMQ6FEKT0kslxWfro8/G8f2hzvO5jlOvSa1+b7XNl2zV3UMRBmyGpqaiB5x1hVE2a
HYM/vAkoIxm41aSQ62XnO1DoJUwhKKiJs6SMfkh538dK8pK28JTrQSI/8x4cZmLBK2Ly+vPWQ5Mh
x0GY7KdQxicOmcxH0enZifA8abxrO78YGyB0NivI9psmifX7qL6Df9CiWN8/19HSWQgUSmIxVkdv
WbKrOeIJgwR7xpFV3OsBhKZd0xkEiYA2hwarRE0OYXzRTXnS97Akisxt9g+WBS8mruTj9ufUS+ZF
KmSZSh68GjxjwPH8HqwRM7156dPnqs4gzrLuNnPqncygbKHyELgELed8jJyliHGKqsBRBF64e8sF
O1K8rv2iCD5FKl0p+CuUwHqUiuhosTbhchGzKRnX9DMh8n7cUKxT163lAYKEmwswGWFKuif++nPW
ADawcwHlYGQZy1Uxn0KecCdrxqJpKUpmm+GVyFuT3fzRtb5AoYsk8YMCILM99ltwMDgv3a4CVuym
sq0kgBgQ4JIr5U8jMpvHQm82Ap/uKKHQd8Jsv0y+LhNPTRmDKT0k/sC9HsnXt9M6/Nf4SzUvJdTF
swObRLsrVCNNhvnJUMFyc1sF7VAibgRdeoUR71xEETI1FSFxB51Yrq5jGLnG4cJAvO6ZwP8nDrHD
yY5z99QHNzZdEYgJETUuXHfD9S3E11fyC+yCiNpZpAw/utD7zAB0yZGIpmY5TgZhFmVfr5bnKWO3
euhKzM7Mczt/kYEAdUw5MGu6mH2ocbYlKrPWCbKuoLTTTTfbLIarS95ALSgVE/9AlkVtNggfuTRA
YsZZkFGadYl02X0uq65vctxekd96Uazt3n0YJBbl7eG/rgNABDKgDXza4ATMA5PsJQE+Ctr4L5eY
WRR53foLC4xjixh+fB9204t/rP+TkdHkBWVEw4Xau91SnSWtvt2LxT7LpXyAaQzD5S7XCLqMee6S
B8XN6C98ueALsMYx8x8afYGvn5xbrd0UWlsDziw3YkSIH31oAyr+vMPD1AvgLSzdwZjpS92XXhBz
UepqrKAoNLTgW+COqi7aEGD8kHFcr62cm0aigK4qnYIZZw+cdQaP4i62otWFVYNz+MY0jd4wFood
DazGMnH7WtlUG714bfh/RXf2u+seMBiaA4drY5Wakgjcx+n+Zv2l0cepyn92praATvlZkfM1nZjE
aa9VTsHcAcb6wLe7vqukj4j+BvtQUL8A+Eo43bw/EPYQf0vyai0Ux+5gnSQYYSD0SKH+O3HfWeYC
7cEKsAEuMeQ3U/jq5hfXq7vjh0k+IXqy0rn/pcsXhZzoF1HiIIG5Unf+93FpjbA6RnaFc1khohO9
VIiO3FPNER0LqGUsYI3j75a4+yvPj/BJYSiXO2y6KfRu1VHGNOsersYA82t23y2usIm5h1cz+mYZ
25LRf6bB1MVuLJJRiweNFGCqpMFtGNn88tsGpxx0bp4Sw+kWYw8a2htpLFJN0lT58LYbZB5FQNi0
rnqIvsjTyXzmut3QCvunombpUDbkKlQRpMht5YHY+b1Ig6G3Dy1peuacYRQchkp56uvT/TTFjDHN
QoKr+1noW+0MtqB6x2GiJkOJErbucNv2ORPSaFDHa9nWC1ZmzGSEfXQ9341UiYcLLA6ZTJQNxlH7
l8D/L8WKsgpw4jbEOcdOaDjqG5R6Jgvaqd5j7Jl2Mh6wZe/3YzUVKizTQsjiK15Gmk/KtWKUajiI
HOlvgwnPwFkiCYbNyQx6+XHVaozQ5PCHa9RPHjgd7K9UoFAIZAgrYwJX0+xJn0Fz2jXXrPdUCRh2
GLiuWuJ5SzbjPdPbwCDnzfx05G8s/OVB8KzxjJO7ZbGXoglrF8BDNX5DdUy+ZzXlJcxIHXlZXsQI
nPqlUeThvMCR3Br/CWaYsrv/Q6U2uwYuF3GMm7feEVSer8oqKW6IlGXVZgYhPT7Fd6XsnHeSp7uZ
Vpj3YVyYzbTLbGGEfQaJlDekmVhaalkFIr3bFKqLJ1FrF4maz5cpTygD+qU1dwy0chSdbqqx0gqS
rIWtZy2kI/Tlq7+owN77XAqc7ERJIA5LM8XvgH7y/LjE+eubvEA5P24CjMvMI/7Zo6gAM8IQ/bmZ
SmTkJjlHIcL4zusVMqfDCr+6AGGeKu4+n8E5QM1BqfYUdNTiIrs/UcP61rdti9Wk3FRR09BA/Z5K
+VGAjaogaCByOnyTiYUSxJhbbrCqc//hiPPlj0PPTgsT7mnPPj86RB4movW7pqd0DdVfHWHQoG+c
hxTbSAO0BVDyAPGCUoyduwIBSX6ixkbOMLAKYb0RfY8X/6mRBfKtAM/s1vjMs4qcD+2cC3y6x9bA
0SyYUBQp+1VMFmZv0DeL4XLnkT1ImEnH2vIwnofd8mqkfoG7zmqaqtIy2wk8QkCqNr7AhakmUPTT
eqGt0XARNeidX0jg5/vNufRQsQ4I5BGR8JpOP0DLa85Pt9vcjvSq2HL0BnYgePdOiLOEA59zMbl5
s4Cambh111PLTE9LkyNVDBf+o+ZEV2SOzhFYthJTBXg5optF5LjrI24JFGS31EjIIbgeHhUeKn9T
GellYXQefcPA3QHK7UAQp923lUTrekNj+474Y9VTjg4TPAmgwppMlDFmYwtHZ/omxHnYBTM2j5X2
5H8LDheWFr4ucPiqhuk3uqVZBzJF5TmmHlxPEnXRYqscFo6pkO+dtv6QcJ1XJsC+EIrlTNdVsl19
7BHNllFHif0OHivGoMVGShqlC4XdNLRPv7Ckm1f4FbcXttrclI0BtK9g5+pAv0Kg2WDYdCX7X0sS
FLE2jsZzaDSw30FIYLnaTL8scjYbeikC3iKpyCatF022t3b6sg6YVPzRSj4OvAjh/lIAnTn3i5ov
AjMWXEtV4urzydYpg6ZZdSKdEH7WumYCYnmTuL6wsI/vFR7M777emvBO9HxduFSxQDAxgBtPKQTI
ll4T6GIcdoSMqV/dqPqvjBHnglW0WEIK0fsTwk7Hk6Y81/33z4K/38/yWg2yUwRfBx308zFd303H
xMDrMYYf5LnmtmA0X6IuwGofbR+KzWpTsCM4MdNVy7oKOfLiiP/GYdiDnET4vLEUk5/es9Nq/urz
5pSDxPU/BRrQLRjTBHHq5LMkCTlPgr+AogaZOr/LQU6+7KjFFMxasMQCZR2iIaOH+wxQUVNWD0Uw
tmH5QIYg1Yp2Gx0nCLo04i2KFB3b4rVPGIf2OIyco+i/ThTf/apuAHRnFACLaJiGcZ9MTj24HzBa
4JiOm4+6iSubHaNZ8c5MFHzt9exsNrgSoBsssFntaV9XySUTvbE/AH5m3DrWOj4ZtwDJN4NnGy0k
AdK5cEWDiyrOzBExf8YdSHPK9NWVZnNnoLO89dwUTu6r+zpdLKdRfQPWYn0Lri52eJ42iNedNcAB
M+y5SnByAkizZQeVn7G3jBdoskvnDr70Hc818l6l2eK1U0sU9LXE2U0v9Wy4HqAh6kycB4q98sb5
pQfoBpKgbOr7wXUN7UA39+Dhr9YTuGz2BPH+Yr/QjKILP2ea2lBCx6bslNyQwUNPsgXPgv/TIyvY
poN/gDEd5R4YmWpFh/S6sWmLqjxnUpkIFhkhF2kVrkbmQToFxVEJtIwv8xcCbjFo4GLVOjoKd/q9
8lzbMfLdHpUhazeDSzjXdaWRoKzSCJZOZgkz9N1KKXmQjDl8Mue98c0Gk8JyN8lAZI66U1AD5gBt
N9Y+/nPSZtyHDKiFaCvehWFGW//hKGcrc8ik/krJ9dQhM4ede73tF5BeEDDt28ub+PclDyo4KbEp
Aed3zgSuZkWJ9EsSWgP0wWD3OZA5B38w7ZXFU1G8rN6ZXwyGrj+z0baVzjMk1ztZMjgW9aouOiLc
IXImKB79YLa729v2b2xWSBMYUCpmmes1VgjN1rsfhKu6EWKMduoOblWGKZ8V6epd5VIqVnt9RQNx
FtHGi7gtTrPAlf9WteO1MS+qDA7PyNEAUmbDPjwXkYGbLKIV7+v0QjX0JG9QUZBre1glPqhmLiv1
1yHRb0bfHOlPikuWRsBuyt/eyThKsI+nYCJlCqS8CSRnbmd02ZQtY1vMrLIDgbUVH75/rUfON51H
pKF/HwwtZPpNNqOHCet+2x9Zf5423X6heEuZXx5ZZNfDlEC1Xk0HQMJsJ5ltlRiipjDT0g74DYr0
yJw/kBPQjFUkPA0bBtZphlSOrXGYIYgzd53Qcwz4UL/PE5KdMYyNxx777xj4SuT0TvR3qyXZ1A31
8Ex1Y74QuahZVBbSs7cjkTJWrIBw61+Wg0gfKr03DpaMauX8Zfb7ppgJ0yX29uxeq1XZSFtQ9NDA
4n5o1T9CB2bmYukZUvfu1vTILZh1fg4QUTR4H+DCPAKeapCVqt8tIOJ2z0D2UKkbwIUFVR7a4rMn
kb7QQsRZsuJvg8mjVkwoC6MAdDlNhZMaNfOzGb4KTwTw8ZT4zOPqFEubO5d0r4mSDOzx1u02neWN
auSbFLwq7EkT27GUrmqjOqJOKrqmW60iNeJlob5ePZ0by6Xwuk2qksJXpxn0lDyhSqsrB+qAUuck
L2avQlhtKq3mwpjbWUk/crG4HdEQMjCWwhgMNp5ny/5JWny17XL2Ylj8Bvy2Lr/OqmxUspksHOan
nvK/3KR1H61Tq1G7Fpxxe7foItt+jcq6CcSCvydhp5DPJVp4m5DJriOQ7v+qvv5ecJgdgysB/5Tq
32Cnjj1S1LmzpTjOxV9/Z2CqOUyyGQPvZqFRNDhOBGkaOT2QV3zCG2B6yYTHGyrtTosC3w4cEC86
dOV96hu5NlkAAV1mvyhV6JdbdmlS4OD5R2odLzUDBkN2TUfeb/wnirvNTRu86Enzx+3aeSuDTwdO
V+0KCpXirUOs6DIuSs9619Qmj+kMeD9JURMKIWAUG0P7HGeIoOtTf8NHJbolY6UzfbNW9L7rODrs
lOD+/Kx2kz1RR2RS4uEO0Dc2IsVg+mRxmOMd4CcbmkDoexDhkmxCsA9q0BcfRbs9Dz6abhzc6sgj
zA0nUnntQWqqMmUhzSUd2/fEpy078TSi3MlFvrjXMdjuqqi2H1J9j5jOBYImHb34iXdi8aP2bNRJ
3o9Wy5l8RtEWkvu/pMJAjcUkQMianmEAEmBpesnddyEZdmt8Onpx13FxKBy7WS/Oq62Iuma1dZ0J
V8YRTVuGEiuTg6KmyLjGo7cwge5vrdD1sH8BkJSIIKtnegDOidYkHGGWO1X7du482MGpWJ5YlbWD
7NFJpLDmv4aFbXQvT4tMHnIoYfPaji8Ychp2bM7Y4yo/UtAThX9ODU0RTLijQ6Jb/QcrEnAxGdBe
JaspKOCv+4+VzV1WqUYD0l3hWZvVYXZMDfbYzBXoaEHRfQe5Vz/VkyIMTnTghX03xIZWWGD59CST
HmR+YhByNFfrEcwCurgFXOxhQWBswtoEgAzJU2Cq5yBNfTJvJz1apAjscJfCOKUmpNBYYxNGMFvq
+DsUsdywBrz57ZB2uSihbNdbtreBP1bK1uZpMcTU8MNXOJ25hK2TWN1n9HgsOonQuZOdNHZaKALC
P4wUnKVvk7o513ZH/f0QcyR8zrTD7bM4tCuyALOXKyh6c/6hszqniHLpWXUQcp9RUswN6SMls1NW
5rYsbWabJ4Ba8A83BiVgFlDa8XuYtC6QndzbJBxCN2yKiXfHS91GvjGiCKT/EpJUyH9JwyR9SHw6
DqkOwKMjlSnjxErVRDOmyfRookxFfGUiBh7acKAzkDiMVV5J8dTWVxL9ZGV348qjTAh13OBrtQYz
5SlLDtUizYM+en6HFPh2Li16/HvN0wjlKSc2xrN3keQi0+JM1jzJ7I0nC+JN/0y5OeBCsY6CQPRN
eIc/j9SexKQHSqugiMKiRQzQ0KWM3gloBTREEicDbGfLkj4Ubl4YG+cs0h0Ei/GLL5q05rkfJWf2
XUAoBeK6s4fOHB4kLiDSoKK68oInz9p4DtUu00MDYyLKL2lwMT7bUM0fuXEqyBXkbriFfT8AK6+m
qqUknvSjoZfBMcxKpvlJsBIVIcvMtUWvT07ita3mkSK8UpbtPUUZXERtPWum6aihXDpsXtjEhZVZ
zXBdRRlGJEO/TOnf++Y0sbkc+P+kN8lt0kJagFQ4kPHC/TPbqGdmL/xvo/TLugR3psUGVrSz96JM
yEj24pE6LlBIFcZOcE8g6jMOPfbDtm4IylUqVXd/2z2ftqgojZgj/uaa0/raJAiMBoesT3n9GFUv
r/cc1g/KAbm0aN9zxVqTYhdnzJHK05WNn2GqT8IkcE8/6xeTq6fCk7auChCSCHc2lx5Ln9Dj+PtC
DjKKgMAkYI2FQnPf30Hd+A8iQk/v6awlkTHJignG7cfW6dYKDqxoeC4DHgzuBa7c8yCElh/r98z2
9nlJjkX129egVsjHoWOteuLsKLsPlJ5okMzMxhawsgaaG4oiidJy6N/NGseaEl4M2Z4dLpyKx1iK
PbwSW4KG8p0AwVWML12AuXjYF6O3ijEOVAxXB6wKpY5BGsuxXIUqhPBA6inOiKv/T8pXkkVEp3kS
bxRj4FC/2n6EK4aU1k0F+Euii3saRewY7M4VidiiQU1XC4G/HnDIYAyhqXwus8FqiEfi5P7nwV7M
vV+Mcs71OYeZFhCDx22jUBar9kpCxS64GduwcCBjVZYQ0Hezy//LWx/BSBma+apmmLAlW5ezIbn6
BEL8YwAB5JKW9hnczbC2Nf+5h2ZPynMe5xn2Mg3piOUYVykOmbJCBd1WMYbPOvkXSGgzuEt/vyAd
QEc5eigHGGj3cl/fmmLlpf/Ax3Jx9dwXr5lIAl8K2Fcv9QA5Aoj4nWi423wQ8H0gFsBIJ0j81rcH
p0ytdj3lfgpKwVVNDpHt0KQSer6gVzyfwdSdBpkWHYPEAhuFHG+yV5k1DEyx9FZ6VxwW32K86Ont
nM1SRysM6jChmE2iQ7L+clZxveEPU9eSv5UtziHhG/ueLXO2NNZtgCB823bYDOewjhfYUyAWzqYU
QuzLuHIkGwoscgooaMVi/pU1FEidTYE4AuTbu299Jtt9O6eYw747qUw9hMg9KasKs2lDPZLC5JI9
ku2FBQ2eGpNJQ8oARUVwM33LfCiCD18vYFWW4nYIG34AJUGWK15scTKu93DSJIInmGHpz4w56I5z
2wRPn+Jdf6xOzcXA6Nn9s56dTxhJ+1xoJIUEeg6ZvyToxGRvPeZRBP5JxBwy/GzEDeBZEtQkeWAe
NsGmuyswS1YThMkNjkIk+ZvTt/1R64IgmWOhTAmWsn6KZb7i1nAu6LoBPrlIKaKOxvz7RaxCIvuc
5OaOZMn7/AdnD3ulffXcwsEyTixz+y0CINJndTnj7W16N7m7U55UBXaXxdWdww+/4rThGFAD04oR
KWPSaO6MhBqrnJ7vFWhEhwnSc1iNZeuTe6Mm51xrQ7Hu2Z2FG+wOeBsFdPGpDrlNxUkEStl+ZT04
EPgEQgNP022W1cY2I9GPmh3caUELRpCmJlEMtDw/nCDVYizd/PlxBApSUCGsPNE67IaRySg6p24T
/ieF6s3e+Qd/QnhtGcUTRfYpLEvprMY9adVd2VGU9V9GfhmglWS076Vfyp7jMYQmBenB3SpMeSlF
PpEXRiOLKYa1kHMttM6LPNOnh1mb5Dw14w5pUCUa5UeAlw8khveeLGgrMgI7WaZZKEqgB0vKVfvj
FTo52LdIP7Ds01gRvZ0bvFyTdDVsrhn7H4vUaiAJSYGy6EFB2xoWjk3cylKsYP0Ewam0hSN29Ij/
I2DmHfh60Ifqz0FF6wJsFqJ0AJ+NC15iYCqPhNSBcKLB7GjG896pk+dONB/Q1mwGygo7o68PBPHS
MNWS9umSNlRor9eBlNtBWACyw5UqGLoquAMwUzrNKdTUY/Nn29dom26RO1zfrML+n0yfMkovQOl9
yG+vaaPIvwo/rqe3QbVn+kC4BRomMgNFzHIhxWv3njEPH4SWMQ/V/wfWiVNpKzvxxBDnks9TpKHv
Qy86QDrSCen7k9ZglY2LNo5/hVqtvCAPlWBx5PV5WfwhPE5Xx60dqzIM7trJoUs3B089y4eGM7w9
TWRF9gFUNnxSDEnX3zS6+nI12ypvAKWJV1HEmu4aecMZKynG88Zq0IFgGwe/Xwl8ClveaOn8cniX
zxK8Bnq0UjE9P0ZHjj4KL3YGjpEQBVGF7uwqy2MYNJTNAAFXmzYPsK7HstgL1VMnUAvf56mQP7oy
R/NJ6fnJYikV4JbksoIFTD52fe7n8vJHMjQNzF7E/wc/mn3hC+iK47qTfy4HYzWTj4emT8UGQSpR
6sLcNggk2eFOsLtJ49J5Mf3lgqTwHpPZ2wL8BVDUFtYs7BpWWe+drt/vSZW0etvqYFvFOFNUYXVk
fS5IfYH3mgZA0NcPec6EsqDAPNWMQFRk9LxvaOJcHcTl11UzFOWAIDcB3Q294091UTK9FLtBBsa+
hZn5o/G4bsM2rSc2FcJ4DaJ9CiC7YGRuTreKXJJmDN7wZYdzJ4HB3O5d1uEtgpN1VBZet8QmzRZI
9VjJQSx5g9V+3GbHQJCN9Ot0PSWhRpaB3jZgVOQJTypVibAA6WtDrHCoX9PXt/YtuEoJd8UHiMl1
1ZOMaesqhXUqz7ECqNEgJHsPWBzh4I5JYBiaoMzrjpnx6ddB1uQ+iV8gidnsxm6Fx6YWhFiCDKxC
XyqpHSUjEkut+F6Wn1MGeb/QXxXkWJTgIw4NVdvBp9K1kH3ENpWHoS/m0M9+h841ipcnFtwCTUp4
dI8IT658ipXPxmpIdCrDqFDii/I83jOVn+XPc/NBOuCOjIuIw1ecbq/kLDc6dRIlRpRidtyIuXaf
MSUVlXHA3SqfIW0Xo6VbjEDbhPq3Fh7GHXFzTFIkM+i9dHKYx5OdTPH6iCjI8vDWQfCnHlQyNbLq
iTmWVKqKip7J+5hwAgrfDwkGHVbrETSS5mBzK04ESDvmlqLowTXp0zX2IYm3+ZPRZgn8tdJF8cmT
sdn036v0D1yazLJFPHpQFRq01G4+ZP57O9tFMSBD/n9UciIUnc2H0qBUwJW2i9JeRRTOl8NZ0sFN
l2JZOR9UOhYREpMXycSVuTt8AMskPy9j28eVhRoZOGhxhYmFPPMEvUNzUi72sad00VqR3cEwybIA
DqoD6e5/VfB5g+Ekp90kmteHQXh5bArbqlBU1mfTx0gYCrMuIGOAV3hEwGcA2Tba7LpmhETh46fn
LcqfPjr5feVSq8fAn7eUUsnvgw004iYUuUOoUtdqPjPRUXfiZCiMmfAkdgxPiSLaewBqTiPLyhLz
mZd8TYPv6B/O+JeKSzmDTTMyFC5YtfrGDCdZqPYCrR8eGY2hAnDHij6OupbjiaMYilGdiijVPJof
6asFnzFMWixukEPbLGlgEUkjdVfskcjyuMp0Thzo/nP68wgDAEbtZKFUL6XAoHpuXskaWCPrSLRd
QmjZuE0ET7pZThGIFIxpu2E53AkKDa/RjWWWmf1KgQrtMefV3lwxGFcWc50ljDiy2Unkwl37ZApV
h/sBrj+dQRUsycvmNFsYKVF/BD7ZAimhqnUzwDonMSof08cGG1HARN46MsEphJEWobEw+gfKgcjV
T+iX7A5WYm/ZJEyDMnDN5CTKozRi3NFmJifa9IqzJaC2YEzHVnlLdvrPhiFnffOajoC9N0oZiFyV
NaNhPwoarSn99ho2i8N/FaEFA5KqgE4qoaHIf8AQfwhbcu080fZ6Y9/g4CdIIM+SAVORNduFdxZx
dncpKADtLImbfEq4eInoYRz2zqr+1C3n1P6WWMOaDfzvlOw3BnyBGRvCjqwie+AYd0HpMZ+aT07J
JjY7XeTuXCOG8v2T+SofrKAWeU5YB/nSy9bIMpctPTt2LN6rSj0lo30v/hrmcvAPyx09ORZ3hmLv
GeyY8qt0/2aiqo2xPnAOg+pqZqyMtY4acprCoe8FBanUkrAteQuYLZqVvU4hHjzVrdfWHVkGr4Up
8LPyADnScmi9AjNCHbJwlS/kVM3nM829GgKmLE4OqbcxjQJFKz5UNfJzekkLec5GtP1O84rw4CZn
tdqk+36fAIxsKs7R+tQio6LuhkaBXWXrCMdt0X/quoVnnB8013Ahf8KN5kQEYNH/hHEElv0mVWyW
moZ109GFMIO3M9Sm1p708IConj6mupaaQ9C4VqPR6Yd4DXuhlR+0bKOXhTeCWnncJ7wAJVF31ttV
GrNjx3ElX3w0jlsk9LypLHt7MGOKms1Wkg0S0/aa/6l5lWQKgYPtbq1t0zmkSdBby3HkwI2ljpx/
yb/PieM0Qpspgjv4aCoh1lFu1chcj3XaTMEblW8o7MS3/tuRTM80cB2IPhsxT8+aNsTPnevlicxL
RwAR/sYTpFILdI4D6sIXpu4lxe30WnpAcbSb0oAIDLMdTvboHiReLT6GX++5BHY7M+BLDXl5zMR4
5fzc80SD4o9+LQae7pxgsUxgi5t7ssyUoNmyHziuwvcVGb8PxzOeHlZDTNbV6B5dq6yermghWHUv
MO99Ye42ASg8Q2QGUUvY9qrhXtXEZHoXxbenlmJ8HYdSWxRRlZfhyV/XzNRhe7z219ewS7TRYBfp
S5jKNBFJUlestxV86W+FO2g2VnuSnkF61rHdH9yZv6yrDWCAiEXbV+Bj7uHvxQWyjBIj8HqG3mV0
e9I95WHKYH5oO0RKlCg0GCq/tTV3ge1uzhf3/SC3gikx3GxJlnIT04iqvjPa0fb0BjkoRvQnSv52
CZdcE3xG2U1ehz4ciJvzM+BWaoqSeCWgc61broiQqVnIGN4NOaRHUtHbMSo4swDsxeO0Qmv8DK5N
lAihiJ7xqldKI64GbOMyBh6umiWHsTopToBmTnq7jz4m4DpvN4Xjf24jp4n6skhyjV3ybMmJhon3
NjSVfEEc2NfYkkHB4QFDF+GtcBhwXDMGm32oCdsUBFAbPo7FE3YkZKDzZpOS77TNDKskwd64yJ/f
VlfF3nn9+/p67WB/lCNXYc4dlKj8MY+UCBDrHQG/5tekF5Am+vbsu2ueROReumQUusRxbuWWhT6c
+wzd1odPIW5kCT4nY7nCr9d3lQXG0lYo16eshdyp65Cxwf/6sFYJG7zDvjUrHi+dSWmralJSAcA1
HLuRA6elZIc8mI/3mJkWXrc2m5+QvrV103UbjuHCbNSudUEsf9Ek/STYdtJYqYMXYr/ehZwAtwiO
GhezdQ7/0edjZVJBbFpWPatHqfMF/3W8v3m4ugphmUy5EBgPMWDARDN5dTIpiOEgL69Ash1VBm74
Ii4GvJKkshgQOQxlwYOSq+ZqZ7M6QIOb+DuoUlQ9nmvTxHDZ4gcU6vnayh84RCB4g7PGlRKaTv6s
+4YwPVK1fTRSTZD/qStptyAl3nf6blQ1gbPKCSf0Oq1YUflBRmbM8F9qdkTsXR5EvQfvgtxEqkF8
gqRDgVVQNW+Q7DY4Zzm0ovamWKNinz9u/SBIDVeMaa5IoI5g4H/qPBeDc9lsxgesioO3O+A6bTY3
nPDEA5EnVL7ulrnzZvIBYQg/RSrLrt/ByxG/T+3wTONKJ5TZlOOm/5dZBPbhgyt2TM3vrjnfMCBi
mmQkzHF8gnWBI9v9AJD2l2hG6jnEVvdJdvBN3gj11VSgJWjY+guaP1Qh9GAnOl5JDvJ3aYtXZb6B
h2JSq+h+8k7XEaq6RYaxs/sdg2TK66t18O8zbiDNdvGFY0fLnQiLm9nFPZe8xGudioz8mIaElDtP
6zdFQH7EZhHwipMCKCHTVLsAFju8OEGDx2xfUeAdFvDLqJ374nmY25fZhVl8JWaYmeLAJjWLy3V0
FOqI8cVta9gGjNpB7V/V5PJE3p18dIdNs+gjKlg4gAZT5IRY7TPBcs4WLHDl2NEtjINO+ngOD637
AYIirDIDZyxqz1yzc75RFf0K6fTH+Xxwmm5pXv2DPHkhVUYIqf5q2Gr9PeXZFvIXteOosi0KtkkT
ZwvtUteorXJaLLxYOhq4Ku4LbKXHp+Tf9X8UwSfiIvovUJVxiDJvwgDS6HqkjQafIs4uCHNolpZt
OrIc7RdvS61qJt2l/PaB+spqVGd2gdIcAqTqN7ySlrA71iBagevYLYWZcB4PdgAa+NkB5lLrCZwt
ynw7nLGGWBj/P+hHSTbgpttbmB9vbZX//p8NDjqU9qKnxstS479A2/pbRfWkxRL4nPE/FsZ5lAeF
mP78Dg4VC3nxjVT4F785ZVVmCWpzCM1tiU2Myxb5LbrVinWiOqmKmPHlnpj94Hqu9RQKkaU0AtF1
RJBCTbGAij9hfzb9l+n89HpCUKvUa+K8As5xCsqV6Wnsjo/cMiyXXxjzjIeNb4Nqw1dzI2eN63Ye
6F6Ek9cSpnhV3IpQMMBqg6qsc0expSaB0Lr9czXfYnCUaCr3LpyVpKiMUh09wskS8uy5fc5/0PVD
0WNkguMXdWOi9yZrJfXmaAILT3CNnoI6T/J0GYb/8CScmIjpGsbL4r21TBhbH5qLcuEebv/ttP2l
BODydk+ZBin8P9jiGvHR1uE2zyKGiDIBI228dtBat3YFaVa6WEtDvJS6AyApPD/hEQtAshTcTj43
iinrG6YiGARV+egPXT6edmsA+wSO5o3rJOMR7OKusa28RQPMg4zH79V3GzzNbZKt1tDs8YD1giyA
00uJekgKEtvZD2KGA2i7SFfgPwa9+1yLDx+KKjR28C9Q5QKsmcM9xcfTZD94jXSLl3NadY9W6Q1Q
Jy9v75pWTt+8sW5qhkdzihZfe0cZor7P4AkDOCzqfRYdxeB8bjL5RViYneqcJs9aklXh1gtWDri5
MOs906eRlG0DPZG4Y9BKMyKj0QoYtKn2QR0ebGd7VZ8MVIR8Xeya1q6QPhXljgTK1z9Jxx358kv3
EmSXQI+raHut9VArajfZGBOkMHopsQQIL2uUqXx++73cEXRdD/GAyUAeLdk/V+EB9a4/JMqOCQ54
Plzubuz9JHBPOuPkkBJMxksc2xErRy61Lm03ahza+3JqkboEKGbdeZsv3RBapJpAGQb5W7RhAbcP
GCgoM91bNniDfYvVDik7uWKxU7+KSXLpGuYoSLzA54hG+6HsLf5R1DgnAzH/XroQ26yjumEer19D
ogPS9eGYgYFMpo/PnHXmmplJKMJDccvS4y8Z0CN/PygLfUqBV7Hs54k14ira06XIuW+kyQ3Xa02n
W4cToPGQgXH6LCTUrhuN4qQJM4A4d5n+YsrMe06VIxn72g7zUm2sQX3f81YWUXkrMEcO1cEELvJF
UWvsr77wF9hGjIWfyf11XILqyN1D9K0m7nMWSh+t1fG1vn2kE3CEFCC+blBCayL2To1eZ80NIwO4
HrOzpCfP41dUiXOOHs2I2BL3xkYbWXkplFfYxNF26/prMgU9pse0ws7e2+N7wqomltbzJ2Sl/ocv
2HGgNNdMN1VnX3PNGisR7WIt1l9QkhHljwN/od7iz/KLvBAVrZaSRIlf090yQxRNBAQ8C7jVI6ka
0+kjXAEcCtVT2c/9PDKffVJQb1aDjcevnjk+tBpi2n5UcARYEO9sTCWvgkqOuziz3YrXehBQrWbG
X9tLd26pD+uiR/l/TTqTAbuBKtkdi/lhO2Ox8ZQ1aCL7PQugxiUUZtKdyGEYgga5aykkSYt5J7fj
TMOoO55dTCtX0JJqqcx7wLcW+IUKFYvte/XENSd+ofQXFVybQeKbrKkeLpqsixjnonpqmQC77+LJ
kkomuVkTovNwAhfTwmdJ5alL20gG5zBcM2R0nlIX5s6b8RRxR5NALsRtifp54Vd4UKH6H0J0rXG7
kwA13Cib5D26mmEIKDlzHBy9tjd4viVX5z01ogzmGFbDVvwkrMhGFVzjD1twbzKkr629Ue3MUZht
JnRLDYew8Gfmk6t+sr/4FYnBs8HH58ZJHCERwwcH9syvC2VG+TlZivF7FNzyV0iDCUtS75MOfo+3
opfn7ubAnj0z5ayae5JyBSGcRaGWrRMDASyxo7Vtmk868H64Y+AnfcZgh+8r83ZuKHbGlz/UrOj/
7nWzr4OxYadHMkrXoEDgoK5pVCgnpKhQGjYudFaPXuEi+OMasShlrPsJ25qb7+2KGC9SsXk0cpJn
AH7cFn2ZPpSSrjQ6XXEclAZ6FfyaGDgrkNf2OkeLsnoK9cLXOu4ZpKowzFVVtEVIgmo3xKR8WQjW
yaLp9A+V26Gxh9k5tSAm6KQs4GEPwQfoO642No9QCVZzFEgAsdT0Y8nztfTxKjwOljdKkstxwp6U
u3B5eEbpGGro+ql5/n2dUgpAAu++Me+l255A2hq5AJwbGuvo57xuOUbXx+F00hcAHnTkQiZGxs/L
c4DmhcZIhMf9WnEMihT+8Sx3/nUcKlTEiawNpvxfF26aXtiiWUCPk+P/qt9sOviSfa1aVf90UN/K
wCUiNlTLc2mDrG1xu/GQUx2EZKuh+n8fWnoBnpHf8nQXS9BJqyvz2y529v5Lg1DO4ICPtHnu5pp6
v8yvDc2hgQ1SzpSC9Inn4uLxQv8c4yYZHT90K05vSq1lSIwJyFPrk76z27aevJNv4FO+u3XXFa3U
m+gGuBZsQCnJE3NJ6/fVH/Y08U5AUMTOYciGVDQ8xyaxRSv+XiTTYtXy90cU38uYEhEm/E21HrE2
51HWk6fEgy6dyqiro41djGTIov6k6F+cTynPNKBQhiweVS3RJvt1lyijDDKqL3QwbnWIAUoVUYpL
Dl4PXYhrD006NxOSdzhHHVCXBmRrwTa/cUHeDHPREtFcCD8gdAT1xVYH9Qs0j1avZpgs1pFUs1eL
yJY1LSaX30gpVVIjwjHP5Aoy941ve0MJ7ETEFgdVihPxDtXlCPVaFykiRThlRYSjgMTZGTJgX5gw
3zIcE1SjXvlssa6IRKYQ2qqg6zu6JMKK5rkFhNzxRCv1p/6jo2pJl/c871UeJd+WH7MWG9T4X+Rd
XZKcS9+mTeu7X7Y5eJkuWgKgzVU62qUjuGfUbglNGKO820Vf5N7IaXANfoM5inocyCehFXDJPWnd
DGFo648UmURWe6K7AFQ1zucpU3U4wKKsibnwlwE0GXA8jdPfwrt+1/+UUEegD7KKPQdlOjE3l3wK
GwIqH0TB3PCN43O6q8YXEC3wQQL6f7y2hI5KKgxseLL3OhzdWALoQGsaqOPGSmlm19VbOoY+NH3A
IAWgQXcIBRhojvFLvzzphw2+Md87O1sMKiDBS76/PRp6peBfyVuqTMxHeMxIdf+8K6NLYAnCDrIO
Un60NlTVm8HPDaWZmaoOUVNx+Q854vFDLDH/gZTQzSn4sO+P6spcECd5prHJeutpiQ2tRx9cwqJK
MeVhXJ+NHIkIl+KW9t3liHdebf+HbnD1R9vrxUIXBnjrBL69E2qBtH7PTjt/FLTkmGpcyH55n69O
vyk9xHnONt5d3JVPWTBkJpaIjT9+zrFVbgqkWvqZPt4ygCL7ZaCOoaSTUlpkcEHcs39h5VzNV1nF
quzgZqZX6hRIAv6GkiIZfVgoqNAXcMDR0eK76v+hfJl8zKXJE48z77MPn2Bx3T8U3zHjuS+V/0oz
GwPyFUEpZnBFFYHoHNcS+Yo9ylRaBLJXn/uiR70XsoH+WVVfEW5X/H8PCwGPWajmKnIK6M+bMjcp
e1tOR4acwPovVomOGSTVQd3s6M2wtplmFIhLv5PqfSWyN2uFO8/3CjZep8Cr4XchLRtvx+k/i/9P
r0upgU9+w/UQok0wpqAUOwC8oRKToecPQfKZML34hW+snDpS8faMhvnLrrNu4wnBhIg4f2Lxa0Zt
9oKlBk3ut3jRDXHrnfp0RMYLsse2AqA9YL7Lj4dK9/ESGE0z+98nqLhCenb4o/U0m6iIF1G+f4Ur
2hG37WNUsCJ9S/+CPOI5+U6/oTzbnonb9W7Veab/DoPD2hsJEbaLHOzIfo19RBXIdRHHKd65Y3wk
NcPNJhpwle0EAIjTDXCnsNgsHny5PEL5UcOviTEvYG/huuBNp7r2/MPgiY6eX62IUE72oMuBtei0
g1GVZ9JX8DtAkc9balLf2naf/eOMBW4i5vAQ1yGkZyPxjWiRzr0FeX3Bh/ujRMUCV/kfHMpv7Gry
n3FI1e/3eB+8L1fHJDkOfkv0TlcyM3TLUQqqhmBoytS8H5APzgeLIdI8IjmgWhQuFln3vrXsd6u7
G4YvOrxEhYDAjd3T5YB9uXLBgj3tkBemDD1ZWRnoG8vEGh7F36OJ7osFzSI7GAqQLlSI9naq/Eid
ONwwjheuHrSTG+EofbbDbD42b6msBVMVt3B0qG6subgA2sVILZY7zSidpvsdjJoiu9nYtdCKB5Vo
caY7hGmFObAbw+vplEh4RIsRc4dNN2e/0s8+fGnVayxkWsUhVwwyWZsjFTd//+vAIasfZLOraMaA
hTAd71Dy6BBJLMhk+Xjj268qAVKnM0Nx2+14Op9uIlFVXOWPAlH8EhAE5KrH20n/qfBK7Kdnj2L3
ffpw0VlAmzblggjCHHpjlOb4HzB2Z9oGdHYMb998JZa69UgSKFXzpL/6bbvpjOLTYjfTLjgzLbXu
QO0FPDP4+8FQbIAaLPNZqnThymWuDbjpKnzWU0GoiSygB0coYRVR5FLWl5M2BJXe4+vQYSMiv+Zs
iPlPMLektA50qh7JiXzPIHYEKGTq5hp9NierKbY0ebNtZpBLwupjgrSkiM9ylFj0WLfn5CE+4FYd
yajZ1UbnkZe3qNPMtogxTn1Jenx/C0Z3SIiTkpV8pPiB6DyYfAJh2ehIP+eqVBiAeMIFA84/dNzh
/zpjz437p0SBUdaHeBbPvCC8fz80Q1bpacmx0h7uHEsgU+f5NDKQctWXwdpLF6P/trMzPQclpm1t
v3eBJ3giiVYRyaPlUuV6g6qUgdONwMPkkNHaKXlZ7ALnD8AjQsGBwCCX4xClXaN8SvRBQeNA4s1N
yWykQoh1EcRaOoWEbPMrzzVqzDY4LbYQH550u8GkmbWfupoEq8xRbF8j0pQE3giBl3pkj/XuPAGE
SEwNFvbS6l/nQTIRTKaFtzUOC/hBYj2EvYnhtROydRV9Q1UYUWtALb2YV4l9DmTtmRN4HtYvW0VB
2Mf6e4E9BccLZPqH1tfoptklc/EZfVpxG7VM90TN9pk9fWcr6h7KiibhFHgFy1hnfPnWmyjDZJi9
5Trap/sQ5YoibQXcGV4aHgbuVuSLYWn+HX/1hDPGpu+G6VCCFjZ9calTIIG+G62Dc+Lyk3ar5llm
JMM6kVmAQX+O/LJtx+fTJXT4lAQcV+K4zoEdZ/7swUzfGwC0e2ulE5mxhSQLum3tR+f/Cv4s5Wdm
VZd3Lsxim7a+rn36gh3jtDmHXdrf0iGLi8al6K3ejtrifSaHLAgHJsKevXj/VTaw66+OsiVz0hzW
4UDzzlSyJY02mNIb74M7sRmWfIq3m3bXrQK3+A/de9WIdHJjzB9CyFGGM4kXiWJyoeqVKkOZMYOV
aqsDRMNgHpCO4YO+3Gm2Rb7g6zZZOE/EhZloxvqpk8pNNvEMw+3FVCK/Gt9xAVzYRMQF52bhpgAj
EGLfAeDQqGu5+3wn/tPkXKP7nRBMsP7klWcjiLYQAkSFlEcTiTO3MJ2ytZtPqhrIkOONYM7jK/oA
fgWJ2YkJn3Ad0jeKxrhEY0rS4KURiPbnVjACRV0/lGcDD2q1MXG8U3Vu6GDxgITtzPOfcNSZp2pz
0vc/X9wsiY1mYuCup7HCpitt/uHQelWcOvu2KlEqyQ0lWB91DZPkLhTiifbyP4kOu5VmnHvQLtPe
duXlgr+CiFQkcwQLcjjosParRa5r3WNcMTtjUsqnmFwyecs4pDVBnct4C3qAVGVWEyR/RVDtCfHi
07GH1nmGzcH3tvWeAqmAgDYIXHqsE//OADS6NfEK7V9RW04DrYGuf+rz/JxeAX86GjlmwDAEsGGL
rdLInRm1fIluVB/vl2XwfU7GMEQ6ur2ZD9GdmOC3v1/lrmovFSsCgcQ8EBZVhFpFW/3PvycDcQ7l
L7giC8QkSHP+WUvOUywnbGUMCPgACtHjghZxHaxD/Qg2sCVvyq7oIcq1ZbPZZCxcz4KWPsbOOPEr
lWQkiwY6HSsGlD+cXIto//TpHp+sBBa5wgkNHULFAITOxjr5lsBCUDadEwiiqRRpRdaBDnot0WBf
HZc06S7yvkCgkMYucbxBVPn1WL+V5N1RUiKiv1LQWjS5mximoeYIUbHkFjVAkmIuqEYuHMEabspb
Xx/QXP7OPxoIr+CkpktmaP7vVn3fRobkG9nY/HV0Ue25bLHyj2xNCzWmyAYYydp37P18AEzC41RN
FmK3c4a/2Kg0lbX1l4cCuy4Gwp9rs9R0t6bqQ8leGfGQcUJNiM7wFzxP9Q8uXkwDjWJ00qTTx29F
19WNX1Vkn9f9iIHE88/b4T9V5Izl+9BDjt1eeNzoj71GQVAU6TX/TJS4YreNc8LZ1WNaWEDlT2kR
JmrVyshfgTAoMCv4xisgUpJbvuQNpINZC0j+I4yymIHaX7OlNl6GKD9zH7KZ8txP/y6Yo6QBXU5A
wMizSf5u4yP5/Y4mHrDs4oDABRrwY58K56UhYlbIs0QxQkAnWz4yhCxBdhteIAwLvfLtac04U/XE
Ck+OxNl3Phadx9DUmflKAccnwqo6Pi7CXLgcxivbzF/HdGI3S7cEydxA9GFJsF7xaCWJJJmifqxN
gJdqtxB6/uwotLeek4xue9PZrCikmSsEAenwbAJho+oVN8EjXgls5ZEgRk49CqrtGRKv3oerDhtH
Gv3WTgWkLwngRvKeP/kshvClzvI6znYKOvqC5TCzKkY9g19Zz+rTLr7gjwVtRxAt0bkvVn4NAUGE
GeeE323lEuwN4HRXnf0/CPWUHgJyxv5m0kVIG+X9MU6Q1qvFCpdTJnveh6qzgANeLl1iYaUi9GNt
iQDhyyRBPtwihU798DxP+yyajURSzBcdJwKVnl1dku2tju/aa6+j09pT89eyLMBo8uWft8aO0+q9
hM9iaawcGkfTh88w9RcdozuVbKP3C2Ms3D8GJjuvSqPUYoG0fsjFRrFawcPwnPuEGdAUmcFQgxuZ
mBBEzu4aYiH5Tf+a4mLZj/hmIDQE0PetFPmA5wGZ+v+jLxFdMoSGyyMYTBf9MuFopzYUWXrJ9Agq
8+uxJw7UCEsvcX0ii0WqjwU8Be2vk72+OCL5IDvC6Hpplv22IDe3F5WONC7afdHF1+8yHP1GX9yq
sM4sjQneLgymwHnvBW7YjNdLwlo/YPnsErWwDjeDZ0JFNYb4uAjbpDjhlnE5y17BL6nbRVyVny/g
0EQ9Nv32e5wL+wRXb24DQtWXeqdNGYuG8O4tqjo6bciibyCUF5DIVaFsphAoqa0byO0H5DXuKsm+
XBwgQ/+CS/FmREPIZ8qPxn22tWPBdX2GPjjceHme/PlWQZlsZsmVpCx9vPcG7T7tWoYu4JmY/Vzx
Oci58JbQrbRBgcTK5O6Xym22avuPpWg8Zox9w+Vhe0ArFHzb05D7ISNZg+mb/CpAWctbrpYO8Hng
xdx/NzHh8g4ajBzmuXhpYJF1+WV0d8FpJZIO+4OxN7LD1Z1jhf/DLwqhjmPNiBcp8kYoGBge5M6t
pAMIY9+T8F7kQKo+X/KUh/Hr/3iyDrc2rjHLMvFeFN6nNspgtHruVKZFBHNinoGFmWX8MEnukd+V
VajGfN2zZm9YjkuVfwo2NjUAd59fa/zjSnG+oG6wwnfVUPu7CKyU6j+nvIvafZDkTMWTv1dbqqWk
l/xgi/MGr/1/vF3sYvNqU0O9JcMQRGK98anYMWGktEOYtaE2CTJRYKqhHwfffUVCqnW4/Bd3J/g3
rqdkfSMTmSt40Htv7OXhasF6uO2elMxAEEGUFvLngopSOqHV+040FRBnRX2gG/ryoRnrVm4ZXwaO
Tw7oJgvrI69a6nVAJlgFuUbcJ9rdw/NxAEoJejtsd5A79YBaiWG1PzMY91SBl8ux789+R4N3pe7l
8n4w/CTxk5v4Ubpm9JdZy3vN8aLI9p9xBZeN5Q6nLhXcGd+N1h6w4lWYWp6PszxALZiqXYITPlX6
9w17dUrjOo0JrV4en3QCW05A0EerFWYrzsRVPUdT0hujAmBotpRR2ECp+cwLaJZpGLZseHDGUtsN
10tuJ1wtnvpxHPreKVtAnsnHEN+BpeRF5/LN2X2z+QiZ7sM3LAHnpo6TZn3Os2Wohg4JMJNmQzzU
ox9OHaYttPqrD06jKy7W2G7AvuWv6cGFIpj9SHj9+a4B7EotkWhzU20p2lwHF1W1KuM8UuxZrhOT
F08sdM7K6LgOXzYeZ49TpaFlvSPPOdqyy+BzLRgfBdHrAsxenu8WOooDtsMTX1j/ouRYSw9k1VAJ
oAgNuYOvbp0ZMKtHMSXvAqc7E1eXgK6aiubbWYHAplBQV+KQdnnQpSZLGmgAvCKzXrOFDP1WB5R0
3i5wV0Dsg5B/zJ6EQUczSEf2ewdPkGpsrUMDKxtlpSFo8rJBeehlgl5rxfTAyTdLxmVfvccRfU4J
zbU8sPDfmjrW9gYT7aDoOrFGSY1iQJf1rJrqmdPNNYec3aFGiTND99TyeXEjcFoXcp50U5q7YFzM
zeI9zZg/ewtYNsW2w1O/z0VykHYVBh9ng0UNJw0mL8W/MTwjzTWUOFgiBQaX6qlN9zhVH8QKA38E
ftA+6/DPHklO9HCZQyeWh8dksXxZIYki79DQ80z/Xj258Y7dAjGpUOBVXQj3Twxum0h0k8CK1AU0
8ruh/eSF/vlQqaavsRmLBarb2RIBtKjTO7QbBqOKbIgXjmj6rlw5jopoM98kavBVYbQ+03Mp3Kjx
6FizktibIC5sGrkGkDC+fTwkY81M2WpspEC5O62xfInn1sh+atgeQUgzqy6iLsI+B8MkxXY75TZq
r5FAR7x9gjeWY9JzwuYDP5EbN2wHQ5w5o04QOTQkdwaRoiVv4fJK2CNRPk4NUvS1aAv0ZNHfo7hE
VZeMorhUodYW5Tp1keCqiidUqDMxzhxxPyPfb1tCmLNtpJCcz9y9Z4QQP/4NeoH0YbNHHgJ7YF9U
d6uPMe5hi/3NzbWuuS4gM1GZvAfMzPOlAOiZPe+6zra2Gl+CHNR6RYzGn4SIXcQ43hoRsQGSiBl/
EHKqNDg0JKWLaL2b5fZw3fDJHyAVXLQbHxD4uHHymDnZp3Vn5QFwZ762dsR9BDI1sEztaI+IH7DH
C15MJy4/drSCWGMwmkcfaN7BJf1SBmSBfLzcgg2U2AuQar/MLJ2FNhwb6KDg+no6QDu7iAEAxbP2
8analAv88rWLGqfSvpc8axVcEuYNXMuLcvqhWXo4Sk4LKdKtqWzdzQaXHiZRLixOUTA9KIQMyiWA
I9gNvtmU6tlRs0FGxsd4K6xIAdDEF/IdPzt+gCHq+KbqP7YOSk1BmykJQDXO8kU6/IhyCTlUBPHJ
+M2W1jUq4mArggD7+kTxtVro534QKov+U8Wm55FVu88mGhpAx6KdII07FntzPZ3MzU5KmybvXA++
9SOQeemCwOXfI6N5dCYupbUnONruLTKA+WxAgiHx1yURsSEfoTHMA5VNHx5zLdpNlz9E9IijsN3W
/Cnswt7Eu+oPt5Mmi7SPNENQZYk0kZHP/X/4DmOQtUjBxXxUmvByBpPsVt6HL6dT5NWGwCS0V2nw
84I5cfeK+vCiLAHdAFYb2ocZz+7ws9BdDsZFKs36opwW8IsZkarptzh3FgvgyAdX/n0vaqmQUzp8
btpSYXSMIOYd6f5Xrao3komPrx8JU61Rungq1xHpnAW/t2tZLWBexjXUHC6FfZWXrxV92M87RMh3
UN9YHKHttnxwa52lhm20cOSpDmwWgGvpg3a2wUcOqK1O8DJStWsx7RN4IqpgZlVixThJxu1gmeD8
fmayAJy4GyguvuwG5Acsgb95+xvZX4PRPHMhM+mt9bB2BTBXG3vUsqbYaYJHBwbQc9HgY/g0TQ9/
zq7ibxi55doPRrjjnKrApiHu8beqW2mAXmSxiFxjOVTElWbKcT4MKW+hPZZ3dB+kO8gk93cs9NZ2
KSVej0iKcRGxJ/u6C0ZsLHX8/MmBjn7MzVBOCHPyS/yxLi0D6AzRrvo3/UG9VXhTR31aBJCT41Bo
QZ1ItJL2X/WQzXCFmMP+jGvvmEd+9ExhddbE1Fl4p61XIIUpLF9kkSyWHFIuT7oOwKfmsJFFKIzP
VfvZO6anInDrqKpufXx5vWWcKHXz+UyQ2qF0DO90HkifhNWUfi41Ar9xWuoco7MTi1TnUUqglw9B
dm42D6d9IXMxkXnl6R8uRI8OhD7t/YCcbYBeBzNwUB89muLqvwUqHMpuyj8GN94vJMTFk7UGdznB
ZD4cDGQvAop0AI7TqKUs2yODHMA5As5esA7nHbcdwbjSXJZO0lyqnPpy7TsmOtX29RWB33MW5lzj
BJeZEJxjrBjPHtyTPXci1k6N6x0aWEM4lkVEVrF4IoqawqxqzPs1aXAAXCEJnuYqhhuvlTrySqP9
Qbv5xbpLlYue6LMMWdzDpgWJuUj1qNkdWtcKK9WdIPHjOtDvIswyv2TZ9WU4TOP5PTxEcCwXSJz8
B7PDdnP+vodWfutIU9B/rUjL802fyN6omA/AUByFCrFjydv+2GBS5I0+a/6fB1QB4soKVMEEhpE/
FA9fNjXHx/amefvRwyt0uvivQJYP3go229AvD0DpYTD9j2hldjW4+MS86E1RaCl+/RLiG7D5wvoH
6589gmMOnI0GwPTWjY3cKgyh6jbhiHdhK7UAF5gQbjBbHyVBCmxlIp2fUOxPLMB2Y+02KDEyHvuP
XBP+rd0T0cmnNdWg6DmNiTFUxo6/9VThCxXeLKBpIlLYImE4YMf5sM8Yt21jiDKdbgX/wfWPKnid
bgGPWU/NUPAWiY0xF+8dleZcEDlbcwAIeAdJmyF0GMqlvu8Nw+CCcUfQttp0uSLmHzf6mLLqKScM
YTEqHpBBRRNreI+zLwBCdf8OlRcf3v+48dr9q8hCDUtW/uxV+HPIl7bdAzn3amP96yKj8pcXYRic
EEF8a2GSxefasIV/ak2/bwvXdg0Ern5INX7k+bm1rP2HoJ7WhaYg1uTBsktlwqVhk+zjGBtqCEvX
TOU5lFde8BG45s5I4u2FWtxv1AlgBHczEohktEhfnMfewt/WDtVVkZlL7uDoOTWZRBk7JXow5ETR
89kdqsQxbIeycAZ22Qp4XyIhziyUwyKa3eF9QDDBnmbd/AF/3TDkIZPF3wJ/Dgas5m7NhBuZ+Wcw
vl9EXpljKBFq0AF7Lt8bwU0NS0bWMcBBc1l1vg7n2Hqeq7QAgwhuD4yqZA87nAxA/iWr0Y/yVWtn
plSbukCytZq7tnyy6sT3HgWoD7cFczvJI/+DA88Xc3BL0eMB3gZXTMrUidQoXe3jAKZraHNJvYJo
4SC1z0nlNdF7ekTZozZjn61WDV7Hbd3i4276Ye5TVwJSjIJ0uwFYainWdKR+P45ZuGdIMPSlrjFA
lJtSy2k1JqjHYjfV3TcJVNdTXf44TYOm2dqED2bc8wwSnwyB0WSm/s5e1qUfYq+Vm4apPboze1x9
vEAg33KvrBXgV4ZA2ZaOL5GwJS0On9wU2qij8OnZGhvFlbWbvKeDPeOtI7VCHNPBZKTvsg4DdRVE
KNJUXWd0TX8t7B3g6IIdf7Ybr85r/GJju9k8dVkVltLIh7FnqjPZvFIuCuicV7esnBtIgBVdl0Gn
4/AWYlSKiBCEEuk2Pb73pbRDYIfITFvAmlfFvdf6rIO7T/PX4DhYBfXekZ9t277tLdCGM74xe/1E
j86EvbemZ2yDECQ87hkKvXFAKbwNf6ugriBZwSawzh5jDQIkzwUjJvLrhKUFyZwG8VAxq0A8coen
JoqHaRBAaRtCa9nnFv8bVuLAUMAZruh48kTVdfwxuObYexYcuS2P3YMt9D6Mof8TDUt47i6Lp1T4
9lr5LYXr697UvweCB8Nag6iB438KEJZ4Gv7asLbId19gLzp0VQ3IM06KVE/nmXxuxyQjPjK37H3E
HmtdOUiO0IN+SsW9sse/eEwevXS8deAaoRyNbOny2Dczs5CN+t4lpYWQne7j57IgUh5AZfUBPwZp
THBPwVuqA9y9ItQ+g+gQMqaKu4gtt8H0MlgCBID6WNCAeEfj6ZSHuh4n6SEegnb7ED/VafFh7eIe
p3sXFpitWYPkNqge9dPUGQEmNpX7yFK/7TmiLKWChg5amKPuXeNOBLNUnF8OpT8PgQf6LqNt/YNo
uLTjKOmNN/9+3WFn9r5dMtxGLWhqmtvsWENhVO4hLpr9BJLA3Vq4sOKpc4yVbrVW66RHDbDSC/82
sPP1QJUveHHtwOC1MDAsuds0Xk3WkhwmX8AG6drKi4r3yDdB8d7RETvHNlTNSFNRHHUuslwC2pJF
8Gd3cuGR8RH4bvD+iRuQxwDC8kVrxtwdoAiT9KnnCv1XYw0wAOMbSiNRsbNC/IDkDyURre/4RgFs
BnNMXon1nJ/vQBqLzPKgC652ZQlk4s9bp9AqtPI23hyvVgpm5qHUc7eahVMIp2zG2mm4gf6Huh6Z
emVqwfxKRRrSlG4cKMJZoJTcIMCKaiq78MuuJXWDZi+jdLeSF4lumqaK3K3ZGw9zyNMdE9rJU5Y/
+1kQBikBw5+h6rj0cXIcw00OiberJQmWbRjkgKOKwAD3NtsTR6cU572nlZs85RB7ZkRpFmWQw0UQ
oo068nmaZhLGhDMdF/B/sQO4QN+nie3SXfB1y7JXH8IOVK+CZEmnd3u7N2u6IEJb+mIAHeU2HSxl
Qk8mqeWJ2OMburvf2pCL/IoCxD05xhYiwQmUHldkzPnKMw2sa803ivEEL/zilJDIZYnoXkpE9e+5
TS5pSdlt45RP87Q7ntTYEwNGpjJc35XQGba/EVq11pD/CqOobWHyR2IVzFqLjRx1O5gxQ7VlY+cT
YL4Yc2jsLNPvHOzHaUTROXD3KgnUO8luzJjZmRnxGQR0jVndOx3D5Cgb66zg/t34sLaGLcqq0AXM
u4KR3aovZx9E+ZeqDtNRe2f/VDlB94ZW91dcOfjw3KWGAg0yHpBgT16kP/4+D72AtNT/kE6TgV8Q
8ZzpYdx/DKAp7gauENe1Nc9vouRPEu1jQTKszb8ib8u6cuVt9CLfEORbVEJVfVqTmRq3YNLfehm7
zRAtDpMap38nRfr3F2Y9nTHbzqOi2b9cm8GlP0CPVfX+UVtCuBGqhsMHvVFZ+VP65NKPl40VimZZ
iJIyhmRFpIcThHzxwDM7HI1yoEEHhFAT31iVOHKzZmMb2wLpSgT48oXSsCktyUo/yDWM8m9lg0zl
KvKDabg8XkuowoYjCq5ooGc1vpf0diTla51HCL+ZaUQmCXZd8jEKy+Mpc3Tg/200yimSmSNq2jsc
Ups0bZVrZD+ymxSNN6ikNu8/xxZgGtCTLJ8T/DIebOvOHaj2GkmiNuklpjvmPeLniNZpE0ZkcE8V
ai8M1izSNSjZkb8URjZs5smJ3XIlGM7QQsIdlFovN81y+wVO28gmxSaZPhHrVL+lj7xrwhW6qdWh
HPgOeH6XLVoXDut8gpEGZlJnMJj5OmlLUUnVAbOnKVcZu/NkeP09rlTb6HlDEe0H3rM2lse8iUj1
Aq2PVOYOw2pkvqOCvlycIOp3H5ZJ/dgW077Yy1jCG2Ki/1Bapzp9gQWNccvHOk/CpxjTNwIALbZR
v2XkQpwYFxpgjxUbhkAuOW+MBVuTUnFGW8I6odCD/caUhkwfJ8kUUTiKjyl/BzT8U9kZMUjd75m+
O/PWqZCkczAOPLZx+XXdIiUWVpcqYYlhAd5CdssT5GtFPNbL5DzhbwpNWmJKgEuh4RF9hw2pD1Db
s0d8L2oGVyLWFOlaC7XbZKa4/lrAd03XDt+aDOH8wJdP4/bsmOA1QEGC4+LaPGzLydjPZT8Pu1Bk
TfEY5EWQFGoUgDxCcspTYawDw7y6IGnc+NAImSs+JxVvpYIXnjA1gimYJiBstuTpXvFFhZ4AiZo+
fUBHo3j/5gI3uK/YP7Wp06q0YRCZE2hcLwyf9fTbGVtyOZafdfq9me4+jsFujsZ1H6S1I+IprDST
G4lWhH0Xr67jHAACh0Of4B+R+cPXNaO+HmqC4y7fp7u/pJMcs6KEDOs0zYgthg39NcGFZmXkh6H9
RWqyKFsrdBwgguEAxb9k2FiWtPKQmG+jrmws23swbHLftsAvNX6mgVx0hi1Y7rxUaYDR0yjCxgEn
njsxiAx5VE2GgEiFsOJ4eQ/LEt8PDxZlVsLT0kogXbE0KbzjwRYWZohvdwLxmrW8U4XtHXGPuJnk
dOyzNQoTulG6X9tRB0/m4AaCRwQBQCV5/o8kA7EtfO1nEA5ATS6B+gCDw72+NG5PPFQUCL4YPnBd
SkdL0rTKy+FIVYhM1VhgI0X15f6YzUmucZTvxe5wfAfI+fPodJQyWItFxpu399gXBRcL9WeexlcS
PxdsRs+xvFQA0EqwLnzp2abLcQd+htI8Sx8STgKlfadnTAC4wiOArQFJm71xDEm7wRvKegodzu2T
3YEqRA37QSLpkdd/C+oa5e5LqYsXFhS5Ht4yHM2tC2ek8we5Xo7kG7whxyWASXcKVrp+ZLrFLSFt
7u8EZTW/IDHoM6vcZuPR6UgfYDnXw33gYRXE8JC9OoCYekIPQS/xzYUV6yZbjDZSlXBBVzSMaBO8
pti8C/fnE1KWsHoNhcUwJqNsMbr2f8MW94DDptE4Fd+rPTKQYqZp8Hb5P8GGvIfY0XxNVslSYSju
8PlvdTqPZjdchsMbIu2Tb7RKmOWCby4UCFnz+UHJB56XzlF5pWBXR7NOIZTL96GkeLiBnfmCJ1Df
izaQrkwEHCvGH/Wd3x9g+2+TErQiW3ENGWL+GjJzDN9d5XjvUD53VEE/6BdGhbK3BpNIHsZWJ76R
rchZSRV8616N2nvK5KSkVHGjBT3aL4OS/68bHUs1IgXDJua9Ee02//jvGTmwFuFVzumfT1ZRMXj7
FebwEIj/zM4i3N3GXFjFVd/k4MdqG4DNVnSRIXRCXFKpl8XJLlHAvuUPamPHJM4HOJGY3ir1aqEQ
K00VWuz+BfM+n0dfT/VRjs8cbaro8oWk+SSXJDxNruBDyOFSvgWg37ZKiAM8PrQh01NNg+buz7fj
Z7UCjkxjQ/lmcvTUbHJ3juCHKb7T7MNYB63SPWNFUiO0dm4gFq15eRpLx2pOdtp7mLN4mcyEzsoL
6BuBIQ8CRNbxLDx4gdxqRHmRFj4ef+83KGm/s+onNWQqmogQ9wngOQZbnlqggO1QUQBBqGG5B0on
G4JpbUwE3ROzfMoAUOTb4OvmvcmHMUFe6kkL878zORAF0teBDPyb2wiHUU1B7USPmu0H5SpACkzP
UqYn1n20cYNxYmb9bOFpRMa59MNDHXg1BSSaxfZN5F8KHbvjrC3X2w3IeRhFkeqTY2vc50MVRG11
IYi6n2ZihiN9psRiEMprTCr20vgS8+R0Kc9lVFz/afcuLv1nEqttBbvaWcFnTs34CZelEcga5L8c
zj2nx39ioTFIXHxVtPMuRU4hdVeIUQbzw/8nchrAaOWMD2ujxoRgCyGh6QCs0/xRmZqjTjTjntz2
+htBF7WbWBqAFq8B7z9kdhpQoW0MBjfEcHQyk+kPepuMn+AVbzfubO7xhB3esHTrIFIa3TG1mxdZ
1e/TBxU5MhTLLVOmTdSMnXgg3TgxFtCR2kX5Mi03+Zq67c7VqQ8XJRYcbEbAcWH+qOGsJl9R8Ndx
9eJxeRyPucAvYW6Uhy6fFA+mAsuf6QyKg+458WRGpmEx1+66W7kTsgsqViLpYJFJWeSKRC6K4Zkg
uOJ8kKlQgvZTT5AYCyAtOsVfwMdclOCsFDk9Oaqhwuqh2XV7fgmhDNmknl7struLBenN1dxRTPX4
piDzN92rFDJyKAHzds+PrgZZ8fADQw+zfsYu+s/dpjii1wiQ9cPGmojsZSP+CZ7VW8kKKg+E854F
7OUXxSOUMTzAIhw5Xjk42PF3Rz8RjKSfI9wVt3ge2QNgP1wPFmiFYtIt6xQCoi7KM6glZ6IjcHIq
IGRVgYTJEMtDOkoZ7+xkJ2s3D/H+KdNRd9kIrdrrCiSicYb11WQUNSqfziTuibTXNxnjS2Sct2AX
VzOm80Nl8omvVXzZk/TTXg+vjrQlqQGgmluFV4I4tOSEibxgxbEiUC7BhpawGTw6+5XZqMYoDAF7
ftHmD+bmFPLPPLIUTI0yx9Uafzbn7cKX/ptsoN+HmQ2h8MjTZPWdCVfeOFSbGJAF9EaLQIX4O0C1
qBMzek012zHvjzVYHLtxnbKmVgGR0z3WXI7aYTfky5Uj/YKCNzzEKxE1oMrfWKwSWDlrMYPr/aWY
SNa0Cd54qnz5o3Zl5SPnTJa1RFCnHLs3HicZhppQNu+id14EoTFUZpc1/j3dKvAzbHpa9nhtcuQ/
14n2+h+3BHMRqIhZTjm4sCfOMcwb7rnHgK9jcqRzPc4dAcuWg5Z0BlmcRf4OblEoFnyFKWYL1ZgT
rk9x66EtlsE0LTbTo2xxYQZqGuyTAfHqFPH/nzdIqh37wfOyYsdCqxpSjCLM5MOm3zZuEauVWNnh
eQFUO0WSNhJ4NqmH2anwdImfRWLAYqA4LBgF49/Yk+wIqNj9aIiYA1300Zi4Jc9LXFSPxpQkNjoF
1k4dsa3ngdlyimU61ln6vAu/KRYOsWmxl0QAL/3XjixZfldg8/BifpMI6+yGqSFYNIfcYWj5DKgV
+z6kECcQWRSBviTR1jCMofYWo1OBoTpYNOUzpPXD+URFU5LjH0w9crIVW3KDhFMICcVmv5abNnHS
xw+TUeaTHHUuQ0VtPynnGqBn40KdwCBqBZoXsaM6+hUVm6c4SHLnn+IBCyjiZS0GPpbUq6No8K/A
mvOVf6O/hyMOBv0+wDEkT86y/7kbVqeSC2G9XXf86IQMQ5908skT7SERdaJKm7W3cFoWv05JgK6O
M8rFzPNLmAagBj5OUd2SY4rpzqgqLbZYnQacAQKcn3xyUwZxBgAcIoR1UCnozeo/rvIq3t6wHmJt
vxIbQ8+yIubE15bzi/nsW55X2KmDBXy/7v8fMk9qi3AerUwrGBP6u88WhZEGm16mJwBIl2+ORXBo
kKwMKqAFro/IPVZ26MbZaHUJumP8VgEesUx0VpFP06VWZWzxMqQx4hcvV9HnlIOX6KC33NeY8slg
ZuVK4byEeoQ/5QczIFUO1EJZKmbNqLbHzlqbEHaBz7FJDP4Ld02Zkw2C9fs1HagQ/4lKwlTq5cBm
oMc0FJfo80PsNxSoaifDAuX92/rwoW0oko2cr+rhhdIW/BP8fL/7sLghgnVgRSYWmLIc9SvyRP2Z
iJ4wxVUZqN9FGUwNY0r2E+oJbb7GmmymmXjz2e4YZsIfWOO4dcTcB93jUUwHlTIcp7sLk9wKB8dU
qDulGmAJ/Ilffs61n2PMbCbpGbdfJocQCafgHuls26VZKAJRi9IX71tHXgnWr+MzSTSU6eWaYoG0
F8MbIZ/sPSFSGzinj+CTRMzHZ+TIN+XL/S9FyYex3Fo8pypeA2ZTmQ8KzziEfOTImophby+6fOPM
YeImi0rIg8quhyp2J9Ktx/gFpG5/cCuSg4dfpaVV6J3T5zwOM6aULAueWc1/IzhiJLsCAbkI3tHm
SylmRNJMyQvdLVWTL+xRZCtLFOxAXLG9bXI0n6FDpmGAuxQZlheN8XZ8TqzV54/KXTRx0MJarbuh
F7bNgmPXdQcs3vYQoqe+QOZQBoXJKbgvZJEr0611ss7RbFG+rtb74BcfZHysw3T2H5mh/iBXF/H1
GLflDGKX8VsrDpTCGNzDJ4FwQm+Mh9iWn7Gh1p+DZb8pJYSL7eKyzhHg3FThvFo7dCSeeBYuSuVV
5v2h4JRCP6aYIR+QDDvCdypHAuoWcBM/etzihunaD1yUQRFFAbkPCoF5BnwfEo/374OgGE6Mckbf
DvjAwhdoNJEV9YOLydBlgEnMZxPz3MR6kBOabL6ywgtRTlwslChO3o7KWAaRpFT1VuUsQInr9/W+
+q35nxXLj7Aj5jkq0/jYP1Lt71zmFzXNWlZUnnsRasZg+o9yba6oYzYy3AKOmrlYcoA1O6kQ+492
l2Intab6nF3eO2wMOzYGWeRYfvoM3k3iT2UAlwROri9/5AZxiZKBlZxpi6NNQAqivFxab+H3jBkv
xlwCL2Bz8v7EKbK6+rPSPKqA//vPxrwuUCXvigpHjNB1MCWP7vBgCqGd/FUjCM3EymcNE85hqckA
41u6aJWzTiwicCqPZIq3eh87ZTLn3RbRx9DsyrLrQLUO/wZSmaeLmxk2Pj7dX1QpiTq2S9y9QP2j
yXveIpo+PPltAKrgCw9GAc268OU0BKgU3lobzKTAnECmbwkNHPf4Q07vNG6d6c0xwW5k45ZF+yuO
NcamIqDGzmLfqJfg2Xp2q2butb1K40rhMhT2jDCKX6LGuDTelNbf7C6iSyWv2cKKxxPDfh0tVBlt
xHS5xk0Ec1vVe64RCZK2+TLSX1EQaWorVGErGOEo5Kd0iWP80ZoP+15c0lRHXhYWmMrrR6B4ItaR
RVyYZ2FrTaS+g/Gtn5lZQJuxNrwEjQO5oEAbECa3mBP3EjptoXQHIeT9qP+qRw/K/yTdQvVBvNzM
Af+yQEmVNrRJsNkFNoYtccuJk91GMTEZZ8LHhAkt+P8Spr3BILNDvXjn11kLC0x9x/p0RVsepMvY
+2apulUyzbVkuWtaH3uP/eSV9n4yAD7sFE1PCNJ7wPb1rxOpb1ovvs+lS+ybrT8T2/1PaJI/CEK5
uqLKsXCGD8P1dLQ4gRuSCyMTECNAoaswpVVTDB+RHYP5R2fHm3SGgXOpk2Ncr0rjLcT29JMpjlS5
hwY+ZbeplsHWrdeBK08ilnFFP/VEiO067ilVtscKyX+vVEOHG6mZpRDJiauRjrY01V6fGzlmdLzD
ooXI2vBe9nfrfChKX/L95+RzUmmgTl3p7T6A+czJl7Y7HZ7aHdNNtYUHqbR0lOMNt8rsQb424T63
8PI5JyWiEMyeoGACcc4x3BL1VI0lZz+UELunexif5rz0gTw0PJ0heF3aA3K2Aix19BRT7vICC06V
eNkNgTqJ9Co+2UtJ+5HLoXtil1rdzyUUHXrmy3dQUjeVsSorQohyn4vHvmDcp/+uOqiYf7gy26+X
btckcAa4Mah3JAtBIAJboAPWcUBPUzSd2fRx//p6TeWp8YgnmCqu0A9ON3iE6afinl6a8XXDMmJm
D/PN2cBMZta4OW4L4gPzBLgLyupEPKVnEulDpNSok7Z8Ex0TuhnsTNCoxa0OU0VRNLYjB73MA9S+
2mpC6nsGylXEuusvIXPpAWsua+am6gYr7nKBF6hnZCV/rmGB9J7FdNrnjrhEUn9H+PESv2XKYRz/
WxlwtXj9t3sFEY7WN6ETo5EPRcpOR/cU8BSJiJUquWdJocYloTJESuz4f8h1vGTOKIpAoluBB0bs
Ge5fDemEgtPX8AdTzklVG1Bjdp9j27fkIa0EyM8jTMOeR+q3ZKU+2UDMZvnKlupfjn2BjLQ+y7z0
YjtDx3wg1bRPdO7lO/Dd7WuJfI0l8h5owijeeqay1IucUnrkNI6lxG1ohaSGM3FfNkJavyD2Zq0Q
sGHfJlx97pLSQavvjgTo4HWpKyoW3zL2s5b7nPGv2bCfWD9Gris51m7UV4zOYArqAv1nWecANXJI
KNtUJi7kyNqRn7BjUC6zJsVjuGR0ATyzM1uoQ7IcBxI1+pTzP6gNB5cSjmjOVt/lYS42eny+M0We
fjSWii/5vXx6l+9kZvKdM5+4SoNwTWiU6fzr3SKJQbuvnF5Uyzv9aOyprQkWdkzT9V957D/xeFnh
AisxfGuRBV5fA9cS8DMbOk8KJH60J5PQ8MjvI2mkGOf+EIykK2RtBybwC3Ehsl8anbFIUrzvjusw
tHZqZUZfHCg6BtJdo7MDbCyi7YW1RWMt393ZdJOzo+W0dQWhz3wcYAIui/QumflK4gm2LTHwHQLZ
0ETp/9ZW0lShSIo7FsNx/xlGImorLlNbiW+UY9ztBc6C4J6T4/VUqC1gaSpYd2FZD8/Q4XAqJFNp
FvV6urPB545Xadr3We2fCxdLcrQePZfDaKwBKsIroNxmeJwBuQ96biFDM7Ivn3ExWv4hO/Fof8Eu
B2y/BAKewR+VC0S4PqKuE8XastrI/0FHVylC+FXOiAsdPUa+U7Ubu2DRL1xXVP5vU1cqh5XEiVym
a3o5fBS+0mBUMwCU8kvbNvkmdKaTrOrvg5l4FWgjnHr0GTG8ugtMQXdYcv1HRFPL5E6nPjFyse4z
kDE0SITySdf5Eq1JhZTC4U+lHlWeb0ffMAE29RSEXqe95rTm4SC/pVocJ7eggtEUXcdx4w0MEFoW
Z7rSL7ocaAWcM8ZsM3wsUit0ATHYPCvqNiOEv7wAl6g8H3VLjkFKEYNAcvcQQdpDtjDihMXIaqA0
IgC3xvaPieTigN2mdMetKmId9WdORRjR3ajsb58kQji+MpuUZKBarPUAck7xDR4VS95vabv5xYCx
QR36cpY7zv1aOHJn3+dxdbygxSRsJDmBNPJdUebklVZamHiZYbjZ+VoBkYMLMadU9k/Q6LPHh8Ac
fS+oKed55g1TavCKR1IgI1ZFIIHqIWXSXqLefP0vy2CsVunVrEshyflwg2k9nRLeBi+BInzNVniS
3HblFK6TzhV4W6UVAxPFYNFl2qU/MB/UKACx5kQOYCUxBfqjxdoGqBEiykneOxtt/pdUEAzNldOK
rlVKz3iAZGh3RlbskVG4J7LNbpxMwF4KFSttgUNb0oNwL8zVDxGVdxHfi3dBGJR0fT1kL8pvOqVO
3JjycFoRMSJB0UdOl0MHFtM3m+4J7zxLOX/fUHPbgtGewLDhHHcTWgWM7QuFbxkdKLVs/ejm0RSk
L6xfGi6FjXoJgKlmG/g1w9hiTN9mOODWiqJx1OeEHli1U1ucvG+4BMYnQjrIP0BKPeIHwIGKjtiI
1JxQtx6URqUKWvMDMlkw1EtaYZOVpTI8MIhPek9xdELoB9q3YQsRueScujzp8qRqGUBZW6jJKXM9
MdDwv9lcIZQVSrV38bFSPGsUuD6N3nwoN+zKF+LhyETYvEDk6SbO3Uy9cugxOcBkbBtxsxJKqFJA
dKj7VCJBbt5pD4n7A8+JmVsXVaROj22wfodOrkIpBoh8OhxGrNuvBWGM8s7lAncMZudhBmIpy0Lq
YVE47i45qICSsBqocy/6Jr6X/eGnIvwywZSmZ/YD7DNhP6mQFGkSwWO2CHmbjyAee4A0C9vsDeZn
OXa8I+o/9ecAL5odAO1OAK1P4G9qFI3nPRr6SFDLFpmsziuKwZX5D5H2z6RUVdEvjYXxRTo9VSLL
ZMdFcKwOElPNT+0iPPzqPwBsZ5wAlBQjiwfOvbB3xg/2h8Lq/3uOy2+7bFjaZCb5jucOSTWlu7dm
9weytUt1Yj9svViL2zsP5dWwrgPQ6xdOFgzAb5NvzhYmtfSp+tDcrL8O9YnIgKF4wtGRtgxXaOso
P+4mH+B+qAItc5bsAgg4fbXOgLhgMfYzcISKvvpl8Ozfig71nAeyHkw3i2lA9fDg/db2XBBR48zZ
NaiZSSEy3u0hQmezMYle+rQDLA+4O6+Pvv7nFli5Z9BWQxOsy7onnZt/9zcDPAsvnRIS4OKkptzg
I7DFUuMDrXq+wD9UFeeJcUyBGUNl1EV82LGKIx3vy8cF6NCSgSZKnOeXosjtaFvELjz/6lWdo7uW
4aBPw0jwatcqwB4Qc2nmsVWUTbAxjy0Za/IlIAd68Ft6+4c9728U1Bivhr3Npn+AgbjmUygxYfmi
BXv5lTQreFfXJUjRBxxLUJZd63siXbVmgRafBog/B0nWUIfCt2UuUpKYC+Plgz4nKGJXRamAVliP
dJ3bGG/G0NsY0h1Ifc9PR1VIzDO4h3/W8jJqGOC/pazE9vIMXmfUK6xxvXaVjeaIogDw5zMEvbuy
GXqEKhP36U3h4Xjz5FU0qsoMCj9xawC/1itm4wItq1ugaAfYx8swOfnaeRJGUNP9Nuwow2XicTNk
WtoY6O8aEHpKyaE9UUlTD8AMrXTf48HJhvFxIP5pzDRCDE3ZpS6zv8FFeso4rRtEOQFOEbwKeTp3
jdHAZI9vvUPyk2A3cP5ZkwOGi+byXkY38nbZ5O2w8adb1Pm+dfGTezUK0ejEP2+GIEgptx85JG31
sfyNVxfVJrCFv4PQx1q0kau7e/NkTzx3LGtU6G+RNgn0SS/hU8PxDL0EisZ+qCZeQdz4ZyQwLe6J
yhNDddwkqFC7icmCWqaQQ2Wt5dpf8jSNnvj06PVDGSuDHvZeyI93zZyviv7cVzR08JAEfmye4kXu
OaqweUu9SAmPfLV0uD1Rzb/d8dZcGyZmHDbE7/2tNmBg2jirDrFWLrVDfpGK/FJCnwAVvG9/tY52
9aryFRJJyqrXb+07ZZN80MCpxrpp0Mg7nde7cqW1UBPTRibWoe+8mUlyk+kFS59E4wAS6/vPsNb9
vewIvJ2YTE98R7JHgcK8zClAZ+/3Fd+bbQx4jKqjvTzpUSDBA2Rj97zBwHZSnveR/rH5Cywqm0Fo
Q15IF6lxQpGw4er2q9Sjhav2/F1Fr8wfwH08uuJy+OnD+E38SISs3jI7CE2SwIzzmDQ+UCx+i8K+
xrsp43AQZfq++Vd6jkU2oyKRXz56Aez03jSZtNt4FGxRzBjwLxzMnXZUzEyMtxLDHEzq6oA+2yvh
9E8yxmvtPmw+y/kAvSbjcmXj9d5cIkJtvKesik4nnZM4K1PJBIIB/pr+H1Sa4wObwe44GgeIwxQr
K/lMuVMhdWYzKFaCfrWzIdZJEsn6W8gcQKc4oZQly7E8k8ivDBctafw7xZJp9bvws1BHTN4GnubB
DBUpW26vlUEjh9h1LfUnxZdHekAYoJreaWQjg2OAc7TxnIciyjdHPi6bMmw0eYThDbGFKQNsM+Yr
7CjynUOmrgswdQK7B9xZi6MO6T5QDI9+kO+xZsAfV4qrSs6ZZY1+wepDOAxCLiNoDLX2AS/l18T9
SU4SP+k0u05/9iOFsg1g/YitagRj9BPi7CaWlfbo2+L9dqAZNI0EQGqaM3ta5AXcKOrwv+Y0ZLIE
XJGVONWNBz8ogGp5In9IQOCvKEjitGY51fcw2fXJRkVk1dOKuaHRylgC8lGV3UriqjgZk8tM3Y8/
JNn8KfnLRFg5/P6B79zHG2EuVEp9yJ3vSYrkyjRebmM49T9Wv4Tqh99nZ9fLYvrC34akjG3LFamI
m+YioKvL0TyrtxaaK7xWftiy88ufM01HjNmzseFEpRZbLXogTKOvrvo5BjOjY/uROQ7ei3Mxb0Hv
Y4v6Ca8hSP3Nr++B00tgloS4waKmRj2KXWMH/91sc/8fpMJHJ8DU8SFK7AKYXCTdgDV7psZQ8Z66
OOb5qtRS8EdtG3jQG2eO8EaGX9VT6T8USwy6dOwLvV1FcBUdcbi9VTi5fy0+L92dwq3ItqM/R2vS
fhfz5cWLL+TZnbDJCy34jfTVBy3un+HLcJ00JozkgeXcKZwgw5Q9S/6fKAFUon/OzhdxCGXV2sjL
OHyXFIjfxM15tpZZCVC7BMFJ3iQZ7eAXLHHrSbb0TAPIRJAeAkOEc4SJIFLcNaQh9AEoUkdMRLaD
8gBsiPnG+6J/aLC7SE3/lbohoWiJcB2lNqeMdXiRDqjTBotikD2erJ3gzjLFyk7SSMXDTncc7klL
n6f16H9UQACfyDCKYQk5RnRz39l4W/yqOWxzNGmXH6zAgXEzF/WIejsZV2ceX+l2jWRm+GJi7/6z
KKgW3uNNozWMmZJMoKhT02PP+Ag1T2MI8KNtRTvtBy0FZTP8+6Nsr+ibgwRgnUjd3v6Asabee5tu
akxUodqE72QritlA535TOnGjpX5u/jZngSTO3J6Z7TL/23gv6AI4qDlUDtUQX1QeO/cEPBHmG57K
RRk1uhHEMV/ecDftMPBNWiUNkIFRQXfNC+Xxhe1IiyhujEQgByf/cJBg0GgZXW6dzBEY0B0rNZsy
u2dGyYdRyBMUqypae+d8s3Kjsh9tzbF9G9vAiDsN6xpyaIvcgXj4NYJ+B+YfmAZf84v0VL7Y8JFh
33TrB8FCkrBFdJmdAcOTA+N/QZDk9qft3TYK0NUaJJYvEDVYboXry7LkNfZmYxQJJHaLFiUg4P0+
XEqpchwKQBanTXw/SE4mOUoGuLBI+KoJuJ9xBzAw2qFu7KX+t1yxHEd/zG5fP0XpD5Rci66Ou5wO
auf3p9YOhtGCaWIKSFpFwU/XxnPLKwVek9rI7NSreNIgh2xK3j7wlu4dVf71zbWEjZKt1ktVf4u3
gVfteWbjdQ1rdkK3Ezo8RvhzLcmH602lEqhJkm8c/q+73Dn8bLjQv8yvvRnYZmdzgkl7rCTAh92G
U60eZK8n0p+OycRc+dzYiNLAF8uNa2SHwddMjvlFx7kVbhe/cPLx9H+lHkwUvoBcX4E+Gb2VRShJ
0z59Uv2sNpW0TO1Rq77bLZby8cRma4rI59swzTKiUeozdhObbDTYT4H2woNKz5HalSKljPn2aoS4
WcxFEuY6ZMls64SuGknCRIOhMNS65azsxcX1x0Y19+ACEQQCq9dMgFEECe1yWSZaltaot0iyo2lB
98BrGSsGBOiIsqtj/pXv64ReTplAscKuuePifAphJCDASjgfzqI5/PAbqEhZDlChWFmIbyDD50Bu
gGFV7yM8WDgTVZqvwJZnVzecso1fSy33Ajzwuryth0pTzrlo53aKys9ik82n4jBYk0pU1Vrj1cA7
je2Rk643groWD0OuJpFQ7f3ujm/SdKooPQPWDkmxoN4xVM0fflaZwuQOXijub2D5T882hOq+Hx5a
25TO5Yn+5dW/X9/T7h2gjldAUmgOi1x/oukq8SPjmSju3yKEfDUmGaZf7J6YDfmG9QhjE2GowVQD
fDoG0WM96mO7vh3aT2UBjht4w/8k5hAI4jnlh7/xXyFo88mHjgmpP2BaVV14culcOET6y0QGHfgs
tA7XGdi9T4PLd8tR5SAPWuBvWL0Ba4GNwUjT06OWi4JDmgdAdIrv/xFVfmfws7yNNPd7sMhwt6gK
vGAmJDMLAqxZJC1pmfi4+wmTRY6iCLg8MV0QmgwrZv9GuDW9LmWESC+gLImLnW6tkttAKVk1Lqwt
g0FTeCSNTAYGDUAwDhjyrAUqcs3JV/EBPEeZOSjBy5ZW0d5P86775fIqjJCwzRchH6dr7aDZcDZA
Br2+8bWAK8A7MszyRFXlyHQ3NBs4G9eKdCgBcI+ZOZoFl5U9hhCwPG4YEALnVsuDVaCiIY0F8sBz
8PsbD0uDiTLDNqL99RLLS/Qfli8ZAktuhKCjQAiaUglRAo3yWAu9RO3E1VuiwOgsdLhBIFqogNhG
Iu9oHWBE7ENQ1/T55cNu4yK5+9ua1WK6d+HE5F3OVaKd2eAs7aUlixydSvL/QykUktBk3b3KxyCC
obatg7hLQhjfp2ZSmcK96ir9LkNjQ44XecNR6+Xr2WvbVcIHtwLiSxdXUWRcYPmNf6z/XYR5C5zl
4R+Jp1b1fUmWovtAfRpWV5xrPy8PUAmkYORovjvHTgUQ4COLH8OSUouYU+Dbg5OTndJstPFVyhBq
+T24H6Kb79+j3WdnK84iP2lEifZcq/aa9zgZme7w1q7Xu42cJynnVzgres+nLelMEGfIVldK+Ag2
WiPrfLjxkhBdXCG/Y6pdFEixC1mCjLeIGo4+lwmxbm/RRZcsgDlnTSUgdxT6nWL1WSvk9dOCR5rd
exINaDcDNLwDuiwNYrjFceO/yQoanwmbNp4fKywugjVqVu1olbEB8zXXmoOtncJ415NoceqpbZsH
ZfdTg8zeZ+zchvKt0YdYXu8ufSnVyGxqYnkFPHhx447317HprDV0qekxTEp1oVNULKXshah84m2V
dJ3RqQi4McCU+pzZ3QKVi9rP5hZxk+pZrK65rr7SYGwEElqpUefXnlZjag/4vOvfTCVQRB43Dm3u
0VOZ+XsVRlXQqdGgiYD5AzVSRthRHS84E3rC52fU8j0EUteANlSjgfTHHE4YpAGg2gOqCDoK9Vv+
sI1iJl9gckbjNBiCokdSWHx057omq2xsGYRaQvjvb7LwFnBpePgpTcW5T/D8tQByD1W3b3W9EQPx
SxRAR/Vq7Vr4b3OBWQFfoaVG4pHseMqqIVAAVL1DrNqF/iJ7T03/CsxJonYPofwJTp6sXPCZB2sW
paw0aRa/o8Y1SB+Q1f8CX2oM/Sq88wPWJdJb5peOEbzDcD3cUxqeqVIfIneCuy1ZIidwBe/RjE6l
Aey2VL30lKbkuhdIYKPM03yQw4JNAcD5V9uM0mWJKk7WN27aCHyyQDpRtubJaiwS7d57cUmzvB8D
IBhOcDNQF7zm4MkW4VkQZU8hun0OqRA1Wd7BgT/pTHIyhPITgsNBldYE3ukNp4+ZeuLRgMQTFXex
U51QzxltnEIo5d9DDkRPLm/wGnHGhSPQbtpE6rPBF7ReEzjElTjHUxP0KoJL8hVWpOCl1UmXAQNx
m2HGuXnc9soA1dw8g0y5fpLMHL1j1MyozO2DoQHdyrmo2GZIYlXD8sEMrAATmnMeEPKeVacVLfMV
YXIsoWksiriYadTH1l/2Wx4Wewa3Io7dCek18gaeU0bvO46eMUDmDwTv8IjDLFhQ3W+ztCE2xMGi
Yx8zJdGjLQ+4V7yPGMueqbI7kmQxpbgNQtO2WtWog7JVTcgEzuz713/+aRvWQ+8+wnolFcivg3se
iBQxcPobva1kVbUCuE1VhqcfFlt9FvwW0T2KLonZmy0HYR8eZzc6gEpnrO0uP8/6+PfkntEC/Dsd
lJTgzfrrqrykDz6ak9oEYQ9ot1GZZZm9o//4m3UnmRtz4lB9I1SMoVcLMgvdD0ZJMl/9TvuNDMam
vju5Cj/pU9rBDGWhW3zy/9WPz9n+OV6a4IrctCF/sMswNyAJ0uU7eRj+qy9Xt1ME4uuqcK9lEp5w
q/FBwcswfND4SYBWlszRu53Y+2pg9Oe7d9sR9C6h+l7aZF2dTsJYLKA8X3t+xe1W8qi1CBY5mbQB
wgZZtNfqj4ZwMf+h9FrCbOrte4tXEQEb8YqjHFxhgFe7ffHbrLNM5VzInG60nv6cQ49naYj6zC2s
3pNSpE/zsdbJHwxBajvc93OLF9HmvaHKwgyZRImkwFqnCdBcsG1aUSgoplf4H4yq6u2escCytMLl
c+OnXOeKtyXDghAEduFiYSpFK0vxmUWFSmbpOCBdB8KvutgBahiUQzLSrl7Kg1hVn6JbM8xDOu6h
NoZZG+YqMwVdsbP1Xqp88sJVyPFIuXRUtrIWSWxEexelxTHKvnj1G8u6OTQZpSiIhk+Ohxk7ilrD
d1ILnWpSCk7tp/bNwnVIyOUQZ1WIPZazRT3bcTemLZ8IClWVN8pvtNpe22PFS/sHGUFr4E/iFicS
/X8bz1Jb0n16+9YGDZT3b2mFCMUBYAoKQDpseQrrxpPXjvkYXfZjEQeH+LTb/ZZ+0rrT5SsoeRD2
CArEFTaE4NIZZRw6r3B2ZvyCNx9MN22nfuk1GAlYAth4eu+ktVncq2HIeBiyjxZw1y86ffh8j0P4
CawaygrmFPpXCNbu4RuBxAMYR+XexVigFuSvUS2a1fI3wv8tdRf48n/KSY9lGA0kHgqTLFX1KhCe
YYvNRXJP5khTE4WKE7/iraQ6ChhVIjWVHErXOPVmUc7W0+qHZ3gMqey97L0bobq/LqvNGAxyQfM4
98TK5ocbMyG9Y7HljePYdG91TU2ysGL6Tkl3yQaHZu8fYEdpbaHNVx28dHIHMVi82fAbLYwckWpW
qma9IKdrQ2Re2HtIICKEFYGv1Y1Tql5fPg2BXg0N9floFNy+wlhGSDXAKK6q4kl22qqMJsnlEdvy
/Bt8QGQyTWOnAQjqLyGrvY69HEHbUq3WcNxX38YCyMaUAab9PvMKMiYkizDKoFtL8xxeKRIRSg/Q
CsaZLKu5AW1Jbsf7JLu+U9iDGoF6plTCNvu7iugjoS0mGQmx/AKiUdQtsj3hkbcj1zc4BL5MNlTK
EfU/ohMd5qCAY3HtE2Lvx58Pe+oiiw23a2coHMoS9ItADPQsU/uth120MHeZZUkTrHWvAAoR2iOm
1hyXuC7qByM5p/YKSgJzJTUeDOC9w/9SAiKf1Axw4bBV5nF7LIhZFnVc/u3UA4i4cA0AtOAo6Wgo
w2cRJXkfh/bC7mSx+AjSAIyXbUdL/3ELTQXSyP4QKjnQy9g+4X7o9OQe2Q3AXW4P5m/tTZnaPZTL
VowApGq/P/sZqDaWKpotMlQ555dqpjWi1T9dtLRsRIs5+eA2+JLTRd05md6Xd+dUOHiKTalv9YdB
4Uc59OlMHTKhPeG2fVB2cAGVAKIVYILPtXUvePpmlFHEcqICTqzUyryqYbk+Tkjf40PflROR1dPi
kpSf8G/BI38DxsXOOlN4770p7KYxhHdZ9mLySSHiFJYJLMKakSHIdU8iEV4oCCcUzTWLgy+c/vse
xSaytzaWk8W4hMm1DaKgbp/O/T0k5oek9ZdRwx2SlpRC36fNbBm2cDckMMsFqznsGEYYjDiUIUCa
sJwY2Agt+b6H3Wj/fzi+tWHvqgrmlF1j81xVCIuUDhy/wd+lBnLuiAgOuCoh9vugWsnOl26aSiDz
8Ym1RVYHj1x76xHf4YzLG+zXHBIufm0+0WjkaH8oXfg8u2Ewq/7UnTHsqmLDb+6RAtikCgNgP3WX
6SKcXiYYPytKV/bu/Sbk7+Dyef1fxFhSzOB7lnDfZHh9717Xep6XVo4xPf0Oqmh5b7O8P/1BWH7H
ZAhzJDBZHteZ32e3RXOceN+AKfOSLDj78eDnhLxOuYBYASdMJh4BaGoVZ3w5kH4Oj/D3wq3i9wY3
HlruDFiC3gSR67q0SMKxJPLLPSoNTb6WVy3VofbM+ECtHHB8QiMGKibtW5cDKSe3NSMRcHpn4enk
Sy+/QyP20LnrJr/lqWzQhwp/JwANXrpQPhnyZZ1zf63zEZ8iNHLyHe7fq2SryfclJRYttns04sm7
wlXwjoVx52AW1weMARdcs3hb0dqVHKNELetecWggrUnlGlANXBEv+2NYYzcEb0xJzJNRu76ZnArL
d9NijhSuQf6T9wgSBTcCBAOvWUZoEBkGoFooPQLK76AwJnRTcN7gAgMQ+wFYqptaOPwJtvrAf8oj
1N1mekI1iKtfOKVKoX0wO6n8EehCHDyvxlaZcgwup4+eSyR9FDvsBmPNsNjFZnaQKDBz3gFPJ9pN
L9L0sv6Rhj3vfn45RjTzqpXi/4Mw92XBZQMiYii2YuPHcYtLLdG+DjDu9ZVvItNVVQWFAGemxBCd
+QT/xl1GZScBG//5Jbgyxsh+lfDOTF7EJlxvgGNQuRk4AzB1xSv/cMucrVbYEGkfnDsrXTlVYcmy
cJxkxLFVIKfbwxY9EvbS9a7qLYB2lI92ntJm/1RisGBILGmB30tcXvitWtuYlhTBzNcSbu3CuXMo
EWwt8o5c/Ihpd45e6gc883TNqSmVZLiLO20GqGHtcqAjl1G/cgSrD3DDnbEkKhxidhFV/T0Kf2p0
tVC6gWLtIemgtP/xuOTa68XuZ1PWyXcw5JuOlals3W7Kl3sL5ZpY9ylldwHZkBBHWEH7CO+Zu5zF
Q+StpSq7eHP2sVGx7FMn6KpjRNwFMhYJnrBv+NJcw3kxMet84VQV5+gr0YC1CkQnFKPYKF6PMfpT
w3PTcNHmxFae/vSrDt/RhxSkDuBk80Qff1gFZ6AhmYeUV8hWPhWvJ9f1cQTb7EnbOGIyAxO+mrji
lPswn2nbF0ZGDp/nym/7vEtPFKmcUAwksOmd81Psn9I7qdndcZRc0M5higrhW4TCd4DVDSWiAqV9
5gfAYBqVag6CBR/uepwnp2S+SOTuB7JVQmOlbehJzjZ+RbCl/EhHFk+fDfqAiWNMw5jCUFFAc2ON
gy1lKBgpnjfA96qkILiBKznZALuIHJJr0NgnHquFk7xHC4ZO/xXsGzoS1uGKbdPPEaZckqWHNYei
CAtkBpD270wKkDsjfSepS/Z5XvPZg8gqgubdTkiFZHP5aHViY86RTDNcpHLLZXg6bsPnwicLZX4C
smRe3FNy1XCJ/9ohRcFH0oFu5XbFT8oSLNrXidHPr9LNn+Ap5SqQi2zrAomq2y4PqQqDV8nQ2rT1
c811N9pfUSHIcOFoujpVNor/sQ9dUv6Kx/ag7zro7vhjQHL48PUneWk4g0nrS0X5x2ygg/IK4O6D
1uiVTXRzd+SDvfOqblwDlZHhB8tKgwKpCyrEaG8Incg5fInVEqbUHMqLwvEom9/er97RIuTysv8i
hvHTBdwrZ6BU3JFm0WIp1AB6Bow1DzQXjRcYaJCAlM0OkqynsihrFJG59njDTdJ/IzFxj3pOEia3
K6EYbxq2eUWEKD6ZRUfFLieJlN8T7Y7zak8CE3AJ6NHOptAaZ8L/370gyJznyzB1Kgi8l0hd7Yl4
w1TgpUXPJc1PfRs1TUxLj+YGqjM+WB+/m/c5vGh6pjX4MvVoSib9hsKIrIHGqIdCaZJfb4f6P5lj
4thEIwKomHaHXXj4P/yPSO5iRFH+EJyFz9Pg5R5/SXYSIIjgzOi+/4IhVe3kvOdJ0tPwGAdYdu78
UO0v7smPgyNDmeRPfGUjyV8/nyrPblrdhrP3d+qKsFGqhPnPN3EUgTzN/mme8XFIpE7PGhCZkesL
lYs8w3GkLRSEsw/qyikOQcacIulNeB1SOi+jjPWuHKd02Kf0+FFv7FoaiRk36iOZgIxA0uBzkMwM
wK24KCEB6rWE1e+dVobH7ttfNEDhH40iAfGMRsyenhnIoVE865WyUqGla2yj9G8v3d8Nz2u+V3Wt
oP2N+q2O28D7LrjZ3XSOU/X2RN2qW7uFinz1uVnC91NnI3OKP7ARZIbWcoHT8JgBo19HvmVYj6Vo
bCyCwW/x/RNMxeKt+QfQvDeCS94EEXWbvSkJEswDI7AbHmXrFqvMI327CQPArajh+4gM9wAWDyEC
omNp7MoDYnv595/vnRcV23ti7MkrCyDpcNBQEIDD7Lmgvdrmyl6Bcwl/9/QKJcmpG/GC2qI8SExG
aLvvFFUuNf6RA0OEd8WOHlJ2puOIvvx6B4b2rH5K+5QB9uhWjRvOmFMrBTZRt4mVeW4ngZydOmQz
ZDUm/T9hj6NsegFQUFqB43LvTFRaN0AJIlsktuWnaRk3n3gBSVsSozLZRYUMPLO/J8I61OXrXTrU
ehhABs+z02nWYp51ereZzuCeRHgEXe9JUHPiZju7XRrwOUMA2Xe2xmUfOFr87VbBIKhfhCqQtdhZ
f9WUl9BG6gmB8nas5GQba2dtr6osDiiEPoTySSwMSIt3e1A1cxHOP4p20GobYynS10214AIdutnT
RKjCxwQmTlv/GjEFXCYi3ssgRpfsODq/ZKDSwuxFJ2pBER0fLarkKpa6Nsdyo1Mf/GkzNnTvIOgq
LNMWj29jqMOoXd4SpB5VjZd8gQkXStiHSAtaOps28cJ+6gJoUF7iN21tzwhpkqvE2HSG19ApzbZO
4FiVgyKM67VP398kAma9g5zIvm2lZ09WthL+CGI+xvBZL7ijwjmv+q7wmnb0Bc9Bvr6j95odmprC
M/8yuEjrctSuLkjzI0rz+RcK2u2aUlHFWEwysJeuqw0AWIeB44TGnvJpIvyzNZVhgl4piUz29xkv
vU2epAuFS35lB85atDDHDMXTF5FbwG73O3QzKBK66UtrJfgSO8Yll0QHatwI/aSUH+UAa2uEYLvX
aa0m0rrJCxvsfkndr5I7fIAId8JCHgYsd7z4n0lX13sZ41fNiejxW8dI6w+PQJMREnFX3k1kB3i0
xH1eonY8CsnBm4AN8yO/1pGyRnrZOfjOW+9xbXzwjsHRkph4k1uUV8E+BpJ2fHOQr+9dmSUja3CF
8hJ5ZUgZFpT5G/PFUjNFU0ogbnBQgpwjpbOKU0Tq8CtYYH3FpSeac3RXAIRsY8ARuy2vt8ArDvkM
hsjVuyqICcTnRDLO24vIdY0Z9a0nd2zDdsRVNED9FdQ0MwF37IwpSMZ5dwtUsDBIrtLfj4l8eWut
q48MxcKKo1X7XyJR1NrwMjJwPyKiEq9aGrHGuQPyeygmtsLEHbwDWNhgDIyI3HmXvP/7GYTsWago
sdHbitrKLwZAcZLJjjNoBFzJ1xI6pW5Endxmy++nOEMPDofZbWJQwdziyOuGRGdLJ9UTakqc1cjJ
MMp1hHeE5DpHF8f2+2uTT2+160wyBAP/5DlIQw6diJ+XB1htiZUybdeSc2MNunHQUawamFoSSAad
PSwFO2XqZPnosBsnzlGyYiM0ZDOwdqSC6woJBKHU2eZTEau2uCELkU+yjB+SfBdgEEfGDyoK9FXp
qXwU8L2jMDoZou+an4SZRUSkNehbSWDDkZ/hfpmCzj9PxzeUn7Yuqi6LHqnXVAbvwVsYNIGbIvG2
uLZQ2XGsYIP19R/4y++dyfwcOiwYSL4fJJa1wXiQO+zuHrPj4dLpKHB41VG8bIv9s5Nz/X7ThWm+
49qEA9MWhtky3LVEFjiY2ocad9yAgIdlKVf5qdWRJ6Z0nI0xT8uyoeo8RN0hLKdidPX5ZtYGec+W
H7pYlfoD/Zgh8dyKsVoqB3LZL25Mb9IQNHQiHvSgdQNAfGxixRFVPusLiXUF6UdZrNiJIeVKwxvf
z4cf1448xdz8amlEj0fMIA/f8Ocj+PO6EAbnPYFJo6Hz6IDr9CpvVfgMr6tKgzTBbJ6TyuBHgNbX
QSeLZavwjM44C6mTttRHbR1i9QqdAqTX9ayMAe8QUYRGlz2rsEhLhVxS/9BA+vnqaz31yvvGOmXP
X4LgLEVoPo8604/x9Y6IHWLYNa3cZ03keNy699T7zRvjGTgZxSnB2I8DQGlt9A2uLYBNKA5uV0OR
dxIE3mjRHHuYjTCSA8xwJOePHJ7nBlMYEgOnYgkPqT3igxq2sIezZl+1qz6I4pXnQEYcZUQU8ciE
WlEyebsyzYgOv2KILL5oXZ+8+Itnqi2twUv4JipIMRr8ozVgJMwCyDI6sR7SZ3/kynnnYpjZdhfg
ABq+pzT1esMmFvewGZ7FJtQTjPUE5+TkHP6KjKpK67f5kNKkJ7B3OBRjUl8xWl+GzS1e/nSkr7WD
YAoCVX1Mcx68CdJpW+in0Y0kkZJm2erFaa3xWjuO7+IFcql0dcKmAsruPmn+VjMhOVNcKHlS8PlP
ABZwt+qLEvgEEMaQewnmtylIV7zVeQ962F/YQqRPjt4UeMOn2RUEeJnaPN/jexjP9hMTnlikQJ20
tGVgEaq3h6s6yNAXN3Y62kdFR/O63aa6rEaiiI+pBU0IFJFH+t1J1WZGuStLiVpyQyiTNk1nPIKV
AesM88MAVo+cjZLfWipmSDw0rGOSoCxjT2TlxHe6Gruqif4gryVsm5kduPu/CufrxLKebgz9j8Y/
H+jPiwlhBx4BhBU89vVZ/p3Wbws2ud7VEP+TzMINGdYGiUocsMoVfzVtIN54nwPawDNaVMelILlZ
TlTieX0Z34P8EtZWuBPc4Zq8CAwHholcC1yp2HE/ItQDYDc8/hzvHghBz+JZOmGSyRBgyC7zOAeo
W6Er3XYa9R7HRbqdYMlPpi9/4f+zef7C20B+G0BzAPBNursizdjHSN9sWxuUQOUJi5DPLeworTxo
/EoqQ4m1kgc7m8DngVVBTdwj+eceXhZ/2DWc0G3TAMSOwpp+Xjh7n3SDXOOSaRXpfDwUqhcAbt6Q
AStrwu7iDLCJAHiwcGv0XOQwD38dxsbaaS9so7LoRZ3CKMhFo/dUCxHG2CU6IPt1hoOoDN8LQsaX
FTgdN3s0Jp1aI2reovikIn/BYToKMuK+LRRYURqLEPeq1yGKoyXrqnRqT8cA2lJ2dlfMITVLOag5
6EbsmhktX1OwxtDuAp47zX5j9o9dlDVkxqHRrpnLkZQmCZ6bkUpW/6/deyQcU3kaJshLQzmyx8nL
sXshlvzHWQdnK/9ai7gaw6xxZGGMTMxqKzIUpAh9vuMTqfEdTH1gE90VJydPurZ0MVj3ToIGm6Hd
Vnb4Hi1GdB7NEHGUJwBmP0qj1+isExo49IAf4XawyXHPD/GqRBeBlZUqIMmDy/4mM5IubmrGXI7W
orZWRyLMGr2YSWkxJtlGZ4S2oRc0rdUNBr6ad9XDGGrTao1MIfA1SleBMdkkizf+E2a7v3SPdCKZ
8qRHBAtyZhgAvKyxLwIDIHeCX+R/hgmUkdOICakrNK/8jbkuOzr9BRAJpSVlRfPP0+1h2f0Qd0K3
kAAvyiIwXhjPo96f5TT8DfcXqULGuEGaIl3evYX86GVd1tEmLh2bZSaiB1x+7/+mkEf1p9kG49kt
cCx2Wyke8oNgyluGjsHQfag7YPT0GQ1oc8WG4m9DuKEDiEgxCwWPQJ3uK29uKo0Gx4Ls0oOtJDky
UVsYMpVOoJpwNt47FAbFeBifKv3E7TboqaJ01+SlNYwHalkSd2texjnSBEb9JEkGFaMI2AuN/xsZ
idzGxwJ1B/MxQzPwKOT9lnuZTKJTkuG9U3DSYgyPgJ80wggh/unfd8RoPd+/kr5aOmG/Fz2B8ycJ
I9cNRo/JC4Ey0OQNBWjSGVBbb5Pq/1n+3nX7tqeLMRzLn+hYjOODN+H2YzGJLL8nSd69XuZMuXae
xn11vkK23QxO6TtaOcm9z3DVOVPnTN5q9k0M7ulg4Zi8nQtKGaeCzblx5l63436gIxh5TASVdraa
Nsb3EVh9cf2YiXWy4i0jU64tCqsd9CEtuef77ROuNA7GyTQQlp5ET9VJ3WISww7cyNZpXqpefKUL
EklfjAq3rbk0ZWqXRZkADUmDiy5FGnk0t1WiOyFW9/pvI1Vsh1OprGXKsAqexSV44pxYqFrtoLIp
EDpu/GMYiB3Y43lYAFquWL6OKp0hUzFZ0tQ7BjOp3Tt7zq0c/cRESCatWuz4ueePi25+CtIqq/J4
c7GC1tI9/pGZMLqKHTWqUC1rDzrYNfWpB6FMvRSojKLklfKZIVQoG3TClKMyeC1gds+c8C0bVZBg
jChQ0B6U1NCpRXbNXFCpilKvfA0o/iLVVcweSZl2ZxD54+qKprFHb9Gj3I+eEDBN1yAlLJrwrV5u
y588egEhx/vEI5vPAGfvJ8u01XNPgxEQnIuV97yoeWCa5UcmI0sjCaAzRiUyLUl2qC71OTApVUHb
08DuDdd0vltaWTjYuT0EemzDHPaKQ3xxzbL8LPVElEXRO/T0j2Flwhj9ad+HTRcT7+xpl83zjHFl
4R7SuafyLxVovEy5vsZg2Q37PUXWCYMFKK0UEtUcDm8a6vWJXMSWXSwY8YJQ5f2iXwpX9h+h/t8T
9HIc6OrTo9g8zddecKRicXk3Iv/9cWoDKlY5VedvsvHpS6ZvCCuoK927nk/t8jT7Oa6uVV/Blqs+
WkoJ9mHDqfVVJ+a2xBbfcHCgnGYBKuQlMLw6FKZQ1YPq6XajQL3qysUnFaDVIrZxNWkqncE+iTvk
2sSHBhBraQ0aWqjLXvxdddAnROvUKyUiiVFLDOXo9G0YmZHTMa66CHrqybNHYKPqLvShdhF8pApA
mWpez3ewgi5NTxU/GJtGsXVvDUBRB+pafz64PmDEpGcDuoo7w5BSBlskNCn7tP6Xj4O9h57OfCUH
Dye5MY9FxSXN0P7yjtzbkpXYl8ZN+g/1wA5xY1gzmP3GPnv6wCNI8OBCQhmAJOo3/ncKwB1QjwNo
KXtdGGjdsrejVp3cUwOWmNCu3UmQkuFMDVk00sFA9vbydhNNRotXGGo66OZOZey36vtU17N275X+
Rvg2YP1S4ztAyxf42C0CjWd67AJSlrgP0YZB4PJyZoEeO8puFPnzbkJPAi/pCmAAOvwzkufmlSXI
3MpwfLiI7R8LoH3/WK5TTKt7MpzaET2QR1i43CHdzqC0nW3YMxxyieQNjfUKUlpi8oMuUwskeDqE
06bTVqDxKrephhWvhlM1mmgXKW3LNgo/hmNgO3ypxix6RRrRXhax1+pykrurRcYPcS1tourOG4gQ
Jnt4Y6Pmdo+2oMJtVo+hS228oxS5MpM5zf8O8p8jw7yoyIE+Zqc2LXSLQFNwYjIiQr9hxECTXNOu
otixeG1GHikEBHQkaySlCgiEretR+ctAn/V7cR3fDAv0BZSSbn+E+lCsy0ixwlWXKHXSNcIFJHvO
M1VO/i9CdFM7xLp2e6oA74GtJCXuUEuQoug2J1+5phiBbYkI5p/eKtiY7zSYov9h3K2dIa0RxGTx
wXRH0J+bu4JDeXkrl/KipW4wCAFRADLFaDQ0f2YCuube8dzy9u6sINUpRivhjqDLaEYz98aEuLKe
fWalYLeaLcq+cHUNBzBCYjXFLegO6QSQqTWQKlPJMMDajkoGQTb2FsFArGiJ8KeZMx4HVmqmJGK/
/Q5iUe2AVAwkjsNdrEF8s6mrFlmpsXxsWCVvWIDZak4nJOLaOBV4COWDhkxyofq5U/BUnBl+80SK
xJxxGwAxcZNG0sIY8bULrv3GEbJTFy5x3m2PdpH/Sl9+b2vdp15/FPmAyrDn/8DpJSMwPubxn4du
6gh18jrV98LaCqWUuXvAq2igVbepk7zUXdv2UgLHDMiJZmmT9JuDUnswi9pS/OYYZ2khEMvEt/W6
5li1szllxlY1Jx9wP+QuaeiWzhUWePPb/XPhRKeiNJ3Yk+IrmZqZUgBD2YpbPQRCa0t/SLwOL0s+
p51ZA15Er3gst1mdj4fY7ZYd4sbN0q0KKklScgo1UApRTZd5b6gJxik7BCHBlTYXyhRdyVc4B3uR
x3wH1wBZK6j1wn//sZgvUP4EXGFqKd41uAmD8vT5wrfN1jN8hIdthA2pE7BaE02Vv5xrJh+M98XJ
cieo4rf9hOF11GLIjUaPAGB0jardnEFJnNnsssPyiDZ7esECASrh/fvuizPrTd+pagtWVFjI4cFQ
CWHCWXKQW5QDw3kOu7nuVyMRhlxxiLDT85SGNBdHplResymAAJa23ZX8xi7vNCDgd251TD3pKpOi
immQk0jvT7b0MpdAqL9DgVcEwHWwHZndaEIXfPCs9Cp8UCI0KZg8ET9OZyP4t9g8CYGc+T4LIVq5
fC5fzdO+RjpBWMbOX9remBuDkC8BJ/bfnYfljQByY7uAPqMgcecPQHblFA4nXCaVvP6d7HB7ZipY
KJFOAzKQAiv7Ogdbta2d4lQBekZ25vmaVj67eYowEIRVKG9UCSJMQmPSi/pNMPA5KuXwwKUlk8nk
VnLyhT3WsvygAPKv6AYPNls5q6GZKN/iOaYcdiZFTeGMS1GrsHRkPrd+3ZFQmnxT0yPW8WD2W2qq
b5Di5COK7N/13kZh3OB8v2kAodn5iTFKBsrIYOiqB//8v/THA0eRgrk1KOhmPIpEh97bIrFcdZ2p
Yn0KVLaHnmgZDB/yYf/39h1V4BnTRE9+FweYcJmt2uYhIkuSJb/HESyebz9RUcwUZx181bPv5KZH
3wRmuHzWrS7zWD8pFrfS3l64spp8590c2LTjqCJSbj+8q7vrYJ7pugMedE/l2I4GCndEaaBkpsfm
nji9+itMEtGgE7dkX4PJ3yLlWMAbSWnGlxnTFDkFTn8dflod+4acbd2L8hyZfvJ2rK5gtv4w5ms/
dOrksqKcALICMglBiRPUWI2MdD8UcWcvc3WHWB2gdEDMhcBefSHlGyaxT4b08bNHdtvePq0NZjqP
Niac6ovfSPWJABSvs52rguSCqJ+3humQZYZXNUzlhCV4X68A+g3rUEihTYM/jXzjUAgQaLsXJXLK
c3NPCLhylLg5IRmq++M2gyVHGg9hTDnRtXYX58p73i5wqddgi+tJmgaYeAMsh1bnToZ9fCjBe0V0
EBGTOTknc8tPAOWkQucHYjCElf52LTUA3xS7Ti9WLZPXASo2trHlMgzjx0TH2A6WnLM73fnj+vTU
RU8nR5bVgLUDg2psvjJRHbNjcnqSeDZf+2y15HuACbRkRdCqGxXsaRqcN9ZueUv0+913qQ2b6qVD
+HRfrq2ffsAh+aVB5c8rrFIha5TkzFxA2XjZw5GaoFJdv60/hlCEdLcag4edC5q2gsLQUwHx/gla
wN+9u4lxL9zsglSbd7V9QG3xOhMJcg680NA/EfxcoKPwgoa3t+TEZEHg8RYIa3X5tYZcF9FpgGMG
1SCT6nMzYumLJOMzrwCL9R9UG4KvPcHDYSE74gQRvYmQkO0VKdg1E4PUc4bddd1Us2e2R/ACMy1k
SOUlk8AihzK9m2377sW8pTklud+NN1LwIdwVJXN8YQBlOlpzj3YB+LaSJyn3rZtHEUVhe1o27OST
kCw2nhMY7RGlskRICCyB8+OSxKBIRcQOcqoI9Qi5yGud5MyGnr+YUdVOUic+KV/uNkCXx/piAMbm
DkK1qe5WoQJkVUufskq2R/BirDgAGiqCmXRhgD9EK+hm8sOdKGqNJ5vU0D9AM/DV0x7Zuyeq6s3Q
TRkpZyhBNmJ7SxTqvelr1fWbH5Ay6fhNCv04tet0NbI59zsi7kxmY9EZob8AwWtXxldcmhPVt/7u
R4iVj2LbwbV5Ny1ybTMXhX4a7D1WWKYq01IONC+4rFl/apnoFne9SZH4GMaeMpnqaqgfn14KqPBR
5Gjt9B7P8u5d0YkIIuY/xSNhAV6l/6/bBiueM7QKleYKc+8tz/rE2jX5YQkT+yMDD74ze8xedFBs
u01iN0ztyouqLXF3idxAYmoWmz33aVh8CsUfv64sebJ0AhKhn+KOyhY3TEtwn2lJnLvhRs++R65n
aE6LH0KYKRLmQF73xmMgAidMdNMk1x0S9mNYO3H86v4Y1IKvs8LJm6T0XPwkhEhCl7Iqh5d/6B+f
gXHq9u9RfUKkXydodXUIidJrZ/XIQX7At8OHRN5YKdVuG5T1sIj31Mv2bb4PPIbSS6cxXAbIYWuY
+5zUx6WCmu1ewb4Czu3qILuqcltk5opz4tPmj/SPNoC/lBJZt5XzCk09kwK0pqBTK3SgQQ3/xFdM
ltAPNqUedo4GfznB+NThr3yfgGDpLJ1KN92myluLl+ttsIgkbeK2qSOa6Xe4k8ya2h9QaL4cLdOc
i20ZKXOGdndR6RQloO14v6ewBw4WyKMErHimhc3g7imSNxIr2C9VR+isCb7vO08LnIemO4z0SJH6
eaFM4MEhROpIMfUmwvFNTncB9Fe6JH5+o9I78vSr7HNLPr6ax24mns5tLsbvoFL3EnBZ5m2xPVp7
eHgG+NXKm0tus99nLFg5PUXqzcFbrbGACd6myxoREI352eWdx3DgIeEpp9EuO1YxYjw5xo7evgX6
UUs8CTYTpAKx/ddxole5BfMfO3Gsm7aOS9Crj/Kq82IW7+L/lX7Q1YsiR5il4L3fT7RGpW+yIcqD
j+17FGu0OmFm3fR2IkspiwG7/JckO28RX42iXGfXY+TMYs2ULYBbBPXfQMe3YnZQa5Pf/Cfr04tl
zwNYS2swR9ap32UPVsaoUwfMjwo+efG+BpXoIc0bDUbOiEa8WVCPqbJaTq1eyNg1vFzFTQBgSbHo
uytFsmn/42YCKZS5B8Yx7YSahNquR5KsWRKqVQfyYqBldlGJvYVa8nUW4GGOeYh1jExc/l/C8OYW
A/UUiy5Ul6uiLYlsABPoHDrCh2m7QsutbfSFEsG2cpkmm6jCVnFb3WQevGBOTqbybhkxivsj4tfi
JVn6f2r3bQQ7LLWEGOcrwR6JTdjWmybRm55PXxhQiSaWFVBC9Ud74en+/k7ut/8T0z/p7qeK9Pdn
cXkqWL4OwkeihvaUj3XHmO2i2O+RTeMYrSCTDLVos9FIJRPkd812j0syUG+C0W0joZSWcqxbZXBL
u0OBcU2ep4Dozp41nn0SNBSpAGZXbIBBtwEPLAitIcMbEjv7N2856WqmmefOqyO5Ew4G+5u3ZTqM
mzOsU3ii84KTKAe5nSc37rmshCR+GN7uvaC8nilT0CP1AV9i83hBb6KpfmnAuJhyTz4QiDhrWnJV
rxmadVXjcz4z+Q3DnumYXDRKgj8VB/79qiGDUSu80VS0pxUYugXhu2ZdcvWl7UPxGleAF0bjSWEF
ytsThL30iWJgrluPMYnMCxnsKuuzCBhSEgIWZFUxiBkRAJoojW1bYt43juXJHmiz7swdTwiGqQOg
BkXab/1NNBOTT2jpncZyDo0dBHVI340XE8iZbRF2cW85eDPpinzckEd0b8TqZPYmjmAScOKszVGv
9Y7YG7v0mvLxhEMyA93IFGHLTnzfx/XHnxZ4ejiE5R3isOgcweTMhUHJZOQLN6OryvT81AqTrl/H
lqBsczim/E7Rc2rOEQm8mc4BiimgOGpjlIYlTgWA9wHcRyquETfsKJXu5q61Ava1tzRWmeoBUsxk
E/rOtEtb9sj/Yj42OFgP7GkVb6Na1T62atu6s4oZDApfW8vEf6o4NmNcQexG0sT29eX5MdTmQ0ZT
MDKQhHdjfBNyDaaBi872Flpmiv1Tz6R3eqC+yex6PFC1FnnNOhAUiGbhupUbjy+3jACcJ+JFitoZ
rXSS1kMEakCdY5faC0UDroC/IJEetXZGy6F3dhUv7pAaaPTKQEDs/gji9Ekky8L2C0n8kzaS75ig
m3Umpi8qDWYSwBmieaDjZfWeJUq8/yWgJEqZN5zJ6cbncEGs9HHyyaGA2zv/uCRV5jQN4h4E5dG9
fghNDut1NHFmQGwTXESv56rhuqjmvcmkzWtBg/If/qxzgi6BoAgZzaSA0rF9IpAQlIBk76dHialN
A3544GPXgsKDKFMN/zRs5Avkz7Q3cpAXW2Hy425Ec2Kr6BSMwaLGTDD389KMdvuAyVxxacvGP5CK
WDHBR3jrSM9uuOfClNuWbv4klK7yTWfgBXSYJc8uOQAKG5e0WLQ/x3goNFB2aNNZbHvtekMXPKyY
rkDpUhaFCIUoezRqgysG/NcJ+8+zgILU3N/B8jMui8hBS9x1D54w5U+RCXeBmVv/e0DY/qfQkDSJ
jcbj//zB3Psg1Skf1HfzInKCEwIXJVzDg3qAvQJ9XBTdUJHWyHNwG13NMO0LAgF73XPFSeLwz6hX
ZGaoBrh+JutYK+dq3tx89MHO5O8Ryq9LvxOlYYPcsJroubbnk2Hn388mp23av5QTanhRS7LXANww
6pFcuJIPs4+TRA2nCC8MDpxIEKHbsc+1b4WFUEL1tVOuFkw7YmHsfDwgL5GDp9dQ5VWjNX0B9h+m
A2mqJbWZm6vi7EJbvMyo/76d2WzQeZcr92eX7uLGAWaW+UIH0qjxfcrBf+ruk6Cz0Sg8VlnJffuV
7ixc71PtqL4E2sGyMX9ofTVPZty7UF5LAuefHp32O9ydRCag1aIP2qMmsSllqiLWrApsixwtchT+
3oH6I74Qtld04sja5JFixTyNp1EdEO9B61dLGjmD6PC+tZWbKkW2TamB+zF2L1mPmmc1b4QuZ/Ri
9fq8ztHUExaee3pwqM1tCK5WkjUOVI+OapupfYatmLp7ZO4isN5+SguceQmBW7kCjYIxQ/YnIOYU
aaxUeg2VHlEo50KzW20/LqVFcruY5BZ8fqH2smw8v3skvAuqAQdZNNbhwVrTAC5wertWEYENcYfo
KRlWXVkfXCqONMqQrWrikAJk+yyrICtW15IsHaguNQmKJVtwAqxTmdrbEWyNrLlkJS3Ung0D5o7y
2Wvl7FCSPxnyGTBufcZukgjBcUeJC3gYLpbl8htxUOUjrC9GSNYBtaT7fR3seDmI3EBsNruar/Dx
ZeaDnkFwcFyH8wEcWYPwLiZc+Rx3YJP3f7S4hn6l8NLeu7FVJqyd2FlmJ4SgqBChNSS/JX9FFeYp
qNlKGOby+tlmfkEmbAfrJZP2HMliRT+eRFz9f6NNYIrTa6Caln/KhCj8LWGVJRBEvnBXfjjPzyE1
+s7sCnSZPo08PRgdZHBjx5RzKuzMUAcRwjhM6kAJUfHauS7re7nxHFWOWNnfTcQ6i8OGQKM4x/BZ
0aBIZRr8PolY4pmYI9QaghUfZQ70FL25PT21Xy3PA78lijOpC2zNtIW5iJBUiIIyAucUNLWwmNRs
Wsfxz86oJFqyjT/hUWLNOPWJw8Ppy+fz9An5OCkc0hiXFXbsa6kDF17KFdMTbup3ikCBY3LhJvEo
jXbMD1wD2c4qYPmKZgP/yQPm43oQ366/NxsL1UyPG7q5JXzpWHGNc6R6yuVK4HUNej/JwHSjHqdj
8a9Psctc2rw91BmUCUcp2z8dvGh3uFXbBmUG84aVR91iOZ9NcgaIvmxUDAFeoVkMxP0OIhF7RZTn
4O36BSd7clPPgQALBqtmkKOCXiadrFLAfEQW4kqvvZ9qOgR9gzkLksH3El/g8NiKBzqTNkmLPejb
BMvYCk9SVwGJfNezyRalefgcgunFHGlyMbuANeUc/4LJ/GvCjn3Z7KngPKgCoRe1SHW373eIqc72
eONQ1tofboF2L2ai461ukDU5Xk95Kr/8Lac2bs1MfYJz90Eybow16EbStUBKhYxgjRjyzmr8C4KL
JXqP+i19QB0uwPoZCidJ0Q3M6ucHC9c2xeH1iHNMqxVsivngcF0wTwQzHHvsyUzleozRUcfNprYF
UsQ72k1bTyDBgokWQ5Pmn8jL1WGcTmBN/RAbKFQxz/Z8Y0MUb0UxY81mshScA+KVM69aZcX1+Rrl
5Ba3QZt7Mg09SHc0kcAaMuQ90B24tzZgGF5w2S+kzsiQNOvoUCZAgP5XjloCNwAKREHaA4XIALE4
B1eh6nFBzT6Y8zeASfipjPfs34ITCNPEDx9iyOOoWC8jqD4qgOubvTVHw/cbvUGe71JAKivchqb4
/zZp+By6K9Z3rw6K/uqmIhNaRzBkY+jwPawpmVkuh8RTh2yKh7CDwKQ9uNb2UoOeP1MVhbxcUIGd
OkQCvgVbTMRYTrxksx0mAoumVPOfMITMu5DFK9gkGQDW2YNBXBWxqh6SKNjbQVi87qWPdLZY+V0e
BktMBQL17KprHqXgNrwsJHhJQD9hChyju6TAH8bH8rHGxCZRk+TClnQYD3hzIZW+FjGvrC05pTCS
xYEtqrzRN0Ty+ryFu7qiSbGq4qtxJlEBeMvvM5bkiB5nYuVo+Zu87+sP75gwpDptJ05xs61GZ5Ef
fG/V1//j6uxW++4c+/Jl2EvunAGdRjEihUeDnVIbNopqhO4s+FpSu0TfyrmrN74bZspUvZ3JsaQE
RsELXV7HQgJdI3qA+2YYOdc9hQjP8X/bHQBQP0FzwlrI+cUGquTzwQ0CPs+4hKV3B/vzkAWWnl7Q
6WJqPomSLUch54jbNOFlOwbCvQSU/CG5EWrV8jSRC7d3i9AS+DWBkOGL+0HV98YWFFDL6mWnvwiw
smUzguNMuHZ8GzrT+/vl68lmJSS1US5mgvSmHePP8XG6gWiZAqXtkYuMJ33KQSxEKsdFerofiVyo
vn9Sv5cutAKdfr7cB0Be4suYD2RO4606XIbx3R4E/pH+2+xYdv0zh6tp5J328YAgchSJ9U88vf0r
pJz5/eKWhTRzES5bfmj2tABAm4+QUi7IDWcuMoSHrY4BggLqg4ZuBWD96BY+sr79yMRq8mo3erYg
XmVdFhgSOfjhM3/0feUbCkVS7bXuJZ4dLhjirMaO5zFELHJaeON3s7TUwBRbgwYNX2384tqhcqag
BMAGs1/5yFGsiey3rSvJ3LHXp5CqW+1aqweid25g0LMk0c4V7lp9MBzJ/EdbYZc9tqDIPGgd6MRq
/TzdNUs40li94JDfRTejzqIP/qiVZnap3jJfN7vmQ6nF9oaKlAVMS4IQoWgzRK1KfiDmI2stxlZE
fUhITXHY818E3uRf8AsvXncNQxE5jXQ7FB4DPw4UA5RPMJXoON/CGizhNt/38AJaacSs0WtQJFVy
yQJlsjbIqIKiZuyEEWVb1F0c4lYti5IXEfeM1CqWF/ua5LTEbVVMxYIWVEe500QkMDkgwzNvrRoh
L6t9ea8YgOommbogexu/4a73XJ4l5v+DgyjcBntsy8Fd2oZDSaIvoFDvoJYR++Muyvwh8pzWXbEQ
itxeJ8RgTZOOJhsgvM5Ab3H2ey0YgeMlHhTV00+JfA2fcOIQECaadKBxw9XPo6J4up2LsfwESmol
37DVSHLwVy/NStuJEMR35V3bVpUZfpw7OTyJRkMDq7KynjqnQG1HMmkJuIQOdPq5sDbYVruk3yui
U6LQY0jvbgAH4O/LDlVhdDT9TgoL68vaEUd7ipCdQ0yhPtjhUjfM1GHq+S6j2/1l6zF/lFWRxgG/
59wOUwZdoApRbfJQ//pbUu0f7DqQUH9rAYdPSdcUSduN3UliVFAK5xzf0i0adjhhIIaTpGg6qyuR
8ALQLeqxTnLWStnhmS3VHmLqeyncBWqjEBLT6FrMz7aEPIvK1aGbMiA3t1TYDi+PUz/z9dGp692K
YnVenX9iaGhZ2rJgPM2zTHP6ZjxUVBXDyW7dCxYT/f7ChhxHqq+JoaGWXRBSyNt861tR9OOhju74
B/j2DfrNNyRNR/ZI2zpWOZaeYnB0GUwPWn6YIWhPE0jHntay+2ciiqLmhLCb/G9sKqZcXslK3NsN
ljo/oKgPnixcrwg9jUcLWJv5owgrobRO80QgkigBedb2yjZCKIhrxEuK/UdR5MMtiuo5fAP7Me+c
D7FFqqXGwNCnuS711wC/BEVvT9uFKYhH0E4miDYpUz5iV+Nz+nKR4Bu9+6Ey7DLPq4bZdFVU5NJk
GK3pFucNrFmcpM2bXHCdxcm/fBvKIYk+Xul9HabNwYUi3jdfkWTbMHVlZcxSADNzLfvcDq4SC1lx
n3/oJnG0qYzc6J2jSxwLVjmC0FCJ2hSgSFg70thjRYVNZbc98dDPrVoOd27Ro0MPO2b3aV2RC6ZO
XxieFZbZ3QKHi0n4ltg0CCQ/BQ5kSH83qqWmiIBnVWsXSOAs3mEo6D9LBrsLBKOYt1+xMGTm9npk
NxMyIOkuPgfFHRB0uMSN2KqgFMxO36HwHMVmmdWftt7JBRecDrCHK1CphmV1hM3F/V70AYJI82bo
U3fQdJKz/HFdIA5qIWsz+giH62dhbTBV5hBlSCUhkovOyMb/U5f8J/me33yuUfy97i9tncfcPXs9
YDealQWxuHtXkCZ5/swDj8iofUUuEJA+75kwDwi1yc/K1QdIcjR9yKAjnw0ZjVlzcexd74quTDsu
whutEkjY5R54zGqdlSIVC1CRqZ618yoxJBLw/CvxxAq5cCeafSHfqQ/KSEz2aFcEAQRPpw/OI44u
pBEHfyK/qQxba75dhyt5rN8PkiTPKp3mB9WokECvIhFRezKx/XZpIxIHcTkfFgdUrg3gNDd16qrL
fMsvOTpHZTskKg5oGRaZtOWHFQMX0QJOP9hM8axOrfd/fw62+Ts99DhD+PliLo2Ysmkh6mnDgW/c
EKAiPicbz291RjIy79A5skqTZ5bBZ41Jh1mJ7eZhVdkyIT/7ts3QmW0ju9HLGm5bBt9eM9uMf+xU
QK65d9Fi7QfSdom9C/r7rTXW6HZxU7+c8Z5ZvbsIglyQU2NVdzYkbKUKADKcjROF4UxgnIMn1jSI
8vJW4yrmlma+xLihrQnxCbtyTJWg3WhLCEn2VWKhWjaqCxBjy/BEWKrtTQPkBWakrdWoNwTH6p6N
kn1Q8MCGPdEP5DcJzPe5zQnlkR1lYpAW7affySCTynCGhHoFGV89SklYwMFtRy5cw/c1+/LVPxWv
jOrwLpoMBbPCoFITK3v1cM55RMZvm9Q3d9yVMLMEh7H7aXQ+J1TfuUC/qE5mPdutiPxjIKuGpe+d
b7zaLp9Gd1RlGNlH1WQtaezd8geh51Kt+9IEqXykMOXQAa20fTmm+L41i2xgRwynp0EQAqPIA0PV
ybVJvWyTSF685KUuOEq27YhKjB6sQvSWwNUOHc1LPTFVUehEfDRnnf5lCrtLu4dG1LXtovXWkJkK
UKANv5NDysgqBaKXzc3hA5J2Iz2lj2b0adJKPQfMtJrHm3BvOYp0UdO2WXwbVLwqMojBO3vntE1t
3kv4mxYXDZJfODAxklObzIER6+oMmVpg5XCKqaIBJKNKye6ntJMASCEt8s2G8d7lDhHg3FyYFmav
I/+dEaEalPlHWahUzKFHokZF9QHrzLgL3in7sH/OIocbJls/teqZy+lTyf+CDFpeJOMcfmLI/cwY
mN17UfWkvoPA9RXoNrcOFmkIpy8meKXwbOTs5SSSWhxkvHd9RaqhID8EhW91oAyf/WuvUMkW3FtV
ntZ610Viczu+HlPB1oP4dih0dbDwlvApGz4MkCEm4g+7NXZAlc3I7yxg8cGjDctju+w3lBUpAaxp
vaIVBv67q+j38T2p86XqJj+x9Q4i0ru/7+dio252SSfXdv+FSeEMJ28Eii3ZVe465WGTkGatWbt1
uqYOH9d5nwgbJZWzodnKRFSjm3VHItUV/qDWWFZ2PAXGNxhmhfrDKh0R3zjyluwZbsVnpJJ8rXcC
gZtFkzgpmqiYdKeN+I7EGa5AqVjAgHY9abePUzWY0ZPm1Mc4dq46L1xBlKl/Sh4f2nHCZehSrNXE
8wYRLo8KMtRhXhbYApXeVApOjJb90+qpPIGq642fxPMBogMSguZYwpRMsJwxl0ZQ5VgajG5Icx2O
tSNEGCQ7EWRzP4xOpvsbb6bYBRpmmbdkJK7MOhfVF0NUvRUer5NBXCigSmxrku1Md4BmGy0axr8D
N6AOjiz+gHY9Q7v/gBvYKkHd+TxJwNnzX1/J6sQZ0/f96L08TBcW2go6sREeyGzs7e4R59D2K0Gw
pju9MeMhCV68KDspScb1s2Ul0HiWwJ476I9Vfb0aYUeWrsrO+ODzPTHscY3W91+v6vpESv23L7ge
yJjseW2IH4yRYj6vOnw7bZQ0WAaZPWCXXBj3s8w5QDw+b4ZDDkXDHPWXnylrIgDpzqkPUj02RZbP
6Ih0miqI/oXBVkS+F1m3Y2ykPoLxQSywBFevQ3VbsdnHjuFG4VOWKVZtfcqTaPKWkiukU55fzAxc
/L+h2ZNWuUnpx9tyeNh3jadPmTT/HCrqvxAWaCTgv8GkmqFSsaBZyc0gQESVrRD8CprLLICr2oHk
7fFoyXXJmMyXOdhMSZdea+qx8/gjhO9jSfMuitR/mywx/Lh2joTZzqW3Jm4j5H1ez6/ET2u/MADm
8p0kXKcMKzHNUJW5IGG+6zCK0O7Dli0IshPsLdUgEUYos/6WQ72XMxVAVZHBwaRNGUgdNkIt/ADT
BkT8/vMhwW4mDE9z8YwASEIM+nVp0pcW0jXAO0mZpv5qI/UdSwma6i3rTY+6iw7xwcTDdAq3S/om
VLTXj1L8P+Wo0O8+np8QC6kzapEsazrRUGpg7lsaZ5s1UI6W66MQIGihv35SBXkc07CBXXLT5jv8
g0Qyaof8+OJk4Qs8w90nuH7sVtjxQa/ZdeDW0F7pwS6JOFSmO7ock1I16IL58H2eF2a5Clj875ln
XJzXY7tHIN9h6caWAs5JScKj72cCnCzRRaRoRg0TjXUbkZmxGqVdBvWIDSGlhrNnkFbadBZOMAok
x2mxDYEm/1CfLZas9zobgZHTiSMQrM44Uy9+3Yb72eJ7lTBtguhpJy30zVvAxTcKc5VlmhmquSg6
d2QG/8LtJEDHr5AdhWJQVS0k+kRgVz4CBMCwwHPO8bNUTb4RFU9ZsLIrKitYMRgk81VAPhMxh51g
hQqDAglMdf9oYMkZ+24KBKYlpskdoTa9nOX2RZ+3Fd504yi3QFQGDkUGIZskZdgcsKY4STQloS1i
jYJx/42/QIOUpWS9quQYEG9X546xF71C+mWLXVYN4scWo3W/d5HYjU027R2QQcDRqxynthcIa8zt
sE7oY/hLrlzZPbQ66j0ffUE46/WPicBZxh02RlOwwRbl2reliDIEr2L7aZXN7Uq9PY4FQgtKcBGo
HyzkjG+Uyb0ZBHu+EcYgjAjyXmd9h7VMjIO33AgQd8TFVnrSVGNXYlnYs99X9X2yZfVd0C89tRqC
jbm6gEBZdO8slYh85qja/YP8EbKFDwEp80JTVr+q5yMYRVjhnR3ev6qjpiREiEIYpB70pSIYv7vk
rymqVBFZ0/kZkqnZYqWUIgFkkCdAU6ZEl9NewElcQmmXy51gMHxRnMsDiRMaMhACdSir7Gieg9Kj
rlGNwB5QzA0XJ2zWSj1un85CsSHCdOVPy8Km3/yaq61c4Mjawfzgpe+jCh9fjk5g+m5LNLQglqL1
Isz5niUxWqlfu8izv5I4eBCdC7r7ADYTSL4tuQU8zIzYKb9RHJVZ3w8sA/yayzcCwdckz7oak8NP
F6A6cN2LjiHYTiPMVH7wEyYKz/bzGfynyN2fNOCJfuyQewVXyf3uODBpAviK1wI91W3230hWpnR/
YBBnlQQCruA9UljeqVU3uQ1zg1rSx6ULyXyYhH6kqeWT7BZZg25bXVItH7/44r0k4QtKAxO4DSI3
7osikm6+3Kc2e5YpVUexWcs4cKq3rRjoZWF4XAbMb3xmfJkvCm0vzKvH6ViHUSgBV0zfydR2bDdZ
J0vvAummFbF1nAUUXfNLQQzhHtXnRSNAs/K1ZEWDKZfsJ4jF5UPBXkUPahGOnNrNiTrQUbKfA5NM
NPX8tBuRi4oTf7ez/j5MnAFt7sTdlgealTpoO27K+SdsETM2HZKE+EQiDKJB31LTIB6FepFhZ0TQ
WMtdr2B31YJGuwgG106pX9sxxfNs/WaQkm1Va9bE6XNBBBXk6ppakkkcTYleFZ3ngQ8JQAaCowfp
DH+hJT0jGcRBTxFkNFhYyQvfT6Y1yc2X+EYI8jsjSezkLCTG2j/Oa1zigYA2a6MQx59Rjr6IdqcW
LyeQr6fzETfm3T9LseOYkptkxt1+OIJXMCAfYlm90Qnc6STfvHYGIJ/FC3YmXcnssAx0AAJJbVlf
rGO2vfWgZd42c1t+dvKv6DPy7c2gzBVIjAKcjq5pkBg4AH/2I6fAWN+xAQ1pL3qbMKnVf0e+mu/1
Qmgrf7iVrszdMKWt2o0cq2uvkrw2lsHpVBCfn/sVIhjX4ebDw5fFgkH9wT3f3V5idiUHwbCJLTdy
kf3snN5kQ2TzUaeWmJQfFp3v9zc1kuqe2BXzT7omVZWL5MmqGiW6yMZe68Lpp2bKakI8t2RT2u+f
tNgNqYAfHaIzAPhys9PnOeOo3H9B3ecvpYhsh6eTtT277fyvBlbFJRjbJN46eanSttae6t/oog4M
rdC1vdTzqIhC/c/CtEJ1JkxZbmQtbfq9gXQQujc7LW34uDeA6F/gt4DM731o2vdLsp8roZVD8WFM
+MLR9JnjEhE5F8H09l4Vg3bwpsvXjq9fmDASUb6ICQkeRVGiWLceR+S/ET3pp9hE874GcQTFTbLK
s0hb2XIzxqgXZVTqmruG0SrLGrjKlIoEH+kmwo7HlPa1SZU9Hu68vJPRGjlBMiog6M4oE/YtG1VW
AQ3qkEo+Ox6aw/+/LT0Yd9JrKR4kP/q7BElF1x2WiW1ubg+KDVwMbzkkVd90/VfW7NdsB+62q5uy
/YJ1UL+Sq17OSb7siVSzJeXXWeRiXhHDPXIN66sOpbkoBCNCF8fHcGMkOmRCMf7B+7EK4B12+Tn6
T3mUw+mOeFp+/we66yFm85XFB8j+5sOvDYByncMN2J8AA+cei9rSXdOeEEoGUhqQ8HskldPllhJI
cPJCUpW7xt6UiR6uzR/F/LhMyUHWTl3yEg4xf9L/ujXrsFmZP5JqfLSy0nfYphZwHiWXadVSVRNr
tUSb6vyDD33bc1EFM/32h7+pIC2Afpu1EpVzyUL2msIwogu8mqXg1BsZ+JJ/jV6vzllDy1JjBNRP
U4VpA4z5Rs+xWo/nsWmSTpc4h6EZps/R4JsRTcwGDWigBQBBK7WrlXlbxIkyGg4ieNVFTWGXRzhE
5CIBBbpoTgTpQKSs5mtnvn2ESer6OFzJjjFEqxZvW5IhmjRj0hs93/hoTZUQ3n1AGXq9vbSlHkgw
kDVYV86l/ma3wkcCyZUAv8uj2WGGqE7TagrGUt3oLJerBdEkq6Sv/WzVCvpmkVhI5tE87x1CwWoC
nhVVdlTNoO7w3502/66r5bvc0MG10UJoRvaRRS+VFBClaWDxq6+nPO/A3ptBHh9dZKQhHCg6GcVo
zJRJi8lHPUTaekSBEv+dKM1OEDhChZ612BxT3nTy8YPObq/iE1e3TVJFVXQs/SLJfSRwPfrZ1X7m
8U/O1rvQOSMyRfS40i0SwjdZEZO9epCaLDdAztdiO0CLU9VgxYMwYZGsQVci6lKVDSXzkn3DicIu
VYXpRAyJ560lCw/oC3Csi4OWBR08xMLtHO5R05zamQIx1jwYNYwOG5/RnRsGwqFtRytvictdvp3q
9Hg2kIDvrvAL2IUFfqv4UpaZ5WPWSxLnSmcvdd8MMRT36Ezw7tQ3ZcAwUbfIlSs4vgMHufWx/0j4
MnV8Lgq9BhvEiZy97w9wyTKGDnkY7iugk6rHFyHf8t9V0a1vRQyjwVYoeZuCVxsQDMbs3wzzC2Su
LLMWE1WFBovoXWqNvayjvHAD6mfYtvTqlK5+3S6sS6zEwsLCgXg/KHkDt/jXpJs/vT0XOBgi1lz1
km6H9NWxsKdH/a866vYRdb0SboRf7QdBJpxIvq7Ui0461kL8+P5zqUvsHqsTwm4c05WP1XDSv2uu
XJ77Oyrq2hPVvZ2Wj9PXU2f5os/Ky4H9X9MM7mr59v1ogl046LLyTBc5yhSaWRaHow91Lpkh7/KR
pzLYaouUjNuenIP7ZIc6Xx7vaR3X6zICZyBcFx1aR5f0oUoy5c1GTxocXzTX7Hmsn2bbkSHHDV/S
OgYxOXAlaZVVChqGPhJaoswOMXAnB7krYgBj23Mrnp/zhmYlx5EmpuOBjcsCvinl8gjVno0bqrnH
q8UZLuKcgQgYgM6tpNi+UZil8zAEaoIRJc/x6/DtMLDAzZEj11CNfBTpNHxya48jBhlOFfDUTuoy
YDIMenYPEIVLHfanJDshmWRub+PC5VxqBXsHhfr8OiCdrQb4Tw3LivvOmN9a7zWGCfvMsUaSudem
0Kp47LCkZ+HKuD9aCnqGxW3DPQCRpW4BboW1MAHrnMGtWGXTojQY7XK87Npp71sSz11VPCfP29DY
cV3F/HA7Egp0H/3yZjOylRmUt7XQ/gvR4Db2i64H/R3KEws7uMtpggyLc/ZuclRS5tIfZ3g4FctZ
NE/DIZA2MsOgZZdqw6LV6iwKdR5HSXQmFBmCe2VxCo+n8V8IW3Yc6S6+TCariiPnkJrjJBouaY+1
TUEtSYrvQjZporD25yLSfpYRFaKxlNkmZfXkkJbOJk22Xn/BZFUKjX/1tecofK30aS2SDg0V4XTf
JKUT7zT5cQLXplqSEp+S6RpJSzQznlzpIL3VcNeGEHqzk8wEN3+sgSJ2tjh5DP6w7AEPjj91tZCE
hCtc23OG1o6toFYFjv9Fznce/GZ8MXbJykB9vvMEGLCb8Zz1xkrQrp168VRDVLOm0IMNWAeTiIII
w+c5eYw5t1F2Gnu3bGDnI20mU093VZOlS522lNzeI5bvbf+rs5RdiM1XPebBO6LGIN0j+boz9Xpa
E0zFc6EwaqsulrN6dlVT/OZncJVq/qpKB0tvzDNCO23y5EqxzNluGp8jjODf+nF37Jg0dmnd8Dco
BLXs1Hg0sqJo7AGYDSQEV69hzbXoO0FnibvBcDPwEM24x1+ftIHCOZ3HgwCp1BIytw4fMrNF/O9b
oHYn49YgE3uHa7ke/IA7BCIKb04yZMal+lkZyx6WP8AEh8T5ImaVEInkZDbk61Yu242/Z9kMeOpD
tB7PdIjS6D4ImjjUWDBeBb/GQsJKWsjyFKiet4SprBcFDctFwDSKsRFRPAXXBqfP6pgN0JCpDrL0
b6P79D9x0ovLP18IvHZyf/xM3nhiPNWwZjNdaCE2pVWAni7UeVrHYcSM9ypZV6e9r4HXS4aIu/Uv
JArcWQm+g2Gf2KUIkpBUMhZO8223RcUY59LXYj2DCA8FOWKTvu1oGwV/kEYTXexro1K7wm8jSXlu
x5AdM59Jx1ELjNc6xV8RO0Mg4ccMSAq3+fNWjQZPbu0uEx7JzbRmY56mf6uK9qEgd0V8KGyXoPZR
nuo1k9fEqCML7LTAsLGp+3vFNgwsnwOO8vtqvFJwi0VjaNtWpKSiaY7Oof/d1q9STtZTFQ3weKMN
Y60bpMnDMIZnqvqYnttqgkUr58QS/ufKgHa9PevprrZ0oF6pZ0bEdu5e7kPkrWl3O/O/W/wAs9Gm
8Nwp6laEQruhlpqSDm/YJfR89jhBGOrmTuM31pBstvBmtzJtJ76HNjAEwUwqgrwbBCvWd+yRh2Qm
HUNVkRRw7t9MpcPCBEm45BDIUStug5vw8S/ZtXmzTwGAFp97MKs8txZTypnTKGDht9qV4SCUGoTq
fwRrO9iV8p/8VoDoHuRtwIvetiluZCkCk5WUpB1T/f8JmAfmsQfaPqgG0fNRx4eL79J4g0XZqTUq
9YHQf2i+Uj8YJo6rCs9xhskVJBDWyMCH4TMivciCTB3INy9UDwoDCMUcU0HQrRF06xJBivdtNvxb
Aq57MFd/bYoinHTqf7LG41DQYflxMRbA5o9vofGacZFNGRtXO4Wy0BBPnvmK/UwkZqHDe+Nfzkwm
s6EuPEekwcSQzAsZ0XiAwjOruNUCREGf7Tjefc0TSUqlEebZnDj9MIhVJMDWvtUYF1d3xq7Lty1f
xumWTt9WMPgd8+ZOa8JUjxuP3xk4h/IP7Uji7UAYAbn/DNr16tl2Vel1s3T7GbEsQvFaoXO2w4NZ
N9PdvYjsYQcFUvG0jvStpIF+P0xMhXLpvdG+CkdgwFoOEcanPJq4Ydkv2YAoAVSMO/rqfQGAhcVm
rWfGmGGFQUIQfD0XcGOnYY4K5NWQQ58fG2n6WujBgCbTJSRwJOb4ywqx+0bwvJo+jCI4jb7Y20Sy
XmYLschchQMMaKe/NnqlHJYaU27cpNIDV7VJmNQU9CeIjPvdMJKNm+Ty302c+A7DM3ZoMmCwlwQ0
nugU98Qa7EYay5MaQY/TQhhupOFavIXSyxrHfwoRknQUXeFk3IPoiGB5EXth+f9fbvgWBXr9BDXO
CgpBvUedskRqjwXxz2/FpETkd+Zp5GaMN7PYCghf9GBDsbF1G6USbBCyyW+mELgiplZrOVZ87HpO
xw6HNNFZcYxjDsGVkysel10TeS1VxAgaXbPraJ4kFh73KYBn76c/xdYoRpBr3hCZIc7W9A6pLJfK
qWTOf1TIaa9Wjv++NNWjTK83H0Q2M4bJ3TfOxhdlaIM/ZhrZ9/P1Y1SjCV9eDM8KujrMjaX4y2jY
IMjFiRU+8dVpbVjoOrF5l7AqfYeqFP+LtabT/iJW8Q2jP92sV3atGC7BRELYUXC3glFHU0sPumMb
ZI0khbaMh7Om1t8GbXNkKW7JFaZIIGBouFRIl058LUVqQ5aUB8HJ5aSu8Lej7GyMMT47ulO26243
dr9MHw2koWWBe1bNUir6JuaV7ZVOGDdk2prF29uyQNR7F3EriNGAo37HWpKBGrALDzKhMEvhqW2X
gWXzpWbdca/2R5dvjO0m8TJqi/vQrtAZ6ss1eZXO589cmwF+2iM4l0lDUanmoAVUKeL1GlbfJJow
ipg7PpZgEvWUoPOboNZJWtIM5+gKi0ukCKr8W2ENYoRVyUTxtciFHY9J6LUohTZlMIVRDUhGU4/n
vbakKLFa6ztdjI4/0AHRXMxJjHeqYt7IerA/vPGKLmwiK9urM/TQmDpCBu60qKFmHwUoxcpPrZ3I
ZJ+fH27cXSnTyDLTiqY+tRVkQsEqyhBvkRSAuj6Pd3/Lq+et6UcbFPFjVRtoMvpojiuBVz+wbxru
fR0Nh1LzlFcot+HCzhiHqhVApRbE5QUO0ykFsmpuDBPPDFDQ/vq5bqPU7pYE0aKWgnkREtJhM8Z9
L4wPKOO7q+VGIQzm6XhQulKJr0lNhaU/RuxWsO0rBQEe8cutHoEVk7QYB6ta73VB/usUruyP2BZk
ZDdRmWfUVCtjig4GZ3jGhqGh663rSj0p9O18GvYolL5AN3IBN96LJ8MmmBR0GoqyDoL3gL4jHB1o
WwSh9TRmjYpxjjuJJxvhawh4pm0DZIVbjChvl9SalTOiSMtXlj2ouGOQ3FYjnvdWtft8/QZfuyQG
XXGxhRKg9/paqlyZmbV4SLapB0Ogw3NnvnzDqiYqxHU7t8JPjIqs3xrZbTe1Qvp7hfD0j2jvGGmk
UAus1r9nAdqldDFr3lYr3NVhyA7GhVevrtSpCufPFiRp611gzFfInIpH4rJujl9VKn6aF4KIiECj
Qo79XyoJBdmSPwHJ1q89DyHCAl5F1To6grSDu4wgwFMiWQmiPiOGYPqtvuSYnpgdKV8u2vTD0nlx
fIYmHXBiQK4isqtGfU3437ZTBfQRuegCandPBPU/YOBVE4lsttjzmdTS3ULIupBmEoTZkJdJac8d
WHhr7Vx2siwftv6ftMmIojD5w2p6zl7N05K6nfc5PBEVPYFgUJgoLWPaEebJudXdd1wu1JOWz31h
Hypg+zfWCBqioxthk2wHPC1fgpPeP/hh4gAsUL8xISIASb0n/Rxp/Wdt7gjl/MXYBtYK72qLagV+
ulqAODOEWsIUF+yC6sHkDyCMv8ObHwd1fp/mnxcJh78bz7UvUuOvEiqIBZu85hoMduNvA8c5gWLj
ov0CqgzwaPjKhO97uxFFxFmDQnxYgjj3z4w8J1+9Y+tp3e/hMHBDvqiKQWCzziSFeNSKPMCLGdOt
ELG3uyBm2ooIzf/Ek1yk/5qmVxa4oGhl8GcGLseynePx8sL2GD0xN5OrOjL97tGFHH8rOYC2MxoO
xy8wPukSDrLw4JzrUo8kR8fDlCYtNUJectZdos8oGzUP9EnJ3Q+Zm/c6iRDt8n8mLfA1idGjdUIe
93LkPUP5rFdM14iR28Q53obT0IlvgwkQ9CpjCTg4tvhSR3VuAsQPABF8NfhQlm52aawPRbmWY/Mb
V+7iL030sQwQLMZW7q7Tg7InLQqG6/FuXwx6N05aW7p4phIRpU/gHgQqFGO02j0N6KlhrtXWgY3k
JGYQix69UtpE860h4E0F08h5rcDhaZun9qn2twM/C+4CaeUEN5w7flFHtLtjiWMH3JI+8W4SGBfS
YbhB3VjHQKbhppBOY7GV8cwgkf4NIxZ03VPuLtBZ9KYUywx+FBRn3wW+xpok1bIg8yltnTs5l/VP
k6SFUs8dM5Q00b+5F5LJ+biN9UUBA75VuQkIHlYa+mwl46A1hUwcG7xhccCv0tBRff3LMg3H6/jK
RRZ/vkAIOUpZpJJLilJSWLOGt3/74kyuZJ2K0RSlCo/iEDMbLEh2q6JTp0tFs5npIXGkCX0ETfca
FET2u1frTG/F0aT41cdLEs6mbBXo1iFU5d5o1fCt7mg2pE4GRd6O74X9oRiu4XiS0r5NLqxc7/O6
8XWJp7Bpac40Bfhjp39jHOZhp0JxAo8ZSpgXRWMUXLq7G/ncs9OGhFVZkA+/eEye8Yg3bfItJvw1
2Vy3aGcnht/+TP5YokwFHUVgC7HUJvgkgd33zDwP2+c9LRH8LZLHfuRzhGHHbpzU0v6VxRwZWpYM
aC1i4bUGARrPCkUkISdxGfqOOhqKnHwwmyCEJmRj1qP0Kk1DqguHyjFrXAM3m89LWm2GKjqH+8X8
PrzHOLJ8ojlJGHMhpiZs+h3MOWVYoBu09pielsBH7ecYUwWYguKHcCcSN4zST6KnkT+oPoA0pfZJ
uKoeiTydRfPIzBLwlb75l8LTx7RJHxO6ymNA5udoTOniIsqi5mJNgin5OFlHqxuDkTEIn13u58ER
BBw38EcgLDavOlcvFB+kVEiK3R+gARU17cV5Fw5+fkcULDOBnrh+QYLLI8mIASZ2B7e0NXJUuJT9
/BfOtvjPOoNqUBYhiezVR7g2xrMkNTeusjrI/eksRRe4uuXjvpMbkf9njfR7+wgON43PAHh6/+Rt
9RIqaozZ8BygLjr2xaWhHxqPSlnqh7wPnhSkVCsa7a3HGrc3gwRPvJ1WsOziOBgoap/68Y/8T+Sp
5jrYUoXFz8jIG4rbdPSKpOkqv4BnbHMfaAe7/Gssk+77Vm66bYX7zfs/NkWEybFs0N8ox6rKcIWf
T7wx7+9mMN0dpcZD7iji7K7z7xNT3kipSYW8Ese1Jhy7CPs4bgOJACdBzJTqsIS4B6AqrbeSzPvy
tWDyr/B7R3VsYocaO9soWgHSaO13+mj0fqmG/N7/Ls3MUKujIGskaKnBgVlyeGBTe6Aq5d8rm9Ts
+cjDKDghBjeOKwNxFz3e51E9s9tJLldstaGqefUIBl7P0ELn8aJIr9Y/IT8Be0XwYIDfqIFqQNTk
wg7tN5ndAeTPkYyxHAy5OlwvcsR7E6KfC+1bJPg1lEioyZpWmaTl0vcBRrQI8edgs5+wQX73sG98
R4QC2WiAEOHVLDYf02fmvd4NG6E9Z1HsplE4RenSo+KLD6nV50Qqu9Dha+Un/AEGIPT4R/jaqs8J
pVGaLoZvrkqOTd4ZfrdDTWqBLnqKk8S7nC6DDIAZiIansE6czBdi3WbvAc5H3v9w4yveifhKXzaq
AQMX6KoPMSj8HPZPr3KdeQcLmOyXlxFgS7gk9NyZ3mfqw2sfDWZ2OKZpom1WvHH/sd9biA2qO6rg
VkTjW67UjuuDuzcjRTay00p8v9XhXcQ7pusqCEgvzkQedGSsnqOQqUsBnadSpACV/51ErGO9Wr+A
aDnObp+MpZEenE5mzOysTdvFfoKUzrW/wXtd8NNYLwJ4zrnepHWKH4v10ZzAvZiVUTFIefUKqoHW
FLS5luqgAlZ5/nMrxOY0zWwXui6qjGGZwOk3LwoBr5F6EWvvQz7JLMlTwrZAq56BIU6o5HgLUZuC
3uraYncZ6SwBLymNmn20v9iZ7nZC9Q+gL2VpYSHOr2xX+Cuc5DgFURFfc7nyGUwGMIAlfB9sojls
vsUdS54acyTeIXhgIY1A5E99G8m9pWcK2f2vSjjCDSdqK9ubNDYMiS2rVGfVxmQORhf65G5LnVUQ
Tw4zrYAhK1yw/UlFPan1xBIWVnRLg8JafikrKJMskVbc50hV63/VanDXTBajqrrZ/pkLF8AQfGTT
Uqq0quDyT0O8d+rRsNGI08+Hf5hJvhOyUtLQ7dLCulLCdeb4dQHH7tusJlZucZr5+O3n1Qv4V6Xx
juv+aPg9F1tLPIvLYqCRibTQFWsMwlGAhBGDgMgBuE6h1HY63fRH2AGo5Tt06yLeWZpQ0WvyuRRa
/WzIhYFRLGJxcDcYsrPdGdesTZqGwPO4agOL0yUPvtoNT/DeklFBAtWp9k4pcNCDsrnfP8JEcGOE
82JHekRODLWELsp7byispWOYOpfJOJw5+sN/j7gafVncQzx4xDJfPn00jZmmsmspwIiRJAaFgav0
WHXJMBaqQX38MnlaulWLA7bgnVIfZAAlwlXltYB7WE7dzFR81u73BCJVKrByFkIrIrvO88xcVSPR
RIjGcmTxLPb05a0IW6Xd/PwqptUKuRrtILZSEmJE9xjEh3Q6Ca4qdB3f0dJVDDjhxK5OzmfW6vNf
xK4Sf3Wj/6Z1G6wiEZGd8DhkVmA5Rqdg1rx31KloZzZbNgOKwHYih/nXRhJkf54YCnMIbuvzDGGN
+qBOaRttjRiWFHO0IshjcKZNvBIhoIQls0KttG6o4v/wiWqolFM6MLtG/jBqyfq7q/SW13bqLsVm
N5aBD21m8Bw/5bSkMTvOABcXRptl5ETyGrrqtwg+uAnU+e2LSbSusXg5EyIbx1U97ACOzPk4oC6O
cu2a7vXQt3lLGzv/Ca/MrDHf4BHljmtXZc1DoWG4CLUuUI9OJJV3RLw+b7GzjmgbO0Q45Z0rK9bW
UM8rWph19L1BOLbmQ/5M0YHg5Latt8jFHDWY1LL6fEdy42HhoOdCXag9psEpHt7QiUO87pSCivFu
begCzJcNe/18IKFovkUOwm2mqHW6DGtngNwKY+2ZDmxhhz+1UCxy5l8PKBwPjqD5TrrPOr/aid1/
JTXPb20XEnItGTYyucatwsNai0CROjaJR7Sq1HtlO1JWX5IbdajyYHfAh/SEPYgp21Km6G3287B9
eeIBlZ+4EZq5T7qz3OKKegBGhcxh9fc4KHDVe1ZSXag7A7YRB/wGE/eCUlyplVZZEhVwj5SUIBlp
gX9v1PRTNQ//R0Msr8wLfLkfC0UD7PfL00u2IOj66LjSjBwlMW5yd8/jcg7IgsXJhh3xXK8wJVXe
K6W598vojfgTbxUKKEitOs6zy84cXOo/3Ktvck3IcdXaIproYhNqb8OcFviFHVfIbYvn6NCH1qJK
0bObJqTPcDihcbENlCoH9zlyZP4n+DB2LSWgu3j71WLuYqWramDH4AzeJQG+hmHhaxYk//y1wGzG
9LnYbzlal4cMxYjsXnJJA6WFyCvXZYL0fwUPKIqU47vMreCJ3xmdOj3C4mWaVRvCla0+hKH9foGj
mnVYzcIqqYHhvDSCRWjmzjO20zIdxqj5Kf8PcQYCOpAwjS4ZctQbY9hSlBmn6NgQhe6oJFO90JDF
B3MZl0BhmEL+Gz+LdZOH9NV+S6jyyYdk36SupJUpPbsF9ONGbBxiOkiMFP4TBtC5apV/iwD23ZvK
Dtwqjga5bPwkMOnav+33J4FIPK8XLQXwFWD/JuCAtn5kceityqsP4cKSgmEXNNI9loblMaGTVEuF
BARWveFfgZdrB0NJoXhhgbfmvBvM5HbU8swqVsFpGqbRwpW38DiWeVkX323EmJvgNgtWm2U1G2NQ
6+xS/U8rEVhxZ+pnS6lqBDhKnzeRti9tbtpL5I9WtlHAu82I5FYvp6+yNi/kXs/KDIfp9GGpoSqn
dFD0fAXQqQ23RIqh0DTvN99SGpdTaFg5Nb5UsjoFG+3R3WDlzygeZKZF6YvSMg5GFMovC2pOAuaH
Vi3jG1GmNl7y3yzKJKO2nWUlOdMZPwikE+G5VrNzDbUsD1WLXkD30RNyA8PUeKYPLx+Lxomo2TGu
rT75x09bCkOQ8fhUC7oTv/LYeAILPRrCiwtd9X1wQ0P/LHsDIThn7bxyWrKa6GOncmp0krdQMJLI
TTUNLofzbr4IcSx+JtZQmTjV+sX7v3kSyAbsPAIvLc7t34XUbrjW/pXKjy6JkV/d3ihrwEQhGrMA
2F0y2BN5WvXVC2bg/Huad5mgWMtFBS/jp5/qsICJqEKWa9AFDUgVUsNZqfD6lLEgmbO+xlL4fgw7
iEz/Z+W4vUt6puW7rtV5pa6gXkSRVqgocjYZA0rGrbqZbHzJGO/tt+X1SkjnoIuNRUQRi5X7p3HL
76+oHu6ImK94vNkOpYfS04/m1bjCRbh2nAEWCmMc5l5eWSQI1meUTumuSwEGIR9P9oPBE1rBYmVj
jv+ETBqxxnGWpqVnG4g3GQNx1ckBIouwQ2U4Lmb2gL8qRbYS8TTsBYTWNPC6NqvZoguigGDR6jcq
yd6QWF1FBGu/dvMqNPWgr4eurOlACeW/ljQ44JjQ1Rlfos8qpk5CvSFELflAlfsIvjRrM//Rn3z1
KLWqzQ0LwF1s8FDyvzj0908CWNpY9ngtUI1hZqcoFZsJ2JQ5D9IG6zB1hmW1aHBCAFNEj/umixK7
J4ywjQsut0zaRHP56Ai08UdjlcQUs+7j+hObCFVToRYP8uA0FhgfUaAmqSZrJdqhFb1y5i4XiH0M
CbAOUhwpGng4aD5FAf7vLOlHEFG5+MQp7O2rcpaFvp6AnEfLNLgpE7V7evSmBz5p+lx40NkFXOKG
iYgzmXv9zwDRPwYFenSK9qUYt+BmrwJuSJCN83TZIFHP5C4D1QrHShE2/cctuaRGkDfWp85HlpRq
1TjAesueshfa6Y8scEA00kZK9qNPCzmQTMyYrItR/ofbf57vPYZum6revD2vtHPO65sVRf/cx63B
c58mctQnivwd1a9tQ1otMZXJxiw+Z/KNdM+dyjYxWzS1BzDyWBTVfKc+u08f+7JdbPccMlRM9LSl
U9zTIl3/2IR8qTuDjGT2FvT23rxnsLy2MkBrWPpV8X5JJZRIi2nrWjd+ABw3WKy3DBKSeS0QtJpZ
yMAsoRXdWw5B/hB3itkT6s1R9dGW/kCnNSd6pqme6CGoDLrAySecg2Magba6kWeKDwIDqmlT3LVN
xu4xwVvnOXh+DeafRM0yV1N/Xwiawn2KLpNl71awDR91iZMXY43MNfQ89LVTbXu1wbutxQEvzDkM
AVMAa0TEeNXPQpYEzjdjloQgiwbGsOXh18a8ZHw3yEAjDwbmNN8cqj6niHTnhGEGB8e2j+Y3ui7T
gPBviUvaTboDVPE2syLLVIZJBMw+cJO5pGQ6uUUKynlKJ5ii1GfYFRpONtmY7woZ6t850KJxnl17
LxfUC4U7sS+RqBK1v+bUmRoEp10vsL7C2nD8s9fw4vWHKant8fF2MS5D5zbc6hLwHSxczzKXQAGm
y40k/OEM15/sgmxWuxX4zRuqpnFvnoIjEmHmhgEUHZPRxxp0KBdG42bJK3A0KbFWWsJfd6FipTO2
8K5Kg8x2I1gKD8h1gqQYehA/8rU9VBMjkkatVDIBs0mVyYnR1GwyzV/sW2Lknb4j38j16xL+YaZw
ogE0VSkngsVfV7c+dteb0joLcE81hzRyJwHEEOigysA3u8vjfHFJ4JrTYNT7FQp0yRhnR6e0W8fE
QCMZqBxaU7DGR55tWUIxKQeBBqAH+y5NzGfmOYwAbJnHbcHpeOfSV6RF4rrsRESaacH1Wj3qe2cD
cxpby0so14IF8ZFykk4WaZduNeChGFP6b0PgFyUW0QdsNZfVHqCkJ84VuZx5lRqChn/fl3wRQScE
AJRhsXrOl1DWmp32XMJQUpO4kGWq9IngiicGaw7SGbWcVZd6pNoNWo/aqDguidb0S+EbRSm2gM3L
UP2JxrMR5ABh9j42QcNGNfvFjXpb+A4pDp4glJza3mdKSGuEeeLOwdk925TGAhzx7FaOwafHIZvd
QSiXwpshTKPVd5BzF7RyRw9QTFvgFsvyDil8Xqz2SqJ3kWj7k4s5IfD3z94hnESbVhov1nP3FzGI
jto0N4FJTyY63J5uUX1KrSVR9vXRhxZwdebO7TMifVAYqj7U7PdpHedpFqlAG4sExgkfEp4hcZ7C
JFx24+vFYhzDoWimaxrgecZKLybe7ZAIAdf8KaYSON7vnEZOWxt27Bvl03pvqy/ckl1oZjWVX1TQ
0eZ3GXpgGsGvu6gHp60BP3khDQgVms9wWf8GK0QZRnWQ3n8w8KnJeVobX5wCt5mcBNm+97QoZ/Xf
BpBU4iFAXfi+OqonB9GO2Jc9SAVBDV5lhBCrsTjLPE2bIXM11+OfX7T7u3P+izj0rHAlhbLxIxK5
JamECYe3zG1C6grIrrpi/P8B1R4j0BdLMRUFXEl6xK0Z5UedG8yklpnSJB2SOpOVd/mKy9SEqT5u
Dp34Lq80T+aXFD7cSMalKTJ6aIHthIP344QuFlqRuzXWdd5vkF45qmvTL/XwQA7nUA/sPk0zOR4y
JPAo4vuN+lNzrF5UWuGPKan4brqWCvsvfHHDVEhO0eZHyCHBo9NiiR5wWKijaNRAY5X7CQFm57zP
fGE1YSJ7wH8yU6uNjyZ5QPzPVTw9+eOv7TVtOHl7GNWl1HuzuaYGKK54P+1ckfMvYD6hGWh4m9CB
8ZJJgyw73IjMfkUCbq5PaXpecD57zkCjMJMc2Jx3z3KO9Bq+IHWEn5G6O0OO8QiYHeTf2aLamkkQ
lHGivciGbk1J8q4+Gj+K8GwUOOjOlkuT7XdLwp4xFNBlIc3ba3emVfSSONNtUf9RFMrq2wo1HD2j
Rdhc9h8zm38CWmjWN2sptnC9ZNP1zyFIhbU88xCWn/aszzDt7Ry6RtGa6l+RK9DQ/IIzWr66pmfc
41OC+6la0y/NTyIVdcbVL1oICSM3D1oWUK6i3sUK5sJ4dTY50kNBP10/5P1lrSqd5JgzLRK3HXxe
hV7yqXrigFbYh82c/zVI5rAM8y0jMR1K3q87H3m64ibfp/LREh5519lt2MgTrVY1b/KqMXpbeYEN
j0ahrTDCYXHQW5pR5Ya8K8NszzDtsdFwKfHIqWsipySVsLGb0+AWpjpXp1ItAW8koydL+cJpT11M
UDOgVLdRRVtbsYgr3GTWHNfriesaBQ/fuXSyuZtmkwf6xynA9Hoq8i2zUioFaRBf6jFkgAkDzoGg
jLqVlzN3DkIRxP4ey5vf682KXCfShV0nzNdYD/4TR9FYft3ETPr/k8UionYpSbyW9O7SyFe7o5P9
O/0wzWDZ5tThm0LBNrlsXRpRiEc4k1ActlEmbrqUdIrZEWRAdUFxlN4qMtLaHnDdMa35m9PPsFEh
7970Zb9oMZkvkwl07fDJ4yU1YGMeedjnfLULwOV5kZD4FOjziT5NZ84KIa20I4pkJiFSjbWjaxOB
SecrAdzyHK70RoV0rJDWje69iOhsakn6ZdhtjURQPcGbgp6AWIguJijPPxzGrpnFqudtfmC5FnZQ
cje0OoQ0U/AwCv1dzOkaYGoqybbIb9agq0yCDkcahNsIwnhw+ncHCUxrL6dNndySicsN1656yjMp
ny7g75ZZKngzR3yR3CowlshKuH6XiTF2GMexSJt48dlm22Y5cSS9OLeET+ziLvKp946P0woQgU/g
FNACYunUJcfbx05hTYtVBU+ITIxFcUB+vK+0yQNAWVeB8GReDkioY5BuKninCq4U7NnRl199SZ3K
nQ6dJh2dXTr9uVYnX6RrSefwgSj0P4S7HpVhyt2ZP5DGBpVC4iUyGJ1Bo9QjpOd4aRhgxThak1cV
tfUjuOpUe5LDGkd1PxCnCUb38Fbfom0U9xQZ1py51WJkWFVm00FMJcfvJ+FQ+xNSanK8BEgWDhbC
ZrVZYET0fCobFLElgYHjFBMWZ2V/9Z3GyqwsYgB1Ul9tvksROGHpZAGutXf729mfwBuRC9vbgf3B
jq+95geDEjtTN9kS/0x+JK2bH0Tdmii+sJlE0utMT+OLT7rCsy1NrdIha/n/G+B0VUBb4p6PD694
vZwN/NZiqCMATnckRUZfGkm7xkGXE/Y0BXH+Y4riuhsKzNrcC6b+H3bvkPt2DfA8kCEiqo/E/ews
5gptyi5oH7OPiDFSVGmf2a4ttGK2i/5JIaLUhTjcaulNWXvGOUCEpxyoIEs9vH4AZL54BzBUDO+9
oDKv6P9D1lccJEMIfFC0fyC9u6/ViOJ7mLhqw1PXfY6Xy6Jdn+rwVtXCeAfljWIQdXUVh2OIyHJE
91lbsVdYFJKSQ9bmIg2/M9dYeKgwjwwcHObibT0gxO1FvEbpmrtUjSJCUM2rP+QHyyRtpLNcoH9l
eecwH8yJjE7NSbCi5UJG6ze1rFlHgMSLxX/KnvUXe4Kgcx+xkpvQc8NYB8xLwQmlV9M85w1o4VhG
CGua5ATBKRfQHzKFjTO2eQokRG8Fv2KCbMGLijrv6Pinn9oKpK4epH1HyzXfGuHChDm5M48XN0PG
t292KlYuaLpH/+SUfcRJTuOEzXs9SwZ1rJsycDleu8G3PyP96uzf+u4c38KWXKhSE1pZlnEY2Ohq
jw+XV3hE6VQqHj8ltESjSl0UXt1twiSwBOPVdNzGZUPBQJxBuwvoYyyPzzqN0GTYLJey6DIGObXU
HDhxz5AuYHBKWO+YY8Ix9f3w8FP+rqVAshhof04+KMrlGBBU2uhsOpQ9emtn6tSAF+PJQGmqo95c
TDv+6XscBt2DHbIpQR9w2rIke6MsO8r5inVbDSe6CY5GRlR2q5/ERmEyrGFDFURuXUOvQ42M7UKz
ZfW/CbFLsVotr+7IQfBr2hiv+6t+G/qad4Z1dS1pk6XQf5Q72xYC/hosqRzLIoPHtkEPizdNtBwF
DNHkdvK9DyHJfCA+djsHrve42I62spqWq5C4Gj9Gi1ZpgVkgITfTFuFhUKbwZYBiFsiIoZxnAqaE
fg65FwzWPAlqQH0WotLRCISagtEfhVDXyYgPLkvdM1BJ5lCpliBelromM90tL0xMVh/Z2ui3feCj
mKjunIYbt+LOQiW1TNtZTuc4DFEgmFmCMEGBTnEY9nLOCVq3s/v6M0p+THg/I/6s1wMi3CrukK55
AkSLCsY1GLa9dUSYILs/PR+kQJOtCHTmmtrNRSsJ0BZ7Pi4RqvEdbOaaqnwuRGGw1lw3zT6A2Jt+
rhzqhmAZsWgdv75Z4IDXzwOhxGItejyaZposvgjxLhK2XmptwDKkUYvBOdVBgNgvHf8fQXN6u4eh
b8gU4xsFjAuoE/xU4WyjsPfTNwmZlnEfSsX57tZf9yCTDT8+AciD8IrY5E1ArEp++0Pz96LCK7VJ
jbELFWjk8rFFPy/raqFgc98PvVcqsRJmhYrC6gAy6YmaooGN1YK/+qse3CXI9nl4ihnPKrpaEYKb
6i+F06FAB6YVds51PhZp230Qbjl5gZ+fT8+77Xkw9Tum5RhFKA91bFQvmgWmAiRc6/xP7nDHKNM4
Za+CvwJqTZyLTqKVk9NaCEBzGzMuHJLu9y/Kd9qYcGx7DF7xX4lblHDhhKRBMKQJAb8Ja4aqmVTM
AILTOci2NGKbWVLVbVgPS83PteXoDPu1YivRCu98JTyx+VU+hAzunuusGVeN7i8ir2cmVcmM0g4c
QF6Ho1Oayg7jWKz6weehmnBrtjXCqp1RxCWmMpJzeaYNfIiK+xsRMABOu0A4kfOrlEa+p5EuqWgT
lZlnzg+I7LdQIl3+Bz+UgMBVWBNzf8h+YmgtDe1s18B6Igc0GweXnTNnJKmJUFSVYbbouWtnBZBU
NvAfmt5yhC3MhgY87C2YTHw2SFQpCzSSMOjgKpCTlDCVJjyOMbC2b232rCIS4iPnMoyf5ojqdO3g
IbeocSyu5EWTypT8sbJeVKiXhsGgL1nb4Ynlb1/0+QLFbC6oe65h1FtjKzDZSLL53LgpB++aOYGT
XndZ4rCLl9goYN6F0fYTCBAckfHp23TU+LagTMRIDxHkgSGoNZcSLDEH38/modT2wSk8dyon3nGD
FQXuuI1PC4XbZ5PIvY902J+krj/qEZ3WkxejU6g0XzEzyuuLQMAVLscwTklra6BYYh68W7S+WNwO
KGk0QsiJ1U6UjemYHFWvsMuAeZ08NZ3YxlR3EcyK5p6BFpvHEBmSi0dJ1Mvh3zUlaTZ7mr03dp3b
8Y7KVVMZyt/uTJFVyhv5/iB8rZXopYjWVW66zTGqy1K6VfT8iPtNfEDEH6oBT+M8DIJigDPdJgKa
E5qsVZZEfm284C9P5rrt54VM4XLeRZfFgutgYIz8e2uSSA9moC+O6XE9CwK+TFoqYZ2JzNvhM/fI
cATigOtHWw5TClp7EIToHjPHgkRgHkj/IiWB92KzDLoTpKjy0qJqKXFPSckm1tPIy3/Kb9qW5TB9
JYIM6mS3eJYDWGVLG3awCDTQ11+4kiSbRQ5yEz39gySvR//q246sQ387T/0t4eGs6OSt1JLCz2me
2Fz1eedBO4A9wpRgXlZRRt6FCnt3opSqA4RtUgLS/J0qEQDl48/MEneUWzBh4RFrU56KMXQR+kV2
ztk0DEQTFCc0wFkVk0GATXcs6QwsTpvNpWcdTB/HYHd0DPF25L8z5jIrI47HkhkT4oMSKdWf7Lpg
Xn1+XKvMlaQ0DN6hX0ROUYRW2dT1MX2Xri7FKF2CFYKkzQUe0ocMJ+EnlrAK62y517b1id5F+wDK
dEUhoFCAFYVQFOIp5ZCFnkw4kvcvDl9i9J0CA5pPdrbEhqmEU3wF02ng7TIbqqWd5epSJQ+ZV4Sq
B7xOiVVhLG0gjr+oxSToeKo7QcO71OGuL9T7yzFKKGvcISaVdmHgkfdSBJz3T4Hv9EOrBdc/a4+C
oMYtMYuniJPQYef9GK4ieCjeelrRSF05OrGvWdVsXOdFQqUTh0KeVgE+M8KR51eNZB7gjzorczTE
N0AdXUbZmWAvHb8K0V8LdPXV+hu2DDbpys3X3OkDxnoqpMPCt7A+u4q3JGFV+BfsJ8Zz6TwNV4fL
lEqGvYPD35k+69f/7Yxn3IVFNo51ev+JAxvPiPJfr1iyhzwEdfQbKJlr6jhqjk5oURwxKOLNVwQA
y7cIfydZLfa4npBws234ti239pJfyJCF/gU1SRvWRcJlJCJaGc7W5a/BoZA/QwNMU11r8aF4oWR2
83IPMU4fmmAQvOzaY8A4h396Zs12ScoS9bbI78oYyncxNz1Q5TLpBOdtFmYwTJmf7/yXvU4hdqyD
HaxAAMZwCjtJ+EoY3OmdoFD3dwgrkZd8Rd1xuTxJIFWBP+k46Gv5Vj0oqIhWbjqC1sXMBJRiZaB9
FIbq9Gb526annhooikp+I/N/Qu4mgM4YH1nafaeIDhhpsULjSYQnjFfSuipmMaQUrMfJLij8gx52
4UT8cjc+tSp5pfSAL+oSEmwMh9QikDbWCpNBGByJi126Sw8c3edNUJY4xVRtFyIVZhZti7xz6guk
zgNKRWEmBJ0ImF4DhsyPc49Ih0j/youaOY2Ts+QzBX7befK5LHsYUYNsa5mEALiW4gDPgpFHMtyI
vMTMNyhS5zFMnL8y0jiqfhK9bFBYaHoaU/ORtuSeGhreNaoAbtv6CMk7hOf7tFdfNKHRXLENzYQE
PFZOSKtsQxdzAWUSqWlBscvMLuuWb5LR1m93B2TpQNdzLIyGVrkviEk5390juij8K9E+AoXXZkJV
KMPtJ6NGpxFyVKQAan800qJPcgBLvL0WgpPn4XKa3HkNWxPyKUqor1odzE8eIBgEDTnLPqhxIIGA
p4B2Oz1AhvAFtNNRYbMhNHSM6OLOvQRksWa3J2ssHgtpp64442F86fG65z7pQud3svL/4z0CIXWi
njDmNcDYIPsevBm5VcuOfiJa4UxD/Pj1CT3/A1k11CSM+70mn/lzRYL4bTobvxvgGVRwDb1+9e4l
oQEplv0VnRlB2hXvgt0hVqKlqOGJ4M1nt2atSPZUbP7H6ji1hUFH3m2CfJ7mvtzYSxcdsiVEnF7h
djoyeXKoazkWsysYciPkqU72q/Out+FkJ5TkyPd5I4KZHTHw57wrerm12I05LPLHcummbT4HXd6g
Vd+lF6RF0tmw5+xF7lwkLeYXKCDbexaywFRI5uYOZ5t/q2UNcKRpHp2c6AssD6ga5WalT5WpjExM
Kf8G+G8ApGXuhB2+d7o4VJtJq4b49dYdzf3zl9zQe234UiB+6r+2KS5zt90SSlVK0MgJg9ozkeuW
ejFh7H4CFkRwHJguPlAZqfUoYXHbFewHo+PooWamQCd+36r4evfIwSFQo6CAdE14ByNBStoiWx/Z
KXQj7Q0TgjS2Tceb080zrRAkKJFzDUHnAkxQx1IJG4My0fYqtSxv/q823sfRgEhegTOcpyTW8X4c
yIVmAHdqA5IeYkAW4SEkZq5EGE1CV5H7L+9mSDok/uIHVJ+Q2A3ZwNV2t5Q6zUB32UodxW7Y0Ip2
YLSDHm0sQUV5TvgTRI2SRb/G2X9FtJ6XCgN9ytiHRs0Tc91j1WuOZxVMGDhSGk9vZttO58YuJTXA
6M/JW31Don38zPVMHtEmWkLNddPLU9bKALztTVx7D0HHiqfUEJiYBT1XHQemKZqHMgFKyAs/W1AE
pP52LnJv17VJS1Dy1CERcTBBeqogj+SMMjDJVvOV2zlLGncIgyIDbjIEIs+QPpth75/YI8FIQDaK
d2FHZqMExlegzaVjOnA7MroZpJoogn0NAE2Vc/WaeWfdeaJW02nTb27Xhpa/qBhBpwDyzCnIW6RK
I4CKwMBb2s05YXbdGG/z/hdjkyF3yg63b40ooQL2RnOIRZwCYC/A9SLxR6B9zbPRbN8xwJsQ57Z/
xQx0RzTnCpedUs7plAKiVs54Yp50IkgBzIkGyc1w5YonfGh4AIsme4Gr9WKlKscH4+xUA+80eRhJ
JhBvB1ota/E2CG6s7JKvIEgoUQSzZTVHuYYdZID+HPSg3nRbG/Q6zQTO8dELofCMjKFYNvDLO4hA
mkymDo53XuqhsdHN4XLqhL2y85OgTNqEVvQpMYM7S9gDrHne+wdxk47KzWh8x0dWWaD2i7osRI/X
40e27kawpJ8Fk95nxroaq41mLX+J9rxj8hWdKs2tkami7jLYBIc50EsTotfwQSoH+ZM5DZKUySUd
c/EyYScMNUfEFaaGdgGY94CWlvHKIt7m8ZFlR+21blszVtP5IL44yDJ333xbcm2YRiZQTJvGDF09
KkyTNoT6zzyvs7HnQI2ot1cQ7Z0rvNanTExEByMPEqjfL0lHFsQdzbfk+/mUo/ZzRpHiNzf+jnlQ
OiAaGK6AIYtOh0ovv6rpFdPEgMYFdtR4GrwzuPFUxGS0Q/Q6oLlLufjuEMXngOtYm3JAcyEPPbW0
5Hy1MmT766E7zjPQyxI2TWQHmkifIPxW5oNiAZYbsJRCgQmcDqPJcbUdmpLZxsTtpetV8o8PczvV
FWyNoH5QUH0m99T5I9S5iqwQwwQLqx6g9CIJoif4LIQB2zoO4DdtVTrCDve1Gz4eD7PYBfk8wSPJ
IS0EwB04y6oUN/d5/LepIkA3K7kv2IFNrMf1tf+Bz2jT9WTgvZAvfPseXlRHhNQod/VUP7O/Rouh
ZhWD4ITNC/0OQb0BGhsjBnx8yp9bCypC1InmU/M5ppXwgA2u5bQAg+ZN3/HoUh+DaGdtlHM+Jdmk
Tna+fXRuiX2mDq44MRhhwcSr05uKjMHfr9ybHhqb16sO7/3m+AgH+D1aL21jqHPWP1/kGTfI1SHA
mP2Q/znd445hWViVg77sd5jg0MRNXE9M1HW9uWZd+y/ZxabD2mpTEiFs80sbbnTne40HM7nQJGRE
RcGLF7NgoyF+JYdOS8EMpbMTGq7YQNQPZuLoWYylzPHdX3ExXpXnWGzZ5hMyV+TPbCAzNFlXaTTT
69Teks0pJVIO69AEG6JFatkbHMpbxbvrXgLjByKUC1/ZaWIaaVnwy0D9PP8Y6Dh27A5rPfrL9K/d
9ocWVlCsE7FfOu9GSmqkizXE3hSuIKtvCpPEi721+TmpGTkZMI6F6ihJ0NCfld0HAIOzITYgBHB+
QMZHVzTCfRQ0xvXU6FiocsDkWiH1fZQcrHWmevQpJOVSpLBA69y5EP3YmkCQ8j78BUsTVX9b/hkt
BMXtUhsbXKO4v0a7sVvbHSFWZiZem7+fWmdxRq/qAxS/kp1gtmK+l4nuqOELl4FMcRSnbM7uUlHG
2eK3FxSUSbN2JykOw9Q0F/IDQTgGbP+rE40XeCTLP/HsgpPEtaw0P4OPKDjdcsvXVLVJFY7EYKzg
2oMxxWdnsi0dWwgpYREucbO/NNGCdzI74qaEE4IIYG2JlCHhLDNyZUJqq1nVx1c/tNJiRQ6vxae4
guXxVAfx3JjdUGYQd4dg2sdlRiQmKCjCRe/Nevji72m2evMxDHEEg/O6GYr91sI8GpaJbleWVQ+3
2szsShOcJhrYHW4pB1iYUsWYnzBvWkx44XwfvOglsMLIwMdmsyCrfQAXrJLhwpecDA6vjlwe85de
ZZl7u7tcyeHWJ1LcCN56eo2qTBA5tDjo3W9TxvwHltK1wcfOMwtOQmoPF9OBIxIVs8kNWKBLFxhP
DnQ84Wl+7bkqG0oJ4F3cWwO8++iVKqLAXU5/2MJ5BaPGrIPFEcvsAK/3v70WRqEpH8LfyfRvSQR7
I5ptxvlB3km1bEgjsoFnQuDHRW9nQxm3hr/Uu62oQQDOoQKKmD1EToTcpvNNHS8c3UG4RbdurYEt
m60I48TT2XJxiE/0ihfOYmkIc/UdrO7taYEdYPJAUouWiAH1rQrNdOhoteHHLDi8dVaRJfJ8FtH5
SoFo6PrnscUHmIa2sTCUUjdCVIDV14mqWDyrzDNIUJ4J+IFy6IRmPDNzPO47SpcFmj9zi5IrE3Z0
gPYEYGjOLaDgA1lfcu2FXoxJn3elUzW4L9RskZfR/n70Su97Wyv5utVx48xyip+NVtFK/aRKQGk5
gjrjBqC7USPi8G0CXp8vtmTC36DcCUja9/MW3DApL6d81i1hLYe1CfHJVqb0pujmw71x2Bnwdvgt
gSMTf/mu9+fR7K/CL4++3Y2ZCFwxTJm1t95i5I27rLhFzMj+gQdxc+sXL+kDPNNTyTWmCtEKgR2U
4UgNHMXW8yl8ZPrII97SMbhqyuRaxpGerE3v4eTDQcHAA5b+IvVLsT2Httf18HnGjJ3YeiNsV37o
SHGlTYXAjKW9f8twSxcuU55vbBhZ4WZrkqr5BHvwP46CDg9s+RcY/0n9swUMEVEU1FL/wVnTiAU2
HTXI8G/mgWalkEBUCdcIT8jix8i/U9BGQsSFM7rvHmsNKD4gXIuJf1Em4TDzUo+zr/KyQMF2m6t7
HNwTXQUiPvpIx2Ep5231Fz30ebiMKVXKwA9AR37CTITFerTLQelKhKEzzVRT+h43EE6oWdD2oMAg
+UzQzl+IVQBAtvfUDiJGVrrfe7NuQV2aOnJXcrPLZU5DXN+vnYyKvlTcJofSM8UmjWE/xUyZHZk2
/hZ2n7i24aCScQHunrQHIA0X6urM9d7vNc5OEZsKLN9wAoAM9t0iOLPiiMg8x9x5grRPIJa11iIs
eXt84sAIANqiSD2eGQ27PeFebDclDZfaSf4qMF7Mej38Khhmi+jhiF9sZyRoLHMf+Mvyv0nvj5cT
h/4K9BxuiXzCvBjv0avL4czYALgRrVIqZZwX222zhmqko42Xy7VsIapwBBTYpjYag8gKGeSLh3+6
SYTW3cpxHJkExDp9r4JrxfBVIhPyCx3E5z0B6ZPW6r9q1SWYtpzNGCz9VErv6XNN5n2Evf3e3785
gnmXOl/No9BZgjMYyNxsq1vFPJZ53FcnEJANTtIIbLEpJUtnf08MFf03TcVdXAfJa391viZr1zBL
q2dSp45QJi1Vb14j1ZdHVhe+r4BsVIAtprcS8gFjEbPpHSfgr2Te6xP/MPNYt5xH4W0ulzbauj8I
hIGoebhCECEewqYFLhCmaomCqZkjvHb8DxODtVVy4PiG80Bz1VBaZ+ChOc806ql8HlEQNbe6BdTv
rMrs70d0c5FLlq+hA00J8zG8wTzM0gMumGhFSePL/47AsjBtXYMlswc2krDm8LZHfD0QqgA7CbFF
63fUnzrpJqRdoBY139/ZrWTQSNTm7zxch6OPbDCAxcG5EQ7KtpQMo0bH5MSPDi2c3vxc6NpmhwAz
dq57B70d4bBERehnJ7wLLBnF5Yuv/rdvNCJZTWqhSoLAtsv2cN/tPiSeFKYLq3rR1VTf41bJViZ9
MvaPHxx42uGdGMwwB5vMT8AeobcEkY6GdCCB1dE9DVaeJBvtkAXbP44jwKTUnS+pAtmCxcUyj0i6
R/DBlSh30g/4wbelZ6t/X4yVnC9/zOBf0EDBEoOahOywbDpedWCKnLmUyn1QdfNeF0VFpTAXlCZn
7u5sTo5o5AqAxPCKFnm5wvGT3Qp1JKyszowOtCJw08K1Rk957u/JM10e7U1XMUKObQwYEFoIbfp3
Pl5Q2N5RX0sTXnglHh0JmEI/druXfD+UFgDLL9PzkxrfRwZe1fopxkRuv5u2YyTk1DMaRzG8vN52
tnfNzfuGJeOypD3yPM65AAuDo43oq6xOYRRQaNaDHsu6mKAHqpGOBysIK0JbwNB1WQcD9r9gYqNu
M6eVHiUhs3NQBdDUMBwfW/Oe+Jy5ivfPfrKGtSv95/Av8GhJoOqnsQrRpfhzRFNphdseJwXfzf+7
/oc5WwpBS+tucOkR+fTFvNp2PZesvqjVigiGoRupZuKFcVTT1a7MUqyoK7HBSR4JDJvizKwn6xf6
JCU5HnB08O8LDpRignl6AQEC9lQysn6aH4ZnZK7C00FwiItYpou9/MZ1E1jNVPA3CtoCnx/28D1F
PttH7LFBKaZX0xkiO/nC/+3Hea8ibOXTslsY6HL5izeN+DrnMIJ4/+5eKAvzQPUh/k+bYNvanlWe
xZCSPUd7X/ltZ2tXHvkUzMZvUQc/Ibn4dbaTHhDIb8lIROx8WVgwuuYs65rYsBc+xWjKV/V4SXl7
MpbpXYrEsWU61D7zidOPErrrPi2sgi/XEgpftpQ8hEwxAH8xa2OPoKcwQe247Z2hBHrTrlRyZRY7
/3mx7YNj6WFTW3sMl08ryWDfZ8V6vw/8WltIj5RLK8rU8x7FjUc/G5Oj3g1LxLcwCjdCHGCKO5cs
9ByRvF1tPh3qlj10qUrI2tvLtaCaf1UZKIr+wszxQ7LT36Hj8oBVOJgkJl+o42pFiq76dpuELFlL
W6ZsLcoZ5m2fm0Ucs281anqvFWKNoaJqgA8WwkK6voY+i9oOsftuUD/xzNw1DvVUPHry8Ce7Zz/d
mK0KL+LB3B5EBBza/DXOcMQ+CZHXSdr6NimQiAfVoWwgkUKdcqmVwJ9DRO2lSZB6Qq6g4Om7aUxG
820zh1nwYDcZNhyn2I2IwpQT0fapaufZKAcpXzJT3Ip1NsJSuvZtAToVKMCnSldjI+QWI6z27/g7
EPj3l6elqg56JM1l0pWB9UBXbuyWPJ+LIWUwcyL5LOw09+9N7IFhRUAyLovuM3fltGgEsR9j6gkZ
Mp2Zb0Rp7vheZ3exnzr3Y+DUSuamf4e2IQnWHi93GLNthcHmfafN3DedsSsi72MPE0glsKayQKIj
ZvJ/pkXUUyywngmJ/qH/jQRWKCaLzYl28yaADiqjjFCZWTVPUycrbiGJzgYIJURaeSvh52trroUg
qgR2lzraxZ9f9TMokE0D3gE8PL09DNULm4IGk3vl2Kvdnp/ERR8zkE4cgYo+8I2vOfaDUSt5ib58
tgzr1dBALTKpVafxtRk1zfWa+fBN3yoNjOdi1mWZuL65W5UHAJsXZz7LjUsmr+DMGjHSDAp8J6Em
QiSbQBG3AWCHhVF1qtw76Ews3EJ82CBQHI5KKRjcBG9ov8yBoR8SFoNRN2EpWyZORDXQ4xiro8Uh
S7cuK9ZZ/oaXO3spbqcgPmlPdaPfr+G9QddSaslpXVBu0Pjy876YOog65wmjfN9oca9kd7ddtOzo
HqJorBao2/KaIvbpGV4LQJAs0HVL/K7tplbUcroOjT9Adv4Oqki/Ztdsh0Wc6Fn69INj5cTDTbo8
VTt+WQ83DtSc0mJlZI0bHsXtAigxqbb1oDux53qjiKC/A9/1XY3oll6WNLtqtsTb5EetWDG8/agK
35NrmPafb+CvMEtnFdk+RJRJ+lKEcLgWJwYovIhxR+7jNbYPz9k6gMOE5x0v2tvcLfHi273hfGTq
0Uy8OvzeVUvhKU7l4L2M/ROGS+QjKnJEMcmbor0jYzKXz2/AUTKGJiTx+uwa2lJJ9oCmg/gm2A5i
k7zxoyFa3NBACLBtQLm9Otvmy6tsx8CoGn3sfYx5LypKqsGfnSZXSfkS+NYd84oZQ4HZxkangEZv
7XkwJdbUxNtwSPHUdn0R/dzkO2oN/579foNmuMABYgE7oOXic6Q/Qx3vGqMQOx+QFPzJFHzh0L35
vP75a0gMXgOmqqn7wMI4I69/2UyrV0DMk/epsbb7ykT5w1t3MdIQiwhLqpOWFuTDthih4SnUOm1N
4GkSJExBcR10QK1r+t5H8V87JmPiKE+Dj4OIFlXLYKCWaIf+3s1L3dVWAU2VaRSr8TZ41BC146U+
yzvOTH76gHZLSjH2o57o9zpnh7K4C0y/gG/KBRrNUPOFeEgZTEHeVqfHgBwRk6oz6OVRVQ0VMOBK
ZDn8SDiTvXybju/QzRmZteGIXTHxbEfIDeV0TMU+CstKdYNq6cS2j1KMhmAuckiyoux38BbsoMUQ
IN4Bd3LQghvY4K6EAvf4jzlJo96JrJ01RFxS5vpNs2Fxc4326KNJsb77/yWZR5A01Sgl8YwKI0ID
5usZUFdxkjmx9l6DRrmZV+SmHD51zcSKGpvLMCplNkE3sntzjYvDZ7oyrEp+hnuomkNKzeO+lWyA
NeMbN9H2v4gIpCkjXgsnSpdqWetAU3vmKLeFuA1/UeB3Jtq30UVOdIzWGk3gWmV1T9gpg5dPK4vR
TSxb4VgR7bJTo3hyNsh4P3YsNvC5ZO0UXw+bvhJEiLn6bWFz1CsiWbHnozEEMjjxwsy2TLZY7q0l
w/4JIKBHcKWhcf1NIBtE2PFFqF+oszDkVQ+4yjftnPJkiYZMbOKKL9rErpVPu7rzRlpmCi3WFwSc
6hhDyPXF3dojOGkV2236s9e7Ax7zGfJ84eypezwCb2+AIUfegUG269r+5tPwLTFRQQMEq+PQt2x9
brhxv6Oq8/lTLaD5iRBpWHfFupraZxxWoD7squcnnwYP5awu3ilsWKnOBitxFKGBSqs4X3I75XZD
IUiQtJ5DlW1tHUZTlIT6IyVxSIGcgIX1MK2SbqYHdDuO/I3L5NH6T76YqBfTgNzBY+3d4ssG+35s
4cRiIBznPkjAY7Jt7rB22wymFYClaS2FUEUegEIPwR5+UpNO+b3EfK+yNvqvAvTVroY65qo7fA0y
zfSHG7IqJIp1bX11N2/eHDNluTcgH0g97GsA3r0sq3cho9hMLtMLXFEo5sGiTCUaZn3ullccKP9z
4zq+7ajDAhRU1iUVUnWF5Yh1i1wij/W6sNgdRf0C6P0rcD3Y4kTXitlL2099thh9TN29uj74cl7v
pHksXIX2FOa+pIj+YL5UQRAipb5yOCKG8+P7qvCxrf33ozvkQYu29Qof11PZDliSAOBGy7xuwKL1
Tx5rN9+/b3QNr8eniLWKVtD9hiftoHL8I+Da5tDGMAFpqNS5HO9tZ0FlR4Wvu+lHW3nde/pJ11L6
QMwZCgXzQWsCU45inL2cWQz2jYHw01B6ZP571JTBrSgJO56jMjOWuVZd1j/2tdxWv18h5jq6TRRk
D8W6A503s8ANNjthILOiSywCGhagfbk2tKQNer7z2xqV6Br5FShF/e3uWCOC8yb+yWfnzWZ+xUYI
X0Gahtm8WenmsqOiToVcV52JEawkQiyZIwqKJ7hwkJlT7ywnogGAZLfStVHW3u8O6KN95PMzpZTj
+XK6j3i+rPOvQqcRgHI+6TugJKSy6Ud8ukArcLNfOStU88cyUL05qKBzzZGPpgs89DMnb7YcB61s
GZkE3+uMURHYxIvJkXE16kfVP1Zw+S1Mij1azTjXJtqKUzzlAMHi4qJ1qKKg4VT/CX5RFKG86+QZ
EZJx6KhiT0rs8yjKZH3Z5BgigaLrlL758rURHSpva7bW+kTNk8wTWE+Mdd5o0lk+0v5aUNEf+GHh
FfEJ/VPd21TUMBUhADVqqm6UVsnQaePncY9buODyFHJ8vOsciTLz6zq0hrvJGmJtNtP6MDEy+393
9hjbOUMRhP7dB3/mnUwZWbLbq2Ld7ncIVaHcrS2Wzxap8Yj2boG6Bxq+MVVQmHAPMGlelJAADPTj
MPjhOM4+03jimHCBweL/88No6U3mDjI7OIQx50o68xMDlN38eU71bTslzsqgc1Vt6TT4IonPJiDK
M+ViArAq7hWlPCx+XWLCGkXh8p3DAcbSHhfx0grL1g4j9iX8Z8VxlwMFgXdIfHZBOYxqmWn5j7Bc
xSdHMyp3ytfh/lZH33Lyg244wNTfSSW9C/X9K6+77Z9zNqaZbIR3wA/GcLXJQOhDPtJNiCkbqWi2
qsXmjlEOpK94IK08P/+NTRhqFho4hx60yMEoym/yoORFgBGoM9zQKZ8GDqfeW+Nf9zRVI6YoREor
N1RTrMkGf653urNtVJbbaiCiPvKW4Xjz9Zgedu1t03tQCyr6VItBXUEYOFKjG8IEh0Awc1f7CLlC
v6AfgTkAWz9r9KpMAahjEWxLsle8Qm5DVn4zpjWVC8xo4vcPy0DvmeLlfpqWoSH1JCiKi85NqtRb
fg0Vs7EWAweVip5dbUVhlbaPPD60Dxevv1Qy2PccNlSgKgiuAK7kdpkxrugtaj8Eqdqyel/WOmyW
qBsQ5s8SoXYJ5dBfENAt/iwtBm8rn06UT/fAg/4FXnJ1YPLhhjBqObQl3L06CErKc0QkkxlabdyQ
b0uynZ1F/SqM96xM+FaeKrA5dG16bMSttz1u7TnW270w/sVb0/a12z+nx4iIZwkoeZk+W3Gf7Kc5
1Rq0MBLc3qZ2bjq1LIzrlRpCWeO+OC33aUx/pWpa6SeVKZJhvhbGAp/WcyPqNcJxd5SXTSUjiVVf
hvHJ9lnS0FdF9MWQ309NEA94Nl6R9cwcDB9HFnAMAtFcTQqxTJItemNjqlpusf2gxJLJ9/wGvIQa
9W+5HPf8EhyRM1a3kpBYcDcIxf2Tg+XB5KJM6YI0SAFyDH5duoUDSVkEuS0DDjHNecRZD/uA0H1q
yfY847DmNffmLTq6l+OXyWeOK7Q3XC2gkSixdIhsLo4zS9vE/jWzTz0Y3j5EwZQjZynftPGjy9qJ
s+wwdYGjlLsr0aWLLSS/wLJ4+bj6QzlswsFKV0C0Aet063BlwIkcsCaNePBJdP19kgNIpySMJDh6
QtJHTlaV9oCOMmokb8vlSDPrmzZy09pkO9S7GIE2AhT/YoBfSqKyloVhs7hbTAQ4ldhb5hVXRHfa
whaW+QmYAVtmbx7Iscv3a9ozsqmFaEEz2Wc6DcflYpggFu2yCFFuq872IEyyaKiCE8pdoLUqoJC3
Fr9hcBVYt2/eah7r2rIlhq7NZFwY9mEAlwasIGUd0QcjrFV0afGCo7I7XM7WjFN4LlyS5fN4Zw4o
8S6fnpNKQl4IYj1sYcFoxBM7disQG5mDapqax4cXSRblIoQl+LdItzblrJL9mpjVQTKoKB5MLenY
/6IMJl+q0wmb4zhKS8pwyfQIfqEigFV1pko9DmpYJ8RnS6qWZ0rau76f2jBhw6rQv0kmhAuJ00MY
6nifVeJmqbnW90TanPMWzLTWxg3T2V4MhXClC/6GE+bJ3lwTC3hrcdbKJ6Pu/P8hU6bJx2BNzqrz
gCqMPjXo0nuCKDga08Mohle/MBl9qsuq+2lFJ4c7hoaPtFqPhsu7FaibNc3+QejZiuwZl6vxrLl8
JSmPdiWUdcEn0lsA3jNHKHtzExrxPVhxGPYayerufNVwGnACCv8ttP1VLmSt6aTnFOeGBiibqnCT
XWQSehg1syaOfuFjg/kSKxqHVMuFsnNoLJvgpHUH8vK+UeuML7k8nMYNX7dKFhShyrr1E0zBR+B7
+kzRMoFad9XiIqc+84bSBjBOmQjgnsU/7F6qTQESVky/KhOdF2v+cCG2T9afn8U7JjqcBnMf4HE7
+CV3JlhVgsncLGoxWBCZpzhfegLOEMss9ZgYAG4cgd52aMOx1re9skz8tan22vEYTms6Y1v/zQQg
EBXyqC+LNdyS18a2cLLJo09ePSJw9ZWdEf5SFj2SiwKQ7nClh3onLxSGYqmbBI4FYDpi/iqq7aci
/+04Y5yBBNWzaEHG6WsngkEL0SZJ5CGORqo2wc0yz0c/+SHVAvdmT9d175z/AV0ezhTWLMHs2CrC
Q48H+OyMa7rQizE1Xp/3n0k5EmKJGJLVKqke7MCeozvI8v2AXoy5rtL8VK+94j9tD+hoqSJfEXYM
PAWtRaRMlRUnFC71qAnDDXMcnOYU6ESSew3IB7P/fYWiBlI6km9Gq+DWcRFg+/l/IG2S5URwKxwU
RHtVbSAynYKKTCNa1xmmbNyzw8bTRqBYMHe9/ioUsX1es+lB7docXbIVmqzcJPRocGLzTBBcFaF5
FcoeDbJD0O3a+Rlx9LKce00+H8Noktt/Z+pOzYwI6T8KWNBOBt2sBR5uDlMhjuQjC4wzDbTJElje
VeJv8XL06gddx+Yfwt/dn66+ZZDIxNqoOasKp2+VRwBkaw8yVpJ2+fEkQoBUfYN+7D7vuzUeVg0N
+ClCWnAMkOGZOkovrNYAbJ/64gaoIcgNYACRjdCUXM5GEOaF7ZwdGTnn8JwUAkasniFCvG1cmF7U
vNio96bn7crQLx5MxCpi+j30YkeRfQRe7Y/0cBEsz4P5EfosnrmuPeeKTqhZrpDs2MqDUvuFhZCo
Ow+WhZYHyyQ/b0fNZleK5Gd1J4GARGFp/9BAj2BeGbKfD1hVX1ckT/LdyCPHrNKF3ySDSbgcPRDX
25KNVMPLxxwItjX6acuhiITnFwCBMP1cqs5DRtvaf7DGu5ykb3CYks6J+4Vz4IQ6x+nVIW6PqRKP
g8jXw3PpKHxPgAx29CrAjqgWzowsErSak1Dsh+3LqsX+sPjVC6V81EyMGvn/wkiPS4UVNn5xkjcS
EoSeBVxCkJTpgHX9EKJZRO9k55a7s0UDmXpZjdJWa8NskhQExDtHIze0xHUrSPzi3CV8FHaQMsw8
vFVNMylsiN7+ltarFJvFOjRfR1vF4tPt9ElSWqiUGTBD3F31Pf9x6KWwF+z+Ne+tYIz4aSYJz4bw
pns2r+QJhzPpGrJbV/6t6LWFxdH2KnZ6YrcUJlURMuJlVoGibzLXNFkeij7mLWAPBGWoMM3kQFxb
55Fg6mZEa+2ZmCLtlNwzDJVWYw25KVRerYegkH1Geu4um9keGXDkXfv9RGR4DcuLHz9G5ilrp/aI
2XYGbwk8+bUkO/bH/Uie6lET5UN7+rQgYFpjC2orl98U6/SS4BHyvR6UWNDM4G843aM+QsMpIN62
qe9dzevfz3lrR5+Az6m6DFhH+nVKwGhQ2VpGH/dCyd6T93LXQET7Z5PHly8iiOhBgU3fq0K2R3Iv
xORPrBQLQSdfYlYdvDXGSL0i+RxfYVVCbagGLA3PnuHH5TVlMxZHr1y5VT5J6R6/9f4Jh/G2zoJz
SafDJS8buVv7ILekB4KxXSd00jlTVVZLqUYdYsjD9NO82m3THLYCNw4M6rxngfowCnf4goaIZ02W
IV/Jcsu2ATIlRuYX2MUpN4gLWSvo9wUAl6hMBe9rBxBQgnERY4XMJwGd9GvnkbcUoyBpNi3GzKQl
PGcXOUM5lXRo79UBzF/hXkyluOFzufDQlY65uiS4sFjxCSgPDpLjUzZ6VETmmnNt8WOjpJkhZNDb
7lY9L/eaUhOKnJw7jcFh6RrdAOHwayyKV1c0kpwvYMPf/GdKJzdFp/FFWpsj0gPE4PjHBtNmJroq
TR2IDCrndg51p6/s+/U07qkuMk05jWHzNEWjDZ7zN6gBWS8Qz3oemddKa8sF7wgon8uo+ULPqTJr
Dnn7xvDnBXTA0DTfpr4xfBuPtOQ1e7dSp8pJhlZJ4Ex9PvKDTROp2me2SpDEK7mcP7f9bEkYcc+X
k6IR+zFyuAJmKICy36YIT9BhmUdepci3X0LBdWIz2KMLi9W+8KBsKAc3lc9+fCygP5DVKFIZnmuV
Rwl7TBRnXB2dyBU/8RUWmxD8sOjI32wDuoxmeT1gzk6IZcNnEn2TkjgLHss83PkAie87NOi5B4dN
ftdAlGsBOuByKEgrhBBoR3HAYKU7hbR4vUf3PZnTw2MZ0gTkiAhuZzWfzzsJuHs7yykMIOmxyFec
CPr76xXWwmuxfMZqZSMfnpVXJ+47rcJovzMMpsOOcY16MyJ3eC8Sz8vQxznOQr8zhwmhqIuCaHo0
vmc0tc0mo1COLD8dvYvpGe93NlfBYX+qpuEo3IYFNiCru7RMI5NVXDXgMLcKYzGnp/1zaVRq3LpJ
VP0K2gLF8ACooyFr4HliW6r5QSBiVyL3Ww6K2BdXEvj1172uqbsYMsZSXjFogJNwTp2uAeLJ3wXj
Gc47PeaS3fqaHgRnkqz33cLX6n3kcYPNFMA0edQAPg4/yidmlAIwht5xnYWS9/56478JTSWw2FId
Cm8N9dO2pmABjUCWwl7P9wnHpV4GGayCpjkfNzxsbvSiYPx1LPVxtrdA0ZA0Ce1cTlvhKvG0Vjph
sFltRz1FDi4gjt8q04qDQccoiJ9svZ0kVXZ0hTVMJvokot35lBdIRv4lwJh88/xGztJOGxZHPQsy
kybjyiDnTURWKKjXiKo0LI1c2Jxah+lfaH4qycrLddyZGYi8TJoDmiyB6qPydnvHo62+hasG/VIi
hVf2jW/yeatVGRtX5SRUJs9xSHQLQvKhaf5KQbY+XaYDss9gUkEQPs5oAuVBV9Qu2ZVu3GMPh9+3
GJfqZJbyOb7qlA2O0kNOMKceBpGnlJ3J7c9L9y5k88/JYClxSzL8+KemGwqP6aenC43pxkgIqIoT
WxfYwgJHC12uuD1DzrlBZBe9sE/BfOgFKIiKWIyM8vLBpl+1Bt7etm3QzDUhXIDLgb460VNnBb46
yqNrJtHI412/bPoQBkouaiKzPJdymgz6xX/8PUUKpqesnLwFTozHUwlo9Og5OdlvFPMJOdxHhQ7Z
xcq11i+jfv8MX5Uva7ynmIIE9FzRJJ184sHKh5ozwZ5xLubFyjCn/uppxuLKg1eKPluGpt1jFcN7
kxDFy30YkYzih8GH0Pd9gefPZC7MvFJdq8K9RJS96br8/oGGjDnX2Aug5Jmsas2CUfCPqDNZ1dp8
PqwFB28hzWOBC+79uTfdxpCSg5ichsQ9Thk5xxSfCS3mSVxZ1L8rRsktZQDFJestbTHDSCHxpeGk
Eqdr2uW8mXweVVfA0T+0PZT4G5Jr8HKxj+LKl6ALmYwJqNlwv5LuPr7wZEdvrmx3WJsbOt3XkZzH
8FSIjHkplfKOeuVeJ5DxGxiJI1UcTNCkyomFmQSexCreWOCwmATu+2qAKk4gzxmCj7sdZaTt30nQ
Vesx/YMjqbsnc1YhFa539p6/f/vXSICqi6MqXxv4DKxznG1lVUh7aeBnoq75yaJ/Dbde8NV/KEey
9zhIyTNaDAgad4fCFvcxqoD7kOH1G5bVmXoitFIbmX5GSv3umulwCzF1wvqvuqujxxoq34uLWX39
mj2hoPu3tfyQsT4CftPjzkK7ozgZwH05+qdC2j/kKXD3M5sL+ZrHCKdCalUbLTW8U5saKPBGBz7z
KEaRiEgCS3lOy56SnjTteXFNINbnEqesTJwgh1Q6YvhrBTY56sT0trYAUBZg2T1HBo66Ecb1cpxm
Mc+y+LN49rVQv0r5HC9VZ5ewEOjk2BTBIK+dHId4+j9JVUVPOfcw7uSrCvbD0/E5rXGsvMwtSeFg
vFxkUNneD/IkVg39A0GMAvEXa4qWYDMGV1ClM3BgsiY8mFMJT5ibrWHimQbdy0Gpgywo9KwtMxzF
K2NMnroDy8RGA+t4wXvfW+pRfzus2euZiTxqgvyqitEEdddUG5bozmaoWePPY2r/nU8wQzk4YqFj
LEQin//aDXo+t5VW6CPkfhaxtQsONaeAip67z4ZBqEPeIV5dJOI25dVxPQP0q6XGg78J9DiIZMkR
UFRreheN2OgcDvflGd2NA2K1FzKU83uhELVKSonkFQWZNoaoB6+mkj6H8v2LoztKRPRJ6W3ktOd0
eEqAe/xF/DWyqRPIjK2zWuhPK1EXAQAk0tHJJFeJEMv0CSYDrk+Q4inG4nR89G8Ip1qpcpdA6Rfk
/2Xn+NbNG6rssNbwikwE/LyXk1aBN5pM8m67eyVuudhu76ZnR8iK52NQmph7Z96xs6Io9rCopssJ
EskkkQcpFV0qxDiPm5iLlt+Tl3uNAnRRPyvJ3pNEFJ5KhmfEWCQCFeEao3deaatHgRVbmsyU+uVg
aBywZZthxZ0VfJk1RSnp7oWlVdJxife/j17tOlY/1uUMn6amFSp7VMsAP86/3SWKl2lLBuxmnJDF
/mtKkiolZRqxLGPUBPt/uTnBRpaX0EOELg1rVkXOTYbs5jQzD4hYkfo1MZPp5p/NEcj9tW/4p4Qc
PAJy1q910F546QvKLf/S6/hJIAZXUUXEcG6n4uCv/0Xl1QhdWHP1XZaURTWeTUzpE7ucwovCW4cO
+dpguhVI0zITBDtbQjs7lJR/5kylnWM0Z9lEq4k0vftsuCH5DEkQ1nyXuO/PHF2jfPtA8A4Ll7vs
RJyM/vB14FJBH57CE1gjknXA7UWpPBxfbgwt8VZGDJ/QAm0etSP4QD7yiO7huW0SOofCIENKxbw0
WcIEXHjq+if28ilTZCDRuWBCfTvsHApdXaM7RQW13+khzTPvvALmhnEXReHu9E1dGvrcrMf5oD/p
E1gRva+273CMBnDgSpCRkYM/TdCW7ul3AURR9ZfUioMi9DZcaeDuz+4LVgrXMtAmgG/T2Bi79gdC
NjX7xTxXArbhalvd+HF6Zn0Wvh3uFwC7f0UBLY5U+7S7C2NLEN3EwGBmQwEOXS6cshQXuDizMMhR
uwThlthYnRW054vE29/Tztxz8ZrxNqslqOvab5Y+9BVVF61g1frhxG6kl69ZiiorwcubDvxP1BaR
9xkJJxp4I0E+TUljuxMlJgvi4zsPpHsh/XpiBITbcfFWlLAPSX8+k4aYuoQdo3BFfApf45w9O7UF
56WjccjW8ui8256klmp3/+rSPC2xhln40Hue6Yz9lYyZEIWbU6P8Qtx62VsdTkXJCdvae7M7KSCI
ddJ5wWhSXHcjBLH/GCvo08k4c7g5PB0CZ4wevmRaYCJsTds4n9neOX9PbupJRDGTWqUj+mixJUbo
3MtAeW2p7XcfP6jDntVlIz+rPK0ao5+KAUTMS+LretfjYkVthYNMz//dbxAJwh0zDJCfyI1zv0oe
EZujjeAWSvHx5bO17KcP9GP8adsi8ETH9j7vf/XHUN6B/azQ6K39n5dYIUCjapVNo62IwyDHsQhI
UszT0kUy0ajZguxH9ZNOs0AFL+F/B8+SiWSBdnnN8V8vV0/xLXL/d2F2GkhI/bqsZKNMrDZkyMbd
/P2TrTorqozl2fnadAbxWUfoIORl7WLUclv29rJdzEmU3pFYPNODFKHBE3dCqGgH4eatGlQcqXWa
KTblgTbVSGXY82S7ROpLv/R0fwwnaUEqajQFvLb+vZgbBoNekJyvsPKa86QCILbtiJcMVtrYCAPQ
OKKnzN2EL0oftV9uzqotQl4x7sqK56n7J11cReusgMztysAvuSluzMfMGgWLhRAuM4Fa4Wy/0BzG
lHYefdDC6ZXpaLOMm5TaQqJ/S87Px0CY6dq7bqm5KmP2AULxwlZ7MSFWxJLhtDk/yToJNAhqAJC7
u/xxPhM2SURRDxJwJH9M+QRkcUlchVHxs4Pv508mmQ6J9PajvQPTXfF0p2kLqN43muxJ/CPXba2+
PQ/uVoWDd4/kY448rJGuTGagt3QyumQ1KfSMv0UKZWrTvTLXUZWD07qoNVGPZl86Wos9lUivYVS7
A4aLZZlU8EunKhN+cpSj1Cy0P8IJ0vJgIZ2zE+ExPiqDy3hk9FSnodvN4c1mYpH3R2RACyCIBQth
sk96D7LQee8vWsk7gibDv4FlGhlt2nN5HXpQRGDzvviSqL35uJumBajlhhfSD5tDkZGZ8BuO9m+L
6xPRWvCzOQnp3iv9LaNUkntiUyHtV5AYzRen7XNqltCxCw8KSugmy+44qwlEpFHQMXeAeK+ZK/Fo
e45XE0x2jawmLczI34wdSj03tnDpDAgW1mh0OVhVpJmX1qTSIXCoRI/vw5bYk+dPUbZ+QN8mBUln
PNLj7DX/kM1cRg1nZbWtMR/6H65+oxwHjtKi2JdwNoGa4mqKJj4uwol8fbCxz1jKqdMlvkknX+w5
aKzh2MUFC38Yn22QjzpA374In4Vq9kSgdPq95eBseGo65ziUHotvwad0uEsL/4b2BOBeTRmCTvJy
Xsn+tNHLFfSNocdVv4BUgSAe0kiANRjXcbpSblq+JHBpyiwhch38JMhGawcAockRapkpbtjjDBHF
w63vtg+OUgEiQWa+gpTRaTWLT15i2M4e1oRENlD/nS/XaS8KkRaJB7DXcgEExKK69MZ/wnlKQslv
+nJYpDuhgfIW8ZFNFQd8qm0JN2NUnGf8IqdQx2AgOMOEwB2488mQNGAtkY06pn2fmSO/KibGc4ZH
9z4AUIEhFIDUaP5hJXRtm1KYsbIbHYXkm2mYQX3bGx5zhTB50mYla/aPYjok2BjmmCIP/9nPYGDi
mWNUUTEoyOfgpnxjafguezvQuSJbVI12GcwGy3hLB/zizLwtuLIWLB76ZHyTNsUhmEepZXZWdv0U
6lyVxtjoXh5LCYw1WMu/FGvybfc3FktuepWpyNuSMEO/P3B+AXb1cPYzwcA6izy/NQ2L/SgPR7ro
+KtcwdqBuwziWwJ1zeiiNc0pQZCzCvarO6q7O3POgXEjKNsKOg7gUmhDva/4V8tNc5yUtMVQbI0G
pRW/scw89nXjqlhfBl0Yd1R9wKRiMmmzxQL5nDN/i7G72y+axJwXO/2kbtnYyM0l3USGhRH3WSj+
pjuxy27nTBNAE4Oadgp7/21ouioEZi4f7gzcFpo50xzoqSFCcY1uyYZ5mVqFFQf7RI/AQ6xR2Rmz
SLlm9hN094A9uxAOfWIjlbnMPhNocRw78romtpWqct6Jh0n7lIIBEZ1Sp8jXutrMAT6X7D2RjQxt
K0ekyga95iYd+JmHAQFu/MjW7dQ0AI0sqdiwNNmyOjn/jnLYSiCXKC6GISTeY2ynhJ/gJnvjLrAd
sRXxhpxDyONMk8c5acVNop9haj2sfvJiigsLAHawC0T9av9jofqxCfkH9t3hMA7PsK5YUljgdAJK
KiBs8/AjzIWYRMj0Jb2HfbF87PJqdRPA6Y/1OTm3drMZHvewRxWn/m66f06Ty3UXRu9RgxEWuYe/
U8AUCZ1HYo7eu9Rt5LGTgVEok7A76lXFlZ2vSF5Uk9LSBTh3G8sqsStvPBfBH8yfLP2Z1Oh2sbGs
C54SVYb0GdgZo86sU1OzFNvPlDn4frGOdN3BbuOAsN68/3cgNTJUO7szfmGnPXWzvXdVSUpgQSbO
vAOG4+tWvINurIXNRCf10ic/QTz3RU4wOmeqAM/IjT3+RD+qlunPMNaMJunT4gfKKZIPm2e+eEak
Czc3lH6WqEsiWSWruqyFtVRH17OFpDueZrdeRVLsKCQQaW/X5Gs7mmDTcA6Fo2AL0+eatvOwvnbm
XYFQ/4PX5iYygEEam5lqYyt1tXu7fT8rKlW45wWSphlJu0uCiSOb2daMMEXHFazdF2b8ZxfTr9+T
z9VB4EccWJLWpoSwZjfhG9b3ev2ARrAnOsV9J7buO3YzYuS/u8PySMLdzFxk9j4vlaZnrIH9i3/5
ipxAQhD0iXuI1DUjTvhdDIhKqG5gSutv25/ItYG3QadAySwEtcvPtlEIaa9NzUL/ClgYJuPWsbLo
jHmzspcJnFkyIZTThlWP6g01alQy2ROo8pGHBMqzLfd3Q+yWhWMS2IZ6VBmEdgouCDI9AaEyGDP7
313AdrKrW+yc5mZPN+kt9CEFyZoRED8SPGhGl+aJbhylYtnVkxwNT3HV/sFMpoJ2ZPkch2s9rt02
BJYm241DSOoN/RjD29Rc+p2eoxswn94/+RFvZ0o803IkN69+k6T4DJcLB9wCUFrvuIwvvOu6veGq
WDA3+LN75XjZDPVC96jR4UT7zHqCsJNqV/b6x3EGfebb/+dF1ZVTSP9IegH3Y4PxsdNv6b58j+K3
xidVXrT7LFojGA5GppkJN3xvXHyDNfZmiXfDvMokg7nFGvW0xFA/PUIvS3+u1Pg8GBTksp04Pg11
zaDdtmgK3XyQf7QxEx7Q8+SVSOyTuUhlPYwQ+tum24ISC6tTRurIPdVOEOhSXzpY/UT1NCcIcrSw
Vu+OBAq5yGMwXoC2kuKcm0E6fz6ccGk8DU9i7TQq2+TC5cfjffXrrdikqZsZcquJ3thM4SWYzJrm
MqZRPVU/43wf2L87OJSMZP7M/JNyHX5ZLPrrGiwpqkvzGtpBvcEF3v5cgwQcy7cOUopExrvIb7TW
gym1cIuDR56NTctOwYNIVFGabWUEnWWtlkyyYFUNNP2tEDrQncAzBwJnBs6dHEzVoIYFouVGXXih
y87igKN9WWWl7sqLp1FH9bZIWYhxYe8BETFSep9wTwLj4cl1uUPGAURXZFgUeXk1d7si9bQ72Yuh
v+fCf2fU1LmdTLuMhwDmE/MG7JskOlJfdjJ00dWZWBC/Eje9md88ZWiwEZV1WfoWBRLJQ04LPtVS
m882liDvirb+ddPBL1hsUFZUv8fJSlQOMzJHRrSwpih3hBIhSEiKSSDhUfMc+Um7AoYcSD5nOUOJ
Rn2sL+MUhlkQld36FeDEkeQ1izxLkkdTuhkwkDLRuJLDsTRFYxO/7pslsa34n1kk/tfybfsByn0E
UqCEcDwNJTea61VTTwDv0WRYH9XIMAwuazjEKkf002T9ovR3GPzOaF+aR0w6RuiLkdnBLVXSGIO4
8NPjyuWSFdhaL5D6kwnAH5cLb2qk/VzNp3jcV5QRy6xp0kFW/kR/GzihLeuuP62HEwz2b8E4p9+K
LzBy07oAoVqHxGyKjAOgM6n1TK2lXsLHikWpMnG8D0FcGu/IETDqfxZEi/hhhqpSxp3agCx1kM57
VkGiWR3Zm4vEdn96oJThnwtG1vNEeLC85kTclB7ikgsavB1D6ChbUc64yXx6rgj3qt70M3A+qXn0
0Jn5OBM+YqrNuEy3wnnJrnneAci2VuqWLMrLouuejs3AWGUoySGnszI6S2QonhS4QQVHXLhJ4Rpq
M0CKlBXsfqKXnF6WE98ThJY6PS46AHxZ+F5WWeocnlp/GHz1p87l47jQ4TjoYkWfyy3QxQUh2cqT
R02Wp3O3Ef6FlpQ9trPMOPNBYaug5SSK729q+JmPfzguXW7g/kw+zYY2dpOhZa/UYVtt5Kx7xz7L
y++5zprJj5SiXavQTKMuv1vh3T+SUHQjXEf5fMZ/nskhj4IYpFZ4oDnN59rpkKgDBViivczj+1p7
gfMxoiFeoSiYKmcD8gOQpjVGZmC7fyPHJxV4WAbGPwjjid835zF54ThfSnrSVeUUPmi6zkYX/MAW
UuBR6sscbUxVu+33xgnqnNAPG3SAF0aFaXFREfbxtm9yjmglfRaOc6oOSQ4bTqhWEZv1X9h7jzr+
64j4i1NOlNVXhIpZFTXkztbeYJhzIdG8Vv9SVKJCZmtK5AXHa9e+LWpOW0KNy3H3FgPvo0GYCdNQ
cuwD8B68kcWuAKBfaGt5H9x0PET7qg7xz8L17XYE3RjSBz+aJqeCQhMUa5A99COo3edJrqC5q1qu
c5hoMN/HfZrrD/XfJB18PMMA9gGxsXSU0+73983N1pdL2VtfEoPTSFP5OJfuhUOEaRkhe8/pmVn7
BgeLu90tFGwTJfIphaCSqeSJDspXcwXGpKLF7juaYV6PheS64GW4x/FafS7jnv4beG+Nr4u+4hKh
thkY8tOdAuhNi/f/QCVJ3Q7/MPHTVzCdNTJBt2VcSzoYbuyWiNQkekuNFUVIfGMVEnBG6+6jKz6+
kATsEce5GoCJFe3wt9Hib9h9wMhaKCPHbLdXBeMktWeMvALXXE4V9aYRNuGP0cG7rmSwzUrLOP+C
Huu7gK1VjO2imMpmMGzjv5+Skb3eSnS1wAo747b0OFf8SA7wuUIfrEAmFrchx8TQye6PXk8qKo4F
Rg1bzua1WfgjPTkDCjBUCihML7YevIv/YJIB+zjov1mUQNCV8SJjgnyg6aMSVHA+IGfMNnSoiQX1
aNrvfYLGOjoRwQ5eq2bBQ9KdVeav5lgK1SCCcXjtsVPl0W4Xs4UDIneE/iMv5Qykfu178S3z5mQY
HjEdWvAHZKaupfVxb7AFm2bowg7gsIdhjZCJPkwKnu+xdaqUNSJp6PlUpXmaaqsHiE5D57CPZfXW
v/l2/hfQuYhcBUwVAOL/QnG/loPY2D71OiQRnpD2KBsftZlAFTbJR1uQnsbjlCQuOfqGo2RA6UBD
lWpvkT5qd/LzX3EtdIu7zv7qbJ+llXhLuUFBxTF5zoYWr5C4Db1xHDP1Q+vII9AmjVAT0H7k25fk
QlKcSQTzWtn7gX2w1IiuWamEAmtU+Bq0EBu3mIyz87exQS6I3pitqEfB8Yjb+COa/K3kILT43wVI
Mjc8WEalVUnvEKRL0EapIvY61ErEe81ktILbfqhm2fFW30pqGFAMu0q4gCmA8dDVR41bWI5q3z3/
VfwHhHLBiz3j9lruC0R9FCHAvbJMxEVNtEoTa8Dlb1kLoew/en6ufXQEDXE+5furVDOEOo0eZshq
Iqfodns7UKEQg9beDQAnaA1MJ5MxehJSuP1x/EVzvSpdzEABJnsYWqWIDHvpsltP7j8awNVKBJep
8o0dmKp8rfNNjthDzkLMYXRwlr7YprAakJNdgNFRVQEM7I9Xs79fW57/7KeRsrqTECe41Qnf9inL
BhfiyXKZovSst3qax3+iofkOFZrhvVgdxB1JdZUQ5gkOFQgDJIU4u6GU3xFaxYBTpRmwWfwOzz4/
jNKwsp17rcNqwl+QMtLHJI0xNInzwKbhvTj/zHuAdKQet75X8evHWJAJcigjzHW7yqVKNl/o14x0
Uwh0CmZQjQUVZJP06hkH0hT4ezjeiGM7senXLkcQNGxEZtbvGCtB5BBB+KKAQ2yNITz0kbRGcDbK
YquYz9abxmf+BmGuEt+y/Kl1ZaS/SQWWBg1XE1pZn9i7S5rW+Ofrds6ijDI02vnHhqIt+Ce698ka
Eyej+xVh/e8i9TH38Dj65z8kqQp16lHrEPCWTMm4AQ8Tk7Y/6RuFytV9xUymlZN6Md/9gWfeRvN5
d/DqwcORGklsjYPuRVpp0AQRVDmUpBVQ9rro9wK/XctY+RokTmOeUlKBUEE/6ODeud23b4Z2Jl+5
hBYMRrpsdNw5IPoX+xoy+funEBX39uvadSj1PFkEnfcd5sG0hxBSA47bDJCvJf8bpyrybOiFJRyB
27T12c/FdjPUw3Hf43Lz7+u4suROjX6H9Ew++IC8oLoIYURn8xlsvxIGPUp+QagiWreggBEEW+xu
gXO21AOQuuG6TUEzMN23aC/8ut79XWWrr5b8FbGkZGNqhMTqHNjrnjqVZgli9Nh6DgrqD0iTn4vI
avvxx9Hrf8qMvaQ1bH5A337HFhcF+eQA3cWsaSV7VMRDoUrl9Q6kCjosa2FjipAhm8Y/7jt35/pr
fVWsIJ7AYNIqchWfuK6dUyT4jg2ciQYCuJU8ypHIrydhH2LvJmn+YnuyCgrkEBKJ55ikGqo3c7cG
dQv2fR7pZly/6V6Gzg9UALoo8cI71XDTAQN+3C9YIYOwgWeHlpGbnJgqB/E2kLpxDSJtNgzrKfuQ
B3Pr50Cg8rxkuOkY9wDJqSZNN108djIlHLmTTwbaJdRN1OAgiUQR//ezy81kIAWHc1EFvg5C4cNu
QhYHfUZe2V7fmqZ8erDVqZWkpxDGnKqYjD3cksuXcGUcJQxjZj4XUol/PkWmiKppStI1SMBqNExK
R/YvxAzsqf8nZ2y/PeaTbg+Q5a5soPJTUPn59r+ojdQys48NGgtZNXmka+3hzYCZPxOu58ktNsU7
67Gee9ZQjlMO+hRLCxvRqxIcJsiHsKeNUpGUmGQZj7GtuZ4IbvxRDjwmKKTUEV5yB+RfzZ80Uong
oBPzZJc3mix3o8Ts/cjtNqXNttuGurPCpe5JkIqqBUgH1AcT5ocxxuCt0nC8ERjLMnH20vnx8S8r
ApZ2GklL+evDQMPTb8ckWLHFgHe1xcZFRJu3LDfTiJ7pE5zgtKaf1KYp26RLGWiMQzhQpoQr3d/7
gE4rjL1v3VFaFZVhD9sxpiKcUoSVxPFcw22Dcuj3sn67Yhv0XW/kgN5MwU2VpEJTjWzAO+y8s/P0
Y/cqAUpt6b/LbGXfCQjZFjUt61qFOKhlIGKHYGv7iBF+TURMhg0XHRGjcG6qbbyI2Hf8EomXSgop
gzjKj0vXCYvFgchcFkLdSskc94h2x/kG7ODt+voL/uQE9EpQDr8lfNdd6C3b+l3VGLBQbCyHMfae
9GDNaEIf+luGmsDrrJbNQtnnTkS4Fae90meTn7Cor//Wa196t9BczozVoTlO13Ts/S7pLuL564zJ
CZ9AwrMebIZf0Q5dX2uQxviAm8DMuwFvp2byXioCEvRTISO+lJ2mNogiW4RMEOb1UcHih+BoJNHu
iBDeajFT/NPxKtdEjqkra1k3xRIntzopP+o3Sn26OAUkHjgPAya03t9w/fX/Sbyzsq9QqxTx60DR
rIwI2lCcl1L3BvDaM4fN90X3VqwCuNOiz2hIh0R5Y7UrrWkic+O6b+tuzfjFuuoCHXXrB48J4EuC
+2VO9vil1js5puSRKvuT8qg25rn6iaisPPUGpNf681YZmwP1h1VRGZ2c4KNGW//J3LYoCNwDIZFm
zbv/r3rjY1T7AmGb/GeaCzI4AXNBF6mN3did+BS6jernYRyM8KFM5WkipVf50ZDkTEdu7+uGt069
Zb2DBBJ1fj++bZc4j8BQaV/cWZ09eUxKoCO0XDNk+Jv6/7OJK09V+2uJhrSxiu6Ao99qHQTJEOpf
fKsXar2dIrqnKx3546QWzSG/RieL1ThvnbuR64AQX/fDt7tRFV6fRcSuPTa71Eh9qj3vhyS1mTkO
OkjkdJmNRfF4rtnpl2/iYYuGaouHrFMhlGLBwV3f0Yg2HWE9GgxIKSCzN4TgFZQZ2fUbI11QYPEc
xuOH8awTfHiOr5JPV9B16elJp6Hff5Kfw/UQ7ZVi5kuhn+OrdsvTcDfO7H/w90ycG7emYQ9DRcof
4buNQ7pVpT+eg2P+XVNGOoRJ1Z1KKwtUOU9+QeTiZ2zG5fgMR0TpFuM9fuoIpYkaf8PaA2mEJKAa
2zl4URS88/fhwZwwRifsTzeABXQKt5im4ao2orhB9YVKFufqRdcMOs6Hu9dxLRQcNJgXeQehvkY+
Acp4eL0GhJdftm6XD/7p8AslyAjt8THkK6cw5GwrgScB34BZOBpgqVK6sCfiLcpsYMoZK2mBBEYa
WArDb3p/7gBIlpQoNviC4fuPvx8QM+IjuPB0PnGrmMs1ZVEJ3b7sC2cY9ogVkfvs42VZ6BQeebZB
EleXOOCq1EmBbXfvcHu67K1QCipfC1c3jYC/neTGEaH5cmZllWqNWx7EDwq6bun8xJcQPxyMul+u
X6doNbl6/+ouRQc/dsgZA1qBm/b4/Dqgzt12Ufp7QGOHC0dQ9AsZ8Gl9HXDueAalTrv45NVatnYi
u772uW79KIVVY8hd7BeR9YGuchh9jNzRO4Z1HEmc2W1Q8q4HYKvtXPhXr9Wjrttum4iE70Ijk8cB
QtaM+fiVtsYiNHUJ37yMa1nlmDq+S/+kcQHnyilWFJ4FhrD/PzAwwLB6/3GzQlIFiN1CFyMS54IU
ga6/4+DK1qbXS2p0+Ljgxc9/64jsR2OXHfsZij7C+o03GP2Si4+f1PdA0pmfDqATP1Zb9gnvBD+O
eW+yp5lNd3Zpy67GqiQyj2DCQgiXksrvWwWy2NN4braX6bir9dAP2Gu2dx6UcKjfs9u2qH7madgE
I3pTMZQ6Pq3gEJQAw+ll5VxBUmPEhSOmJJVtPN3urRu6D9pMbkxnklcmNqtDQaJm8Joc/X1oKamf
xMy1ggg446u3hCIqqt5Nav17tPC+0AURFgEo1lSr1BgiDTMr8YhqugawQ1zZrtOa5SyF0JaOtzQl
9tX54cgOA+dVx9Qea957jd/5lHY569nOqQ1FwzFsXXjHRRkwN+kHRH4InLAq9D5Lj3a5vZBSlCSs
YTUMSAtCPSP0+2X70rEkltFUE2yFSpJ6YkwO/aa7BpoQ+4oWuGcw4cPFHY67JlUGw05S8aJHvu56
u14UK8OZ4kya7eqMg7tGkCKSRiJaZmNFiq6cWKNd8Ox/7pJ6e1TnKvAoSITVfIWnnNN/GTEllMTc
/sBRfMfPL9xrFnsmhvaRU/D6nKnzfAzXrI7i+Kp0V+aZe+ZFQrZft3bbGPccKxApBTSsztX4fahD
mQuki3BO0jeogStWvFx4yzfN09MHJV0+nY2zm21ApBScK+dT6CqWe39z6kBXKqPzzeyG0Fe6yWrX
v8bze0u0R4NA/v4/vyS6X0KvbbIYLlv2me5TPCtAin5gtANb1x+gPtmFFcw21rUNFKqj0IheNLpv
mU3a0ZGNegKf5O8xWNwojUmrEeSnVxIaMigDdd5WDjc8qJiKRDCXDz07AcTTjgz1Lb8etExzMSMP
+1ie73m4gBopEpzkipPuY8NbPN4myyF3YRoS1X/GCsLaJjwBjbJxUJG6XuF+iYJ7LLilepY+sGNc
x2l7dp33vcQJIR9ZETQcPUdDbPOv4UrcoVuphU4GNKDRksZdoODkizHdtyzNXDSCG3sUsfK6csOW
l+k0OwZfqSoVSVkKozt0jndI3Emh8hXqqrzbMkw+G9rr3qsiIEbCJOZYmYcyykr2/E5WD7M/EhMw
cgjC5ADJzEqfeH+T8hw2O8LmzA9f78O9Ewls2FOl19P365Nk2H0rMv6QRYwi5HTuC9eUcDyuXbLM
RfKN7F447oKohiXKPVC8qiFsl5DOxdQmQw8XoDs2ZwAA4TAlQz2xbZQm8cZlzu/fXxacMW/3Wn5V
fJrtPRG4vFB2yCTK8+mx9WfgHW7PIaAGA0H68WEOXWMYo8hZH9qpvjcw5Gc1HugfMs/0PTBXWn8U
9VVTq4czI3qd0hYQrqMIyhIYFzB+mA26PQZXCh+l/43K+bQ42k6PU+FrAEOjYmFryMvp5p9eyb3w
uWwSeK25knKZkLTvJn0pehNqWt60nqfOEMQoDJsJcBTvHwJiUJIWhqYojsjjR89moQdMpaMwBTK2
xIvChVGAj2sXdqkBc2gz0yzh6tq09pnNApW0w9P0/N9GnbKS5McZrZN7bK0My1UFTNP5kiLMK0qs
kW4wT0dESCrNv2l5mkrMEI0DUn3zGa4+KrG06XVeFu9I+/3gc5MH+w2gRIKjJeBwebIG+fUXX4dp
wPhBj+Zf0fa0yyw11E22xAqZnnKz9Vl9rrjoEwfkRlCuEtxLYJwg+50QD6Hp8v9NNJ+daaA0MP2L
JVbZgUhtQErl/QTX/oM0zxislQty4hdv7M78MT1ApBUQidUWut3jMQKJWycbqZr5g2M+RQs0JrRC
050jKO0N3TJHswzedTz0i+7CppD90akBQho51j027gZWfaVZKdVtQR7W9rrPKyci2kfDEmNKZFBq
DAGRWRh67fpysZ/TyQ7bD1FAANkDWv6WMRZ2ctus/mTVKNc2N34f2P0ml6Zk9pjddsb8nLDQ3O0d
+kF5nV5YXXMdt71plU8MI31w87ck84FX2GAB+nTt5FkbxAgocOZLvC6cNhIzHXM6hRtR84AtDbFd
J4rLm5ZVPrEubmscLoFCARnWXOdTTCrN0XSEWdY7UaRttkSoEXvOeDLo3Fcqa/+zB0DMzt07lsxd
RAMMugxZ1FN0YOcSIiMIZ1bAzGW4Sist3eNiq5zof8HdXNdjT4drQeNqumGNd6jZ67O/WqZhy21R
DTpNkpeZNILmcmQbuAm9e3VA3S2fjDuUJUpkypwC2/qlwSp1nslSCP4x3eIcW1slHD+zk4P76Ql8
+7kGpMc37o5sleUZ7GXrxGFStcP0yyIbq/r6hjq0E0ZcUnk6baQ7VDsNiz1Cf/mGAgpuh41aj2n4
1oqQ0JyRnkH6GXxJJZKYaQGM/ZXqBthyPPAyMBG3sTrbpQFwk6IR5s3P9Lr9yAa8AHpxqtWLpoNy
QMa60HOl48WC9mADlJ6E59dIdA5+vM2W7Kaefqpum7Wg7x0PzTA7Q/1gNtrn+twJIJfqXNzp6XMn
GqFHRODRzjvT9hl+woXXYqZXMBmhyQYIQ9AGFu+5yIewtanKIpAmhu1h0Ox1ZsdRhYLs9cU3TP2t
ODYxWgIVtOHtb28TVBY069TBv7Znl8wZ+EFqSzfG6hkNfjRXmVd/STf0M3SNVE3ajihulvAYzMNe
KOsLBh8SWnCT4SYfvdGhZgyvwEWn1BcDnVN5RkgKFvPCQ9vD+Oqq8kBFRoqVQP1qzujjZjg37Rzv
285x+ajjzph6e8KCbuCmJP8EVpnqK92Hxx78sV8GfFwsfI2o0CGjeJa0g8jKTNVreFP/XjRyBOzn
54uRXnCf0JrFpZyeQORBIZE1XB1jWT+F9E87SUslycwixRyQksZr5Rnt1xBJeMRy6DR0TIqohT4b
Lqa6s5PZkn4L6OSY1voAtKDqrDD5FyINKdVZtCHC6ZyAhdJqqGE9yl37Jbj18lWGbRJDd0CLzhZX
lnsf0jvm55uExa0GnfU5QxR+nFgFyHddLaWYtqRAEeifFtWaYutPlW6oE3ynzwtRHUs3dR8FHh2U
QP285dBquRokVi49voG+VomAttfFDB/2HTcNDMvnhI9PmUAaYM+MZS0vRHZk9TOSm/VfaP4FeeCL
2kA7/AvmAhytAyAYVcgy3G4zlaVvVmSEh49UfGIh7EKe8IW3pnLZEGq3rjW20AbrFGv4aSO1MoGz
c182QpUYTVWNb2WB77b0foGMoRCViseDIzadHbQGkMP0+FczLQae3cbj+E1tg4z7aIG8HO40RKL2
f+W0qPL50XyZK3NTc3+o61bsEAdjagvagal04R6XpEZbUY2V2ZM0TLU8Ho7yBDH1m1sV60oImxxY
p3ZQrO9AFYlhQcAmfhbutJW7npkFtbP6+96AFDenMVV5B0z2r+LeF7trwmmooZ2esWhkdA9dhu5R
PrLe5+hWQ/45o/K0RbJyHPPhptxYHgARQGKW77z0GprQvJ7aOE1uvuJ1aXKXfQHPxrMTNhcV9g3f
CY1IE4QmXdx4YNEqWj9LGSfbxt5whzcXvi2ax6ps2tpFq+xQVJPT4+Dc74a0NlSXt21RrJa7LDg/
89qGn+Cyy5M2CkDkWqbX/Ht9N2Dc3oyUNt6Dtm6UAXZUFXamGHkTAO2B2GjBUoK6RfP7kYyefOFD
aJORweyf7iqk4ecXx6xId0S4vEoTCRyx7rvAJ/i0fUVfIXq1PjvWg/AMF9S6cxUKAeQM+KuL+YpM
LrSE7hwSseCrjMH/qfWRqa9p9/7rkkmwuwtF3ETMdaKXBln/VzBZm6ZrZ75gpdI+Tk5o9ASq2LB5
zHID3RG5FfAt1sg2PxmO2o1G37QdXy78uU1gtqYZ9X4F86Fk5ahjOKsUNc3Nnz+acR96ISf9YTx2
Q9bmjVJd8N5TLVTjWC7kOwUNKPeB1kMpj37nOhx6KT6BfV5RH6VZVRvo9fqv9Ax6HNWC+56EvJmU
xDk2dJ/qvCSZGtd8TvpKbcjdXu4bTt1oqSmssMUuQ4e54wpTiE7rOpjL6oKRJd2xEKa10zhPmFNt
Pz4bguFGEiDMnh2jyx4O3aI+9hE7njmjkMiFEDa72VSkJ04V4Aa4c1E2BBAKW4XCPFRLwscSzDDd
cwLqITv4zhyZiO8niM9VBfIIIjOQ0jtlM7C7T3q0W1VEGgIOSw5OR3495XpwoWE4YRxFWccvM1Km
ZauPQkJ2Ndd9GenSuZZXzcSI4T4OBkcsS3Ture/6cshEaWrk9D+v2Tqx1uYh319kJQxOBqQ6tAMs
wn6pixyIJ0E87S53giUIJ4GzkAbnEvTTu4V/8585UXTBdH06x2JPGNwJ0aMH3+iTQQmWKf6ar3sN
fhU6KjtXRprSUL0hWnsLJlmRNjpx8/h8iGdUZ8nddc9omftQnENLzKHYeyZfhjDia8Jjt5yFWLDa
wh3gy+TNfjH+dMEomK/ERxw0ljUB3M9saLLZB+PP/OT80kc/NEbtfhl4tgCQlzCoy3CHlkR5tyaf
vu+6B7yjWdMeJO8TXgQhH0R/GOPjYor2NySwAxMy3Dqk6aJnm+kGlzsBj6stjgcUvJ7V4F3UPu64
fqC5WkkomdrCN7ZuaGMfGtMcj1gMU1Oc6dTAiOkMsjR0JaA3T2rjoR93Oo54xE9pWU0XpnicmgwY
0xTY4qPHCsDoIBNRVn+uCHdPJVpYZLSzOSpipbNJW0d68hEix7HTZUMWdafLjZ2kczC3sdGaj1XD
jgyQXZ8GitxUozMjoRDX1xFVoIJmCuVPfL9s+UtoWUhlsib4fQu5uGv8Y7cevtex2dtLJ4LtMwUx
82QRV956oOu6MdOggvI1e6Zj2IBjIoBmIkvtC/y2NkRXwrOXA3IMEJ/ORHBVxQjwrdX+oHxz6x8e
kJGt7ukAfKB3QUxlhiAhXjs4EB8gCFJR6YWuRAS8ElCftqdr4K1qGnUxmvU9a7A1t8PBUI/QXphx
ZNIQAtQGxZSkYoGoSI2WWZKICXnmCIi1EwvbohipmazTSubsWx8MFeAdLCCqtcxCPMX9Xs1dX4bs
IPSYtykSAzrwWiPPXFCi3yt19S4xhU0U+D2xCmkf/EbpF/6hKtgNVbf2w5va52cHj+r+diLi21Kb
OqpimHolq7v1UivTqbg62SAPXv5IbHNusxYQxcUZYG6dWlzn7p+w/50IRsx5H48BZ95VYu7xvt6A
7UnVwKKScD66tSxucs3cs90eZ7Y94pGKoPSSNK/aBcgnEBQ7Jww6tTotzAPxiFW20rP705poxaRW
0zExkrvTrtKcI/7Q4PYatPkH696qTh5a3YPlxRGIzkc/u+qcPQkMNG+OUjumN+Cv8gvGz1UFPrx1
0MdSS3llH4ClyRsuQ+GyZC83seIa4gcvgziapVAELSO3ahbc0uEW9kkKfJJhuR9RWLd+q8g9FGhS
I+zR/F72TDSAzvdmPYY/8eVYNoCqi3gyCXrXthNcPp85VNcRjtXdAXWetduo9vGKylq8ZWTdVjD0
bKp9gZGs5yyn9ieIf76CSTSdl1jAdv2szG0r94pX4F4XMFk044PCQsclwHZOQnnyedZE42+d5vvg
hNaAZLs78G8gxKXaRyoMUpTu5Ig2LE/xNxnoRln8cueSkVNnBc4Pd3qW1/oks0joCxsYHxH+a0DL
QQpJ25fuHK2TICBjOAWKZ1JLR1r2SDsUKfXV+SrI3ZX1PKSWoDr1ADn/CU2PAVQRw9763s2Xm5Ev
dp51wckT9Cq5a6Fb3vy7acVwh5N9yGcWxv2Vr/Jrpzh/sx+fTTIIrdrBEf0PCiSY/Mt1GMZxDI9q
m/8liTclvWXmApWNybDgzmz4s2vJSN79hDvqRnJkb2Zueu0Fql/rCkGH0zfPsB5jwc766+vpg0QB
z1vuHxmmPdMnWG1L2KH6MnMtXbLAC+7/DTuGBpS8cdDrJEZblo2ADSAXYwzKvwjNXjZhoD4cwXqz
bD8zGiVV+FjDUG34Jx+WlBrYbF/ybMVS+LLJt5aPifzhyfNzDUTxSlZM/wejUgxEgk/K1VEg5VHA
cfW8yLJygA9ReXwuTmp5pwIIx8fbG0FBbvd2/VTyl5n58OX/XNnFh9tO7MlWvqRRX83jpVRG/2s4
F5jcsTl0ev8WYx4uNiwBrN7nQSs+xHS1/9kcu4hMZhHMLaPRWIH08SYzBLBN+YNfWDcLU4k6uJAK
LxNXQstE5AhzAus7/4mojTvRqfZUd6nTCFtDIst90xFHcr3RTMe/pvN8gM1CeHV6s036jqG0cssL
dYUi3wVxnQk0qkC19neMq+yDLjHy9dTJ/VAp6y16OUhZUdQMFURtXaVGdecHJXL0ebmuv0qF4H4C
mfRWw4bTE9Oz3uijhLQNQ+MiXBZmdmtvqni7AHVWz6+4vZILoCyLN5fZyqvxrccyqpIDOf+fmNje
56w30bxYb+cMgjpicWKGaw+u5xavk27Y/DUd2nqhG+oVTOru33PJHc4Du7cXrjuJEr77Z/6pH+jb
fjsU+mLrlt9YD38cUmqA0czXu8HF/Zeh7meFWm/iWTMBVX+Zp2czSOG4+K/ixHApCPP4pPb10MY8
xJNM7GZdqUKX941c4s/XMEFLBjKTEnQHSqoetIKQ4Q4xAHHDKpouvfeOODwViNa3eJVNQ5Zr3clA
EtfVRYPkuJVpN+zA8pu3al8Q1wS0MXnqvUOpOjoeIjnjZac0p5BiexpDVQUfCSqHbuhZgOlUOk60
AsQrza5CX2JQ473GJtlETb8bNZRVCVXPs0kwG0Ef3tQAp7o5cCW/C06I2vPhMVMsggG5mvdsvfMQ
xXJhR0LLk3Cu5wShZsmitE4L58azzd3X0kmvsO3KUBnUx78XC4GaEqT1vrX4KiWq+ghamwRGAn00
XeWYaGoPYoGLdHbhgYgEJAwpBW4QiC+jJ3+ObBc1LNqRKnY9yea07LpiK5g8bmgJ75k6UxXXCZds
ttgRUFZOkoQFgJMBmFbz6U5ZMMIQ6J6/n9Va4Nb5AGiouX+2ttd6t2W9i/l82or0nU8rMN8gqrgo
QjrwR2P9Dvws3BktG0Ze3X2MhB3nU+pYtywCpFEsuKgWaPlflL14wBMtzN04aXwvduLj50P1YTNP
9Ofa90Y6TDF8sDaY55L3Aip9sEEJRQ/GjMsnuAKkT+zNEhmEfkZjPIlxlgJ1vHTdHyfdTmi1Qtw7
P19hx+pXAuWZN9guBFkWYuGYFK/gJgz8+H16XcqB5pqV+IFKlvAT8z/A87PA4uVlZCfKCSXhrPa2
F4pqTRIKwrT13Lslg1l20f3mtnDtG/WYxb3/nrD/Ub4WFONoIMHe5roM1bsgIbO9JQBc8w+e/fG8
3mPxIN05G6Un7SvelbGPUAon7ivGh1Y7+ZZRZyY6T6u/qsqor/2iz/x9sADQ4JYzNzp4JVdUEJID
1Asgz5s2j7F4l6qjbWj2zlkE62IRPV/2aF62dZ69UiWp/TYiC/u+ZAKFSKL6UOyIAgOsSnA3pu+8
QVyc7Hd6P/4UO0iLddKFoYXz2/4zEb0dh6Os/Jjly0SigEFQqB9r4Oup7kMEtxjbNlgWODxnxVyh
U+NazWhqXjFEnS11mMKa23BqKvsPe4VlBxZdENKc5wQ4RGPwKqIgK0U7O9XaVweZRqdSZryC+X8+
SPE5Mmv2pmX3p3ckAqmpvOlJJ7F5gWrmgBTl0ZUxXAmoGEwxp8Iq/g7b4phpip5iywTn0PBj9fer
wYuXrSX9pGytFdJju+SIIGckFE4ACsTMKJ1dffU+VGV0hDfSLT059iFKUQEi4wOrG0Nx/sbFawPl
38aIcPqPULJNO6cUXGiasJw1k0i93bOMuUz+HKKpENyRMzlUf1ij8azhf7eYdg2m43lcz+VHxL3K
/3o7VQttegDKGfn+0rNZvBvr9bo+0MJaYy8UzMjE4SA+5Nfnh+OhufB6DQKV4fRvClCA2/QTnUET
KV6M39/KkPjd/DQMigkHJzJBAd9zhIQZF1hnpJQFpOrzcnaALiHcWt13X5Xz0uz2Y9IdqVTS3LfY
8wFmUh/IIvtbYTZISvC+i/ilJ2//qmztk08osyK2KMhYKaN+gX68SWFvq+todMtGYKQg/Oh52eo7
MYPqrsGcxZHNfnRv7tJjK5UB0GlC+LuwMwxY2RYu34JwwQcOMPQUrT+qC7/xXCw1/LpXueN5qeMT
TAOnrVc62bpHLYR14+PAKOkGJNCsyY2CjdroPMCIjqa1MLzzt1wBGUNDiLkyVOVjtd8XtMHoszAA
zCBm1VXg6nb3vAYnP7/ybDYSJwzp+UeqjDFjL07UTVfzvpwMz8atgDVeKypjyflXg9dBt5C/k2nH
WL6dLAbZh1yu0uTO15AjnQXoIItOSDqRtnYLkM0/OYLqnMnA6Kr3WqNhB1DP+7prYb5ZGAD1BFSY
7WU+gJFecHWVKArDluWsnoopaQ70cnPvpAEE+MKiTMo/QBccK6yh+bj6UKnHjBiMyu7zeCPI5tLJ
kAaMknDaPNRvs9EMjHe4J5cs/jBjeaWfCClAO7p+1MfCnoNRLaqSBcfNMl9M77g0cZcCojUg7oxv
zofzbTzve7XLwgap81tyTNZtQx8bYVbwMaFwDu/4ZWZLglGFLe4tdjVWEsRclBkF4NX27BwFnrrg
YZj+zcdxiIWjrB/ZcHeI4FGj5biKIc6fv5ooQWsfT0F/OUKc6bewO9BcBzh7k/Y4qjKs7wswHpHW
Zgdezkxj8nLWobtIyKsJvFMeRCmEDvO0971oHLUZ44p2y9EipoAViggrjV+FPg4RSfh1kyAOBqCu
8hCl8pXCJuiVA8FInRuVJFvwXgAcWxfvvWmnfeirCFXrqkVnHKHn7VDJ1uhmzrCuBF34bikvzlrx
rzYjuMLBP4MR7HZNxe4DYPOeOK5/g7u2PLrTJ2jgSZqIq5n0J5MgTLtb6Js7d9JvIqhPfwzM5pSb
l4EB+LBjJV8jiDA0e/816rrlwQKIX7oosMr7NU2rahaf72dzvrGBiSzk6mKcQw4bN5EBzsroZdWX
rAo6i7ZxE9pszNJiHcb+AvuJMmHQBrkcFVbBMcB8pNCbGyxdxhf2q9kRbdE6Kw13z+48SthNpy/l
DNc0qeX0yLed2LoRsxacS6DgfKpF+n2nGop3K4j8/yP3E0JNhyE5nLeimcSwGKxFzbhgialPjqL1
UTLA0VKB4QeFN2O5Dwe/Op+QqtXVbSZ8Ks5BwaLFEJl60SSTQDAUctRZGt7QUBam1MEw4/brH5KK
wNu0BhkdeE4XZVA1iv7fzD6NqwzifuI+Zcmczc+bRsoFx7ze/M2RozcqUXjis3X5D3qrqGUkdsdF
cXQZWnSK5bklXPsev6EmOEZigmV8hhThbo7VIYMhyCuJK1n+4XVd9a+QVS8G47n+pv2fSTL/BmzD
41M437NAGgIOxUncKjQrN1AyBXO93DLK2ooW5gqc7zfhcslVHnOz4wfbB6SEeHEJP12WIK3hMQfm
UYheOWPIPzF8e19D/YwwcXikq+c1rFqPKWRpSVcDlKDwmfD7NW5pqeG9VJymQgo3SB4pqpogqbm2
z2ISloa2gUYdvMIjH7+Ik5Rc2PnxHdFDGD1g1lWLgm9gnEzoM7hMuk23EuOEROwb1zorrTHOJlLg
JCOB8eC8Fd2jR8sV1gB05s7KfnWV/yA/GXnHmVMnpwfIjPXFBQ+dnO1OFBcg/wAareoJvTbxQYKL
5bnnVvdD/m3hYxjLlI2JbeEkhRcaNMrLSoLL9KV8SmDbERp6BIWSt91J2129twNxFLiqniKf5yHM
ehotqK6Cj6Mr7g8emXnMu1TNFwK8dFyqmHsCT7ITSnfjjq3a+TFfRRBGSvX7Tmq4RFILPRE8I3JI
vFtchcBn/kTIjC9NFiTFXXKoNNvYyEk9nw1rsjLQ2OejJq4CAvcl5fIyjJr5Ft9RN3JMWaYVW5/B
61Y6UxQ51GWVJrcpM0mV6TROxKzI5RIvkKS/lPP/37mGImA/zIO8BVfcNr9CFfnUWU7vX4MXWaS+
NxCieWw9upc/pBvYLP922n0FDnPCwVfwycDGAcjYZeqt1NwUDzGRq+nuf4bnC6yGlf8Oy6YvHLbc
Fj9A8fAlk2yZzikgAuA4DPX6rAgs2ECYUWI8jz6qPS8ZX87HEQ6kTGxKurihUZGhOiHn1xoyJDhF
9vDYVT8Pjd0zCmot3rp6Avo8Gym38xN37d9WyKt7/4W7KcTARrjQze5iSLlnAosv41q0OFwqCB1o
W6QqxYBTstseeElvizJaEjrZ7Vq7W+7LsNqbyQRXySZgtqApz44PbIHZ3DkzvU+eJe3NcI+bqJzk
8C5KLXQtUaL00+S6kOg/j87MIaA0IogYwgX8Y9ww1IZUDZFMql43mklw3IsdgGxko+J8DwcBSA22
9exFCxXV0UCYuKHunWzOPUH2NzRfaEwCWiPl0Z8mmhsJovLjsCycOYi67BiYEvf+IjgGvN6xYlV5
YOGN2Pia5QjpxJjP/3QgUJ0n06MJ26BeBrXqYobZAf7c45glzy6g6ne+EhhCQKFR+buPMbZ9vh1V
weEPrC1MTE9Pm0MmZgqq09CFpy8ayoPUWPNU3X/dJ/bkTLh5fJbA05hX9HXZXD3iCiZwRctGnyCa
YpXqwVrbskFceg6s+aJKadek0nokLX7mHJhv90YMSH/Yv/25loEXp5tuLvzoV6rjGki0KGvBUXtN
1TqNWwaG17DnSnEGBXsa3G1qUip6VG8q1kyUyBzasS3DM9qkHQZRGGnDkar5zm4YzYC4xpHUdOuz
zLYwaZkWAjo2++BD+gKyKfePYMM/f08SdqLFNq/vnDotTprDycFpTZXiI2z4hri2BJJ18Q/IOgqh
etXA0r18C4tRsKP/MBiB/oqcjiss9dt0JgV5C5MexLm2VmgJ9mRedBoXMjv9FVTqFmZ64yOEnWpi
hpNw/dsOPv3U6up+6nh5PCsGLgGQQyrOLUyfISVtjAEzlfqgT9UAjpkuFfo8G6so1cMoW6S66Rfg
1hH2pGUPHyUIKdn8UfPDto0H4y2thK5tG+gE6X0PAuZu9DpUwEKFMAT1U7jz6pSKWnLyq5FCyg3k
bqsY1PK5bm2LfKwLFQCwH4GFG8RBH5ljR9YPZTRXOQ3b8tpqEn5g7pqQk3SDRGJIQ/5ZAn5543Sk
Sp3DH/WlgqZKEDw+2zJnz/9tbEn4e1vwieJvf3UeCjUcECYVpagm5HkdeZLXw1PHA0D6WyeRWQVM
WuS9s9PLVupTxOcWIE3xgQXatF0OdlC3hCsPuFgYJwD5qpzGP+2KAH1MSlTb0WdPpfvyZu6raqVA
a4LQG4WwbhSHgqHS0PSPJW+oVMErqj3/+f4V37VAFQW4RuRlfxiymSyt2GajdAxHf4d29HjqHA+f
qLDAd9o0N6prOved8s+wiWuSpmtf2/cLUZjLumwg8TMaGaq6bHXqYq+Z4R2UZtqtgVY+lyE9XKAj
5w+OdqnLlyCfnT93AE7FCdly4yK7/MwG2qR2P6eaWTDDG3P/k5yhyYEAXthqqHzv129Ex4HaZBV+
AfwQ4ffTlj4R0leXWNNf/Zkdo76kLCgxByIg5MuwlYU+5OmHUlqb6P9szuk8B5V/JfZtXzw4TkOK
pu+cwKYAOYHMI4lLjObqy34L5pO4dHnJ4KyubprNrnPNFmfmSNoyD8nmjDek28xqwW1n96zjpdw8
w6rGUj4NnuyS0zLevh1IUFZQZwCRJwTf18gTcHpLJH/xAl04KbxtNGhkaF7+HXp8MGxKwrkTRch5
Uo7SXdWqfjLN0n5jEODrCbxBWbS4ySj6QjKNs/goubET4fQR7XD0F+5UblZIb4Qdd2SYF0k3YizI
Q0m5YfZhP+ATeD6TZCLJFQRxL/H1rqKlcOJqBiKj9ovxOvt7+ywrEgZ5avSmVZGVjiYomAw76Yug
w9u1umJ13KLAiJFKc20GR0bCQMJaXKm2u5OmDfzEReNPXs3crEpcg832Wzk+TjSF9hi3vXmJJvfF
xAmxUeSHSsOE5WJp9XMSZtmvXxQTlnxovDyNWzowWmP2Gi72+4+KnTcDYcTa43Aae2KSjIxfRYOB
L9pxLx2GLXjm7lVA6aMJXFsdk9Cdpg883oOGtVUZDlWRQTXt0Q0INKoVfn5GX+k2SrHutszHJyY9
XLhXlTjpUthMdbzgKO7WKP7oPCcqYmMNMC/dcBHADS5KUldQd4lKw9D3YaK2JF8FuqxSaum7Jkur
XasZBVvlvRwzf79E1O4YYbxNuqXnUEOskLusZAJjPH40NuijP9hqQE2/DydOXopdDz+Wr306AtHc
zulflOkNbR/3o+ycHMF+lIKVmM3VHbrYGYMv0kpPAgEqrlnYNJ8UUAQVs8Psm//JLzwc1PGJhaXi
0+95Vf0V87ggHRN2Hk9hesAulDCrEKVMQQUabFhMzVmlRFRH2eSp+G21461zPSgiSqltpko3JG+v
mNd1O7Aet74QyuAgrrGXCLHvF6q/5Ms5TuV0d4hRHtqa/AzAt7MCDOsV4Q/QzJHmSe2VdsEt49Jm
vuJ0ELlpAMFtqoUO3buPB3nP11qSJ9ByGaKsIH39wEruIetbX+HbjjcNxk/YePE9nEFySWm7SkLd
08E7XhQGtSt2JY0IUZ1luYfIyqjslTj9m09xWwIPrKuO5tCi+y9GwKGP5/193TjwdBhpc9XrDjtK
qe6XmoLfWZMif8Hp2abVD2IFrAzZmAn4gO/wiOeol4u0VZFsmCLN1pe2VrhUSS9T3W4AcSM3nOZ3
d9LytH4Xvwub7hT3xVcKjgSUGajcvmRFL3iq2szGIrqakVbtvRIemvVDHumLe6z0j3bKpb8ML1fj
oYuia3pUCIxpDHlHkg0jFUceD7LO/gT7VW/ZljnnCOo2LeMlT9JR/eoC/cO91RcEhIxEHGZTPMqT
5+vD/kewC+tTno2fIaQgVDQZgPn6yFU0LKt32A4SmaFj0HBOzuPbSYIG5zdpz7oe3pYNjP9Ttjnr
yLWkjOa+iCkugic2txh9pK1VS8raHUYPUbORBacMzsk7d46qCbuhAOm13Rqs7t7lmkdCjVbNjUCp
jFY59EqTkaCGYkAZuKXMEUxVkbaP+gGR2H3G0CCdBbCdBnrBHls6vaCyqmycXK7VddQxC7S+392G
Ik86ScEaAUcDl0Y0coaslxvkefrXb5oGC8nGJK+MuLslybag7a6IiviCc0TLyRRlS1AjHdQ5P6mp
k7cq7IiXuckBfoQQjHVkid7aI4F9xAz+MeN+UH2U+Q7tKQxIgq5ZkzDBWr1H5Epqfo3ZaKnOz523
PsrFOC7jKsAoZNA5EKF1slEORa+P9BrKZ2v6V8dIeLvSEsXiUhlTU8uxz60rX0Cl/RyQobNr8rSe
g57mgatHMbMC/nI0yfA8yXOj/cZG0BD4FmqgsGnqT+j9E2RFBLTQuynpkmLYKi4yW1N8rWVSHsat
YyR0JHDdUcdSYAv7bqHVTOw/8Vj+2qupkqGIL6sR0yZC/JeNabDmcsPwDyS2wkh3mAAx+Nda0I4X
+PZWuuShRCpHpcI8Z2d83BlwxjUGxADNl4pDPEKw/EonvD/6gtisDF7a3To8ZbVQmO310MQyL7sZ
p9itU/nT6Y+ggZ0yInUD3hVqsmOXiGwv6F+kcvd1mWE9uL0z2FJNX51RnplxVKdUBnSelxeCO8VB
XWmAkg+ZwuSyliOgOTd4y25fOezfXLGi5UdfNFhH3ie26Y3xWAMIEwlLvz9crc1P6JKAZKhsw4Ay
9tptZtsw7zYYmGDPLsW0IVO1nCV27IeMHkWqzUbljt9L63Z+8WVHhBQVOyqpNRZiLQ8qsv08zgtT
OVuD9VYQ8r0WjORrX3gkRHskFZzK2a/DmZFOwU7lN0EtA34k8w4UQVccgEVgjntHTS/gJ0JSKrPf
Ua1Du9AUCka+InMUZCaSGj3rYN0nnr1TIcMGfZu8CVQ29iZ6OBZKtIRTf05d2mfhVq06FvdS5/aO
EvEGejET+XvmcG7bJwLlBg38CpurHSosUyjanDFEs32LD0WrfltJvnm3KTeCXQ2CN8w/678VSqPJ
gKq+glBrSWkfyLhjVCbj/7OAGyHSU29IvHfd3UCRIpDyg3VYwNnkmJqSStLpvsybEw4Rl9eb1RGP
6UIk+r/Gxl1rayXKQThK9Z6Mk34mYn51AxoOH19kA5UOB9Q0wTElULJ71lRenihFEw4PuoTkFvoU
r2HqcddjzMzsU/41t8kxoFDAPsRhYuK7AMEbXhwoJsMox/D3Vu5eXjqgqrK0oY8iBhl5bZWNxfsb
Xt+uza9mqRxhYm/SquGGn3t2Bi/IuC1XyYHxNW8q7jQvQIsy6k18jnjgpJpwjiIbWb/oTr+kWhKK
lYozSy9CsZymkZ00Qj4lkpHuwBToDEvZoQ68H4ekfyW+2YwsFQlNCWT1hYIgwpNVouiDSABP+cCg
5VYRt/5zISQjwNRZRqg4Jtsc9+54o3jZUpBEwfS+NmLlEUV50yIz9NM3z/ZqjzzREGl0QzJd5OOb
QsMXY0CwYNk0hjZyFfjIu1sZtRnfwbq1gPEPVeKBeRTnNIZTuKec51kuq6i+cEZIeOznzXOxHKgf
7Rdqk+i/eq821IQ8o5aNoxYfk5g8vIbWlbt/V/gOlDCmz0byrlE8ywzUwRzhVxv/S6WFIpiVdq5n
zRcXhyXp+wS3QzQt9lF0U2+B9b9wv9K72yoYKOIUcaRh9woELP2QEFIRq+j8wZ1q/XOVkwuCsDma
B0uE3hBD10WUcubMgt9ySNTR7jx0dx7H9wsWjOFp7IPuSqx8vGNXQWUwWNW72N8vJWMMggRXsPt9
ralX8wtteEyRwpt32bKUa7i2bvt8Dg+GFo0KU4M/nO/e1dTG9a0z9tlsqNwZnjMQyntlWoVDuQhT
FQlMMW+/i/Qtyn0z/gRDtIQzSGPGd5K7v4mE1fr0XGWaKvfHqWJWweXwXppF79CK2Zm+91JgGij5
bu2THPH1c4fRwtXo4Kcg7TkfvpNxa8EhXoS12XkDDGH45NpyuaMzMclJ2a/dW2asKU8LBL5Vlyen
pVa5NCJ60rAssQfxvvn8IL0R2doqDACwhr1zeRQhKzdNzopPiL1LL60j26Y7DaDgyC/pftomG75w
PWTSmX7VE4SJT324eXyfXLNndX/mpZQNd/FzjWIg9NPP9OqID4fKdrZGv695VwXF/S8Sxo9NoHS6
SuwNgb1ELgjZtatYxMkGOSCLFC1/WxGuDKnTd+pmseAn1zn6wJ9YenhNCWuxh3vI4enD5aGs07qa
ZMRrOSYvtKonkPM5hK7EX/gHzs33LDJeaQQSSIJE3hthKGbKxuKuayieJi8npFH05HGipb55Ws2k
AKID9qH7bKxemyduyoWumQTl5XU9sXIHypGndXUSflEOi0XIb7uXfIFjYoNAWBVNGNO1sdG1kz9m
ptvZklBRqiKNw7bW6V6JI6g7oC2CFdLsmhO12Wvnk27myrRYxl9Gx2rieIecH94tG1OKD81a/pC1
jAtW/hEs8Cm8yS0hTI2RfQEYg2Z5X7Yn1BeO+zAuBu1Wmhx0+euIziKFYDm09lbPrPC6TMZiQyPs
GDaPe+jS/Ye7FCN3Ee40u9BwWVdqy5kME0fiaMpgJ39bhP9ueThCQCXMczDg9hdPDROPJxxUjne7
FN6lCfQzxsmXK1GUy2/dIbVKsB8YQaOWmlgAcqDdg3dVOBKhjt3mT6DpY5+Q0//J8SNA2Ly+3Cqc
qz8Mik6qlTiPAblAwd7TQKwVQlc1Br/LcDfFsCdRjZ+YUev6vh/qnb7Eqc+X5ekcaZ51TWDwyyXm
OQHw7O02wHkh0+39meCWlGAYl7EvwHO9oW0xLf1a2XRRJQt0STLFrBBscDr6edfyD4tzgzwx6h6e
NpqF7UyNaAek+pdSjWXjHIYOJTmzRHSo7ZXcUe0/2VQHUvzR4PaYdN/5T0fMkA8IDzQXZGfQXBAE
/jkwBHt3WCyEqILefq724w7LivuFRrlpgbzYv/7xeMoU9jh5d+7fzYWkLRzu6+nBsVP+ugvSe+bQ
ylIYvqC+ee5f2mFRl7RsXULjZm5pPnuOnSJitxloDNGko3c/sOHTMCy+MxEv3xqPexdEYFRroZvE
fIUCS2eC8a6L2ALjficMDFk4Qf4Hytr2ZI0ClHRKXh0X23fbent3CsjV5vWQ2odZmRk+o/TZ9sH0
kDIaJ7I1/+7DCLGu3H0bLe1cQtDd8IG19kqML+MN8vY8E4nlnSYzGzuvrSc0ve9bEnmH1LyZDkZm
mml26WSNrzg0zqMK3GLZuYNsPShLc1GJ+AifrOt4SNm+KwQURx4kRh/1z/34i0oWP2eQZ80+UU2B
5NdERA19csRhZLNOziUd0rS0mtF6Fu1loxGZTc9rAZ4gEtkjVMVoAgqonFdNmAqK8YCtQAaD+1hr
58jtaRZ50e4a5XECeVV35CaReeEaYhO0fIS1Od34OjQjQhva70kqA0nnt3UNGRvmLI17ww2fPIQV
AJMUIZOApU2GL6ENaNGkmwMuF6E4alu7SxbMb0O90tNYVkCyLiruYo/D19oyZ0feJ5iqZRpmGNAq
AUBcYUMiAg57Nre65M1mkKm3BZPGSqIMHhkcrq0AZGB/mc+d1SoIM0f0VrjGEDX+axXkIFUBYgkq
gdpYqTUyb2fmrkab2Mq+SzUL1HAcEke5eIaDcUJUSc09BcvGO1v6A4/PXuVfcN2msohIR6g8FZzx
Heti3airAWASpGd5hfuedsFi+vsXpd1czCMg0+G8Xu7OmEK9jNzTtUUIl1BqM6Udt8u6FLkaHyed
nxVO77pMxeH3HhGI8L0tlFXQgklHBYv+mnZtjsdEQkOqxefeht6s/pT4YKHUguNkBicEUSE9Ghh/
Qdallzff5Okf5ABXJP/Q5knBdXi8fdmoKBULkJE0c/0SJ5ZvfwvjEcNH9ZGKs+reDeGCFs/yZqiM
+pwL5PqXIt/VXPFoj+JqsyUg0clg/bBT5gpUQ7h6bsHI/5K244goMJLz1/jsIDpqScu4z2erdWui
r5KhfTizVxOQp45w2X2QoTn3kE06ufZ++mMejkLyhknKsdNTk9fje1O27BCZAT+2eBgIeY2f9/cb
EsJlRjMGAxOChSAUMJhC4ilnWSthfkgsBW9dCOMZo1E+cENlYq/6o3MoXgG/azjovpCC/FPoBHhi
ObkQnhjmT/K2taHauxxYmGt6rAPf3l8HCSlWKsJOdKhTcIY+ScyhY2yue5JgRklTnRfW0AJo5zRp
ro4eU2oeZsznsGxLtWX7lykKPGfbPop8IVHhsxtKXtLAFHj8sBnJioaarJsbpJqe0dPmHsMRdQa8
JOLNTQlG8tTAQPsivpoDw1Ug+5+vX9TeV9oLx5dOp/SgdQ34zTLzU7SRhkQc5zQc0UXH82F7/CGE
rOeiaFKM8c0T1hH3Ao4MLMviObvWrNTzD85wKCIH8mAWmHPHIdTj6DR/F132cp+Vqg0zGombKRkR
xblbDMCaNK88bJ1Bsc/vceXLaFHek2V9q7I2ry6OmTnVoIRftgu5yKIiNzAbGj3+LKVBaSUZGgWM
neOFCddvwURUQsgJxvSxcbkeOgVnnLt6ltI+jmngySllO96RD+0oKhM4ch93uoTkAwv2jIzjZ7s0
7jZqJfJMz4agUM2wdBTgXIZpZDszZKBTKNXfoJmTxG3S+NExyVSoxU95JzGGlYGN3qDDA784C38I
26wPOPRzunIqnrbF/usde2N+03DrGHjE7MzYD+khk/FoQzSofHwmC2Lna8kNZpAaWgAM4H/3sV98
UdeQv0eUpYhYoKttxRb5kjSsvfhNSiIaBInMB2GEW1sGqQJpjZG8mjPsEdQhl/sGdOmBPkPSht44
d/Lq3FBQqBerH7Pd+mOCdE0ntXt040vWXqkMjnRCSuTsc4PTErQ6oX9E8gQ/Fdcknqt9RHH1ZsqG
lx+0YiNXjEYlpSOtp//m5P4VHAnFz7+qegUt3K3myg2hNykQqWNABC01K6KE/tKerFQHEI5h5gEF
q/6zecyeC5qg7DaF9tOIJ6Pp8ZFS16cSZURaP02AQR80ggTeoXPb0Rr5j5vOxepOTRwJvb9i1qhT
eBH8Q2G8Vig5O//NYiD/Wd6XkrBAJkjiERJ2qf22ie5uHxN/ds54GXB40uysYCS+iAWk3h9W9ZsB
tX69zpRXm434CNHi3jNwrgCuToi5ObUnQ6ffVb6gBYXOfL+PzGUctviNP2+2p9A012L0J7gnw1WA
1niAcq5gekm5SVixHgoE4HbsaUcbGqFxneS11OnCNMkJrQQq+bLAUor0OD7Goml65Tpk6yRkPp81
RJTWztCSjdJeHIcd1su7C937lEs7rLkRLxVuHN40YO4oooqnmzTByOxsnM17MHrbaUfJKzRPo/jg
3+Mn8Ck3UmAyXpnaQwjhhbpH16TlcWSmuMaU4NE+gKVRqbOHiVVxbjB32/BInl8ntn2ziH8FciiK
s7cUuPWAiEFWXhPgwW8ASChy0mJVM3oY2EKbu83Z27dfJ3ujIpQqMuTnmgwsocW9ssFme22Itcuu
UfI6jr+MJ1w7uQgxxJiNszqQ/vp/jgYOZkxyLBMkia2frW8Xf+20kxEm0VgdCrLCvguCdHIRFTM1
FWlOi6s8wKAnvotUMz9VCKlUwScxRZN7ud3QT9yL/ITU5JzP7sX3n+KtBwbXu/RrT831fapVa5iP
HTW9iGkFHykUfIb8aPx8adTZI9kZPA4WMXjPqkSNVc1EZ7XR6BhVWcvP7NK97RtW821QkGTQa1OA
taG4ZnI7Sn2PG4oyMQhL+nAOJA10+qU9z0nixtfHAHGbEzUvo5dFio6ikycsh6geHbamQKyL6vzM
nsazGEkffPaGPhZh2kU82pJzUoADk9bYGxUTrSEwYPx8Nv3NN0slEsc1/e2/nY4SKCembLje2RNx
MV8eID2n4zzrrTHtmBWrLTto8+NkfGzTsgp0vUDHg8AAdJDFQ4LKl70mcxF1hz6QSJWLSpHTghF5
kcZEC90dKui3oW8tOkBUGf767Cz4QD6ufAHbcTt1SDF+yW6tDghjBaTGfj3sSWqu6Al5lCKzyze7
+kISIA06IpCRTtAP8RswrLOnOlRCscp3ioKZ9hqNNcu7cECP9FRMcW9jSWIwsAPOwFUeORZEY8vu
2V3PVjCcBncP9nnfn3WFFe9kx8L6aLj92nn0ZyfX2MrNyBLVQGP5VcMnIJZm63j8pSi8uDqUQ1EZ
DbZEWf5VpRfY3mjXRG/Onn/DLG+0xDfS0ravADJcuXcUhb0iBFpQixs7BDL4WFX6Xqi8dLn1nMbo
oqcwPN1sJh4G2kKL3QP16cRJflHLxhswW6P1VNv45nGdPLPOvgdOm9D9RNT30a6XmbynD+axk53w
/H+ePboKFafiAjZunMKxqT/r6bqrCN+tu9/Sr19Sj2zKw6UNrVgmsR22AlzBkPZ7YdzS9CyURTN+
YN3AtyPQ3z+8jnyXK8ht/6CgQ5md3XkZGq0TbLyS/gDeC++N5xLz2ZQL7ziEkHyM6HWjB/FRGz0k
nvHo7LwUO7+MBnqpvwEyObE8ZLCs/IcSV1FwnmsgqoboV9O+/QABLs19scPOWUnP7E9EjdUJSyUi
lO+6NC2trHSW/FO4llISmKLhPO1eeNkO4kCyJPBt1FPOS1Q2brPkXgfSxLclQeh67SMOhU0jdH8m
it4caWgJtp7s9oB81xHhAiGZv9syYYDEtNghAbfMXtHJ0IHNn7ZLb5QaZkIE5iPyIFljJQFUbXHf
jR4V7wrxHeHr/cwHGf6hXxJhDxrAoylyXd4SH+4vX+kzVEEhgo6WG8+9WJBT1nfuXW4Fbf1JsXoq
vKitIgCvUOAfj+X6zlOo5gdppXgjNGkugVyhOvS8DiW3oI4HJRKzxc61OfNYTfRDkAo6/7KddNsD
9czo3UGafntYDT2GBmXq/OEG30BaJiq/FbdnirFU5YTjmxP/eMQwxGoJxH0mEBip5UfS+5GC8Ojy
VO5OELncEiHJF015K8j7yJA4cYnBTcLWn9Tl2W8Z3jMzHa56vSwb8b6+DCzk0POr1XtJ5pQ11+Du
9DLia0Ve0im6qscNXRmVZRIutcw7GPdRCpDi1mIFKylC/zRaMOHqWdU3NXgQQSTGdKuDzV24BMGw
5+Y8/QCNiRvC8ooMYaC45kKC1fTEGMsXj27j2zaK5VgXsDnJTZMcvRZcnbVPbHM4ad0v+t8df510
hXYr686txx2gn1vRs3/l+P0Sosd8R3XjwkXAKBBgyT1KtQW8Y9nqg32jQp7WEyz178KTGLMK3Y7y
Anquq/7TtsJQZg7HnXO/0prVMpk8ycsygbOvg0+2geIaz4/xflOMYUf9N4IYGyFK1JUAnf1v8rnx
TPbpo44aiCTzQl+hfZkUA1B2LBc1QvYE3y7qLK7D7R/uAcS/rO+pTn9LrJcT/+0PzkSsWUeotZwH
vYLUiRlThEKFZgg5uWrwWXZjkJgRH2VXURJwcFopWUV4mddVCtw6Dp9aExXBzaZ4SkBE0othQh81
O3T5JZGfMCPwr5382+kgl/MpsL+IFQRRsANQJ7wDJ99p7E5NT1F30U9G2iMC6VFheOASU27E3b49
131E+0THIkC10qD1gxB3u4bw4mQcuJyrBqmSoN9aSgqSXnqx3XVq4qHIKmhh8rSfliWJx2UVg/HH
yjmnB/DQop6uPYtFC/U7ZWLZFYLm4H56pGgM2yhLkbEKxY2g3AKJrOrOESlc1EOwsps1Ir9h96Rq
fQthnUo9KhkhHoX+/HGMrsAinVK93nm99cvuMmkN9EA3v/CLA+JX8SjFnGfp7OtypeAN9HOuJo5R
htJEjdc0ua2PzyiBDzpl7flN4IdqadCNNEhpE2FbRqg1SPxzDKuOUgdJbcZG/5IJfc1Qq6NvGE0r
e9NTwIZF+LQhsqGcU7uRXqt57UUGid5lyMnw72B7LDBR+RaXAvU60AQhBjI/4BEQxtxnKQsbH2OQ
LnJZi2P7GuAolBQ6rNnLpwDYJOXquEV0fatsi/KEAIzn53XYwGWcaoFpPCPx+BIXXkcoqJnqlW1Z
DyhYFedRHJbvUm/4MrQwzSgcPg8RTrhg1pw/g7HSOMj4I+RvAkU8lzQqKE60I4hQOzKfvfWc6pcr
3/fHCJqSLuMbVS+CLpUyF5HsF8Hra2TPiN0dIembNy8SJ1+WqpzB+1WvL+udw/kQAg9jjdPtWvkJ
v7d1aaqkJ+hdR3kDTo+cna49fxwSt8CHKXBFzVe97UQ+jN2hmwsVf+PWwBfJ9DR1EorrTMAGutZw
yTOoPNADnFfvCdNWtO4RbI+NythZVQEKz+cO46z87xDRiHgvnZqZLJlxVXoVfrq/MoQOSeanwEFE
4yjs5u/4HDd7gYYSkeqiYcnLWEToOrRhLY+0pPRl0WaLL+VllQPnzZcUCiE2WPizpOO71MVQ6gc7
jEdDMUtUhEos7PArwpOfsA9gDID2lDLiE3/on2Gdjm0m1iHd+CsMzu50FM1OvtcW+0+JxxNmkMUX
GFjKppx5qpDr/1vGobVkmRPKLY2R6RliKfN3U/dxqRTdsTa3ezknVnY5KW7AujGbG3atF9CstjlY
tUz3tb8qNr37dZezHu8Z5LU4nwhWwzZ6OrXCzR05PT/8739aSj1++Yv4qLM2PlW69RXx5RgOTdpl
g7vfg5fm+3CpnXYPaWrXmZCi+8bViMl6Ce5BGsVqQghfD7owjcF9WMp8Ig1jZeTzaRQtweL9lnHz
AEtAV001cSLsKIb8Y1HLYYVQC8Fatl68PVK+6S+/wi2k3KkIZu8cr1p0P9pWms46chb/wbNKUQP0
UJ2JMmkUcQpSUMZ9KziE75xxDnQ/laBewM/vHLBBnOygP1B5+WENY8wYnt1krIe9lUkZUha6Qu+W
WkLJhNnm4+XaG67J4iUgpab5SYzq2rkB8quaDkF7WIFOLXxbIuwfy00eQ83qpaTF8XCvDNc1W1vT
Jn0/h0FvT6T5JQw568rQZAIfbJ1QHi2tEpt5BMtxkkB9HPh5DlRCKSPXBkQPpazPmZtqz92wtD33
E/FHsAbSVW5DjbRF0liTJ451BSbJbs50ho3sU1H8G2d2tiDivTwwnQhick7t/asSXZDhPcegmRXB
qmeQ2FmoxjC8DT3mE5ZdjWAIjFxNq8Z+WDACYbbsRwV8bCEkQvLuuiMSpJX5PLeZ1CrkN8eJLarb
PX6FOeNQuhIK6uhqJMIALEIUiMCX6qG2a2fCIMzR4v+GuIe5UXOZpRVYMHaeqK+UkhxeKruVYmGQ
qGdXWlYOTQTxvB9buR65tx8nI/7Pacq3EXNRUX7tFdGQJemBspRJqiUlFqjopkpXWhaPMpu6dxUj
u2wl9ZZPECjRAu2J9Yhds7ufRywCJGJbkrHe2BKhMFI/H/Zwit4QZr9J5SRuRrLNs3CiiwpRfC61
yB1SZcdzsLpWnXlWIDuoDhRQw8thrt4RtUR/LoFbfrN9ctVB1CQ6AUGrIORIbNlnFqX58k3aFI3N
G+BECM0gG4Xl2JdLNHMmxXwgTliopdfB1EiQ04d1TY1zhaSnXMrFxLFTxEGY3NeQnzE1Mgxk4co9
7GTTKxmlnPGxWwdgZhDXgSKu7TciKPx/WAYMMXq9NnEiz6wIvYwnk20Zr81MYgSJuifTDQ3PTDfi
jkn3IR30dpHl21Wni/8SgKSdr/+LFqu6dMyR4XP5O9Zh54FdVCFUGbVZ0wgCYVnw+KvccMAbG1z3
fhJSbqvNpU2+Q/eFGH15lY/3dzyvfJySlCl6DNfZWhwyyoUeUIWdWzfMUEY+j9iL7TIFT0V/jDcN
I7gOIrIM0iMTa1ud91TkHdhvEI1f59PC2yBZsRJQxKO++Ow2y9GzhAkPIEo+yWlyg6BUALFbaYrF
sutFTTxg+B9qxXYkn1vFHHXsz7kV7vlTPpkK5kxNB3QQ7KQX4Qv8Zb0zHI1uopQin8hR3GGk1VpY
JSCAneSuAY/zyj5ljaxLkv6afU46adEhCImTI1ZZ38lO+lxCh38+j0YSeggNdJISAP8dw7Vwfu8W
6kz/BCybRTX+WHIzbN2Kv12Hn6S7FLIQ/SlBlGBMSJcuPvJM/pncQOgxEni/kFk61fAjpNSrAGfd
wHP6GaNhkPGrvKg9ihAY2NN99OF2iyC+DBjrZ4w/P+aYxrx0ZhvrviXVmrUmfnTjIyROviQPDp6V
RQsS2jFyuS+jvIXXTOFCvabsYYdMOjfg1vmq/zAWqDHitXm1Tqu7HdmD2gj5FoyRgq/bXidNPdiv
yb2qmnp6c+kyCON8djkI6T9UJIPu7gtr1YOhdrzduVVj2/H0nn5uAiRJARLM/QlyMoyQL+ix2z2P
t7wsVYSjKpyHUcJdc6CiEQ58ia+zaAXQB0Hw7OJJd8vOm/YYQa3izXjmgmn8way3glVV1MnVrar1
lu9xpjyRjFIqTr2d8+Tn2YzQ8adCjSnB0Dyb9v8lKUlmETGupbzP9H8Jkoun+ZmMF17FGqp8lW3S
mbcsnFQfbriqQnFnLxrZGVZaBAaO2J45grDUh3evgYWqp5Oc3kAQnwA9Czhkw77Lj3mjtpiKl4Mn
XW4IvogFI7VmZVo/qgMkpGQFowYv1CbxWhpZzCCqaLtrqMlHUPnenTloAzWCRSG5wF6Xwthhi3Jj
6zwG3WBOdq6iGsx6S4Ggo5n9HAcpexjcMRyoXyDRoW1gqXuDVTbVMm3c7c51bza8KeORoj/HkFg3
a9W8sWsmVTICpIpzCagM1kefX/J7FQRyxJ0sv2gWChh42UixyWov5fCC87gebSkZtaAI6ZkU8kJ1
zbrjFO8ebf8LoEbklhdyqyoedODv6lQFMt2AAnTvZcLnqx+WPQQuoag2jfHL6wmXx6os7GXrqdED
rXBKF9EqQKfjSnyJ9YFm5mNSjBgVsJ1OmUss0HErqWcUQXMxiGfSYdIPJMC6ZNoCBgjsPcBJiZm9
KxkQ0nNuTKg2iIKOtJaBVQQQjvNjf5/JiitiM45JCdx/W/8lTffp5+B9glF6gcaIn4nXwoiJLNtX
Vn0xMjurkd73A6h64t5hZ7uR7Ty+2XinN2V8JK65s9fDWXg1pJQpqxF4K3Ki5eCVtcWrvNr2NltE
MyB5S41lz+Ik34bYteXy66EkRK7ba9T+WB6oT7IKmn9N2Fhals+7Z934N8k1XUV0fZVQLiUMLYV3
9fvc5wm2N2yQURPMNLGIF2FdlzwurifS5mBNiUv55nEnmayDvjIFLdd4NqeExgBfx3+mSXXHk/SJ
6wx8Qi+EZ/xY+EREahr4MkMI85Ugxb1f1x+Q62/yzNI/qbsxSqHBPO4OyI5q6AUBiSDz5jpCDp7W
rxRwG9pPsWEebimqVKPdRxObFFqnFk8fIPR1/F08dKg4j+1Gxkd0mnVfg2AYJ8Wl9EnE8tC0oRgS
/1NwZgIJWINyU3pg3Ge0dzHzalHB5Izm+DDh7dHIPAWjjp0nejOCb3x1l+XPx3MM3AgikxWlm5s6
CJu8zLBEVpiqrQ1X7ekyhMlPHiP+MviBqBGMJmEfmin4g9XfSM96WaescN0Muw07B4mYiEf/qFlK
aP1MJ5GWTlDmvn0EFqbqXstkA/vkXSh51xbCmfPhK6fWlyfNwLGocPVljWiGmNjiVbIiZPdVF/IH
8vkalDv0yeXmI6Iolu0Wdm40hB8Ej0IY6riHgA3rAVqIeG3alkIevO0c4n3p6aaBAdPnX+K8xERP
1qKEzGp0RWym4D64MBdHj6i3uDSU9Ccgs1s9VFjqHaaG8/DwP/m7Z/eQDuqxLiJqkgQvn6rgI3sX
7e4SLqXb5R1o5ycx74eBWdi0SBphWwcrIbSqzIr1bIj8eBZ512O8IR96krCIE0cb58ptejMvxP9O
pJ8hiQG2m0RZ++EXTgB1cJQRq9G/lQrfWOVJJcuZA+wjrYKGo9tsAeKWQlh88yTfJ8NzKkKbL2ds
3KXCm4w9kYPFQ62zYoWtbZdRV/50C6FmIChg8NAz6MEbI78QyklCUuFcgrFFa3clN3h6k1QW3mN/
hBZTc5r23SaniKvngsyff+zqXhA9jqiYK0BbK2DcWUC7UKyIMVrLLCDRuYGDFNkkn+b9Nc7HUiuo
AgCPci9F1NPiH5n0PBafLBtQmQuh3sP8MRMNB2LGmZ7CIE7Zf7VVsdyL2fvVOWeHXt+KLfyIJjb0
hS3N88Q9eMIQKMALUz0yCA+8tQ1E5iA+OCTb5/ypKkqLoudk901vcvx6j4ao63W3pltp1BwQnpXf
OBAzwtaECFFJB3KxOdHiswIWFoia1UlvTvH+k2zG00gLAmME81X6Dhw09V4e8upBRRDdYXW9J9Z5
9HbzU/wPVjNnBx8oygmWgobTbdaaEY9PggTkUlBBeXbb65zuj0m5bcvmSGC/XyiLDB01gpwle3Pg
LexGW3jvSk+SBinpOb/KPr+NhN1AsdcF9cFCK075Tmr6GNsCEi1aGmthoeP71zgZ4fkfWFEcBn/R
7l1joWTm1MbCQ4PXi8+KEqvgPpH4J4WlvLJVKcBv9IQWit3TTbPMrlu6F6pt3yaA6fo5N0n0LZ8u
/XXVyz4NCZwWdHXv80+XyX56xHEX+AwrkkVXpcbv5FmQfySGDUTdOYrIwnce6o8Gp45/Oqo50ytJ
KFImmSvdfwjZpC1icN/UZ9MVC/7OKndZT5fiXsk++t5GOzod/2B0en/1icxrzXPbCQCVEwrrzBbs
b24cTJ2l88G0CncBKn89gYEq3g/T1MQWCkfRIAbRSDFsDjd6OIybFYvHxSN7ud9wpPgylgrUE089
31X8zGo+vOYB0hQ1yfLD1OcCpcB3fn5PPHGc9r/fpWKd2hrYiE97ZkVOadXe0wKjf+xrrY4eigtW
4apTks4GErWMfW6VTWqYnuaYIvN17xyZgD8dpEsyick6soh7QIE3V5fkMuC6mPi+zv4CSkiDhS3R
kOkDF85CLY5wy7bZOiQRSkzHS9ae/CkLO7Y6i3yOUOS83Yh2Tc/8dACs/iBTwwd1zXvIXDMUNvfC
KCPINuVXo9TkcMIaErgu9nQyhA79TyUExQnJswQ9gk9dmN/hUqv6F/xCHC1VL3Esb/0xwsUzTWTa
a9s10z6AcvoLAP5oR/qFKo81P4sy7mmN+m4ibpXLkodKpGqSo1g8/lE7rwdXkNi4pftCYG2zxvwB
K0RMNpKkDkGdbvcbIutlpdg5GbPBB98AIhfuIUMkIHSwk4wcjZjkE516WqYM3MxT4RQamY2TasTr
jL32uSuWtlrQNsjVW9uhN6gjyS20vVefu+et7G5EaWU6XZ66ChBr6rEBTCFGRqGp7oLedKtArFFQ
HOIvgACiMjSd4IlpCc8Fiml+/JCThZF01SB98aLA3v6UjXjDmG5MFyh3RtBra7OreCjxOhHaIgXf
7Sxma0nrbdJpYSfnmgajUY/BjqoBt0RHLuasSXp1wFGh3SN4snO/TGyzmgK8ZfFvwcCzh5D0vfSS
o664g5Jy9zUckTMSdEMNKngDi79h/Nol8zJZssU1qdApPCt9K2syTBZU3ce8/RhjF9eeTWPq5C5b
ef+YYWS5bskxWkkYNgX9O6PdmprexCDL0mrQbVwegd+pECEs0b0EynI8iz5idbzC7nSIFQiPFLwC
rHgoAtWLEKIxhbhkmmhnUs8DXOmQtv/AazCqfLAYCjbYQ9HAHPHH943Svr6y1yp+6XROlPsPZB0y
/oPLcW2uLFoKLUsyMizI5V7Vz16wxRhHp5KstB59V34+yGMDqGxUI3MxQw43DP6Utr7WwSLoUjUp
WLCGlG/XxaM3BYdWKx34EjfrA5qSUrsSYCZwZMiYfHebyuxHtPD2aTLCbZbWGzzvMnnmXymAakvY
MGXqI+XNqWo/DHqqZ0PC3IPhB8X9opsO3Qm/i3ZvDbQ69/tqG7RLGX+P8q0ErhRjdich2y8NE8+T
R5BSe74po1rNpofJ/mOvRY3BlOn7rcDB4IrpSMT3aP+lyRwbaotRo2nqyfgjHkBiymmByXXYuGeK
i5UoUoPUP7eqMJu8k5CaQFb7Z7IMgokjZEKOYJ44iXCu8+AyMdapGYNNEykvcS5VyYcZS64/YAS9
GFSsnrFcSBVQGvIUEeCCspbYqBIjugXwRD9JPGFuKqRJTAdgevw+opSXf/q31hP+d84ugC3eF4kn
8kfp4tBicSeThew4XmPJVeGDOdytQ5oxp+mRRLQnpzZbCyqgwtggGLwYAWRvMf9vgPo0q1LMdfkc
proHoRpu8cIBGFaa0i+zdcIkT9S0pQG+zeyzOMmqndxloIhmjYMe8MHoVb7hdif8i3C3VwNSwLuW
pUGDXf6y2xrhzIhtmLImxITv11PQ4CMqCPv648ed6jrgowtU5dpI72vuo6n/EKiwPpCeWXx5jbbd
Ku1g38H5tpgVO7TAnTIcdSERwRGfnwpGTcBIVMLyV+1Mwni+TnXaMSXDUh4RCy1mPLYmaDlKfvjt
gBAqmfQliHUnqeBrP0PuuNt7VHH/GLP/LhG7KuAATU/I/tQURLowPcAgCrjBpG75bQOEloA+FxBm
pNr2wVhZss/osgXP00OIEPQmtd4sfxB0mPYmMRXN8qKCD7mNj59Npt/M4jcg3q5FNAz/E1o7d03r
KjIS3d+o1Z7RcYJ90wtorjmkneDl1LCli0v/uQ3smYxfQrizwQVTQ12wQWLWHLzrf2HUoN6swhmV
bqBqj5vb9rVUx3/UYjy3IT1NySe2w4UrrTrGyYUOQubfIb6ETJCx4u6cBKKuMavsVk1gMEqj/F2h
wx+DHCZiRm3RPh8Nz1JxyKSY23A5V1zvw5lD84rILlP+181hgJTs98ldsgymK0SgL9ypb+p4gh92
gQ82udS6Jbid9uu8+PXfu/0/ufPaElyO/N1P0lueuj07D161nY+GlGUr7vWSBhqaK5+ep1CU+yJT
agHunql+CeADKoFVeiDXh7H9c6uRQfFYnqK44mUFMR8yU2hlmUwraa2RbMJBteerc/0a/PjCPLRw
LbNFxsBtS7XQciUr0n+QQZd1mhXoQQXPKj2PgCSqCozDqTuWne3gXFWxtLiwdk8OB3dLh0ZCHK4J
TQivL15KaYXZpyEgJLaO+DzNJrL/1ggXGy4tBR8HvTqw5zTp0X3u+vPqmGVco+hKbLc5okpR2QzO
9NUkd+CB/eXm8YBAJdPBwOzOxrlfbZN4CGLbU54JxNcGRfRscOIYhO0e2dcn8H2G0cPhdfKxkHIp
S2bxbHtWIQQobzG7AfJZ3+sizZRvM4y6MeUSOrhwzqpdymZx59vC6E+fC2W/R4v/XcJVT+Cd7kFu
DDnVJgoCnxT/fbKYVYdV9NlVb21e3tVssK8LEj67vyO6CJ0F0YLPgGa+B2OiPhtXTU/bv6FV+AA9
h4OF1cLe0b8cZ0st1kkOL3+hDmcaLvAefnR1eym/ybsGzSvR5We+I090pq+JIwlaRBQoNv76ijXb
3ySUh21WQu6IjkILyU39Ts92B+1bDwNRFvP+kYNnWS110FGe7KG+9DTips2YdFPjbOoRTeMMo2n8
cqOAcfmqZJ8ewwuyqjnlYhJ6HmjOMSfDpqIlRk/ISpXMRx1w5EZLfIRNyaTZ+OsNLAFSqHqmcG4L
OP2i75T7Fpk6TMBi8zHK5Cc0O/c3yEyYus70jY2ipUFbK/Ug50Uq6eBMDPFFH4IjupX5yfJ9/vgE
OifSz47tvdvO4W7BNYCKKP/k7xuWTCwtwbB1nlONAS/twd6saD5evu7uGL/ogyp8mXHUc64MZdM3
GQgZy1mluhPAOpS2z6CsOyzNxKiAnh3hnJAG5o2FxYq7r/vTXm2aZKxzp4XWU+qoSA50+DfeU2r4
AiMnhBTiqdH0GSkICVutBKaBBF5dE50mw4HAdjylu8qOou80Ha4JZFOOs5LpFxw2HHdLKqiGagfe
+ZyClTz01lUChVkwaWITMQOh4zEmVm2iDuSw245/ANhmCwjda99A8W3dXTPaXfm75yLDn7FSGY0T
LIMsx+WjZ7Igd7HJ3+RNvmO+pRvYj0oG0+jhU98N1JapuJZ38C0X0Y6D4pqif9h/9Z7jWFFn9t3i
3pevUFVXGVvSPcwOzt5Ppio7eDdIkFZd8Wm4QcaFgkeGGCBW0OlIS4Z8+Hb59L73w9TfGcQZ+9N9
klJPcCBbQvOhcz3HRh03YqJ7m39l2XEc0ibKGwYWxEj/pJ80VpkF48/3o4XQWoITDYs+/I2YamRg
gHiNrHKZ2PRg/+FIBJSFlSq9CPIZ1wGAMxhAQ1lsfvCcbDwJsX3tt2Twg25myEz8KQ+FllwqCmGb
I8y1fYQilQO3aJZr8jSMzj8hEpVu2eYrkwvePh4FjOkrnt9KmOnISLgLugAEYG84/7BnMvDMisHV
Ow14XPpvjn097hqp19y4klpRP8Rv0vxPmwGech0O1y06O8oiM8mt1200Va03ZPvbJX14l2csuXIq
1Sag39ph4RG6DgVLvwZ901nI/g/p6EZ9i49wlqu4g3rkqXjUuInl9yoX78n81W/ig7HhsJ24W5a3
wSW+3Hmn4R1k8Zt8iu4SGIzOfrVpaT36tWUBnlGqT/O5FYAbqtZWAaVNu9x2MtBYgzWcIHIiApLO
w6EwIB8q5YFx6U61vA9hJLuwSChPBncJRsLsYtlGFivi/6Joi9bF4+KUFypR3502ByaUM2jzQjgW
BD4KO2yi3cecpugutga1QsClOLgkNlmBw9+nqAD9Xt3y76F7VFtKa0t8Iq9zcgm7BBpxllPDehJE
O+N4B0xYDaSUFlZOxZowa2sSqnpHodLJCGmZCKL0l8HceZlewx63q5xl7aqBA/bDqmC1G3CucWgQ
roB4rwKFO8WNEA/0CBh0wVFijdUwdXyE7pP+prIlcXDu5CBCbHfGIQqcP3XjNL/l86Qo86ed5SgE
B2S7qxasGRMRpgtoaNjDUn0o03EhamGSmanuMKoTZNqRiuBwhZzXAa34lP3xDDNoB3Mko+4UbqES
OZUuRTokt8eV5FxbnWJ7/NTbSJwaFVPIc0TnKsBEWLV49CI6bVTVxOjMD+P+z146EbVqZvBlCuXv
E1/aVISdZAB96gUuP4a1phbyGZOkU4HRBkq9lJY4rm4g+ALkc8qVTAxm3En//PiEGj0wM47BxJH6
/Pdu0DxlI3ZW+kRw94Wp+Pdrx3g4uVFeWDtnDzOLXDmroQecVWHU9vc1PHPHrqHXYHNK+cT7Dy+m
qxz/iLHKb+4azlhY3E67lZshjNfB03rY52SpU1OmLrxft9emy4RGv9q4WifKRXj2UN1T4AMgtEPA
W5Bgmqo2JWwYOkJeswzt03FeEqrWTFdT7Zyx8TLaAcfrE0BdNMSsjSkSAeJntIAw23MPwXbZcQrl
ZpF70w45RD7UdjL8DmhutmLR9mlQ9mW7AM2R8qWU9sB+r1FT82RKMvHJB3X7Ur1L9wXdKfpaIWof
Dy45YEI0/1wqiMmwK9YrniBFWNGOIvMIPtm4Jbq3bn6Y4+Gb0Sk+FEi8hTcpHVWBdp16nFeA0QCU
WB4xgK50zuRBk8JIP7K1X9DMeKrBDbKoMP8+eXw+YvcSycmL2zkN1uKHjOT2lWoqxq/K4wNFVrP7
cPeJMVx3vrrHdswUO8dJgGTVfUrF+OmoFyZq/p5iBG9nESieXYFp/CY4Ao8Kc2SLcPI00OcKIKt6
wL+XT6rtBU3kmos5vnP58dyGnc5S8tmjD8GXdpD7u82JgizjJkR+RjIIlaU/FdpbDNnd5u1pMrGi
LPOm+f6liA0I7OVXm1ld3Fla560o65PXTROPk/6wK27u4j9HBRErTxaX7vMJ7J8DY04Aj9PZfxE+
doa+KmEIWfmj60nEoevnLoeddTLwA1zrNLO6PoJoYj0nxYrERx7sOb+4GZzyiBh+e6EbaLKd6DJs
CB1eZy5oOomfq9dtqam3Gri+15dOXihulB+9Ld4J8fVmoODNxlYF4bBuhbeppe59O2agSuS3dAcR
lerjU9aSJbBcE3lIQ5jyyuCkKi8f/557Yj46YfVAdEK9wLTYWRb8SNN52Oh7UhKX1MV+LaHblN/e
htvV2IHhisApYIVQ018hbbwEA8f5kDZ585O49BDNQbTc90NNIoXkxjeoJhgpo1x/Y+FK/gk0gvpz
vMAEsY1CldJQCUyK24wZ8egjB7h4ttV4VQPEuBTgG/xB/cxHrmydSjfRtIWa9RcR4IGIdiwc6hAj
pZ8gstfJGiHJpS62mUv4/Q3cYd5dcmfzCQGDOHoTr0tQRmGSwz8hA6XjU/VEdOU/Bu5MRB6RXBJb
bDTrRLCnRZbQISu/KvJSICtr75E9qccB0gWxPCWVhWBF0jmS78n27p26EnOWJKICtcQNrdm2wazC
XUOgWcRhaA4R1B7ccclaL5GU4je8Ybc8eO7PHHJddGqPweqaTgOFbzo/GZ8ogV4sjcyrAvCFB9dI
7r9ckGOK6ORkvldh4QaQ4hdWxtrqtN0vpC/EOZsOkAcoMYtUyoBZZ/dxni/HaQnZ6wnqcaUmdk/4
cJ2Vwft6D+qzdU0KpCbG/2cGNYt4RJtJV+KUBeuUxkPCq1P26dZp6zf/+sQ7WKZ9I/cMfP0rz1d5
8f6PIE4XZDirvvfldUoawgwijzoFLr8dEbcVz/WohwiV+miae2GOwgvxbR0TXwVY/0Ya6KlozErb
uNLVuCfQ9WOETxxQu8jB2X+XA8iDybvqqVtq0eLyeJnODNfavWsD3Hifg3zkO54JoIWgglCiLS3n
JPQsIEvQdZi5kPutCKu47sbM4JYFyUCNGXEgB6gz3j8bsp62fw6cUsQJGf9cUxALnKwTFu8RidrD
Vhz0kHmH7DOQ1HIvLfta6Rs58l4BZ0CJ+h2W4vVf657V/H60d3REFMlKiJ3Q4+gVM3AJTfMnZW6r
6CCv+xasPIeypp7XEBnojxN7YHTAAMCWAN1+PNpekA9awrZ+11ZPCUcoWlzWRJOcBnccvg6g3iUh
EgLkZCeS2MSHptfv52P7rSNMXaclGkGuhBuzuXdUp7VH/B1sYc5GJmOhKQgTxjGFSCw2kQ5uXhyV
Kr99X7+oH5zXsaGHawKcOGl6CifDBHMLpR6bFStJMtU0fr4ciX8oTOhZ/FDpSIfJqJWlpyvZH4X1
rKAM82x5FWsvWYvnWTF0CEpX1xbRqNT2MFoBIUe7ZfdcuQg+Jn9WdiOf7VbX9N3uzetAdSEd8okY
6R2xMjRtv6q9f9W3UCnlXSmz1WLjTvWFZZCaH545Ur0ojPgdRIK54g4I6XvOD6WaWr9hVFh2emwM
rnpO8eDxkBNoXfauPMN3kTNrSlovgZAUaselYG4xpWE7HVjNKNZ5Tvc7m8SeVndaLWBbrxsQhGgO
mlXio/KuU1A12sFH0OP5kg7wj7JEZO612eIOxAcNt2zjJ+XmudKPl5x7e5NhgTFuZqhSawP182d0
QU6WtBSOQDP9eBdnkCfwTU8hGklwuvwBZ6P3mjcKbhkCV6ztMTkbURS9vPR3t4r0jhsmjClX1AU1
24SwN2B6SJqiphriIxZhVFAWSGxamKGuUnigkswXaTN7yPcpZg/LgUZsvYcMXdGTwU172DcyHIsV
/KlV4y/mhtcUCTb50GarAX+dJT2j2nOWsnKAdT/OK7QP65UisnNAVj7+07Ly0EekGrt1rEFARfPB
ahl71yNtkZNzc5yQWk201gPiTUJIGp17BT42xFwaA/MB1miboThuX9bSDHA2zsSs58eN3wPQ0nPX
kU6g3f2XWcyXERiErpy1M4U9b0z9H2sEYGglJUVoj5jqncxUYrTdYxXPX+tMUIZ9UbbKK7S2xNZt
o9Sjy2SWXZIDVzIBuz3ZhTHdQMq4/dVRG+heG3Yzu2NQgrCVQxpDWbQmuYTxOiDjGgRZHuFNns8y
bUwYF1xzVZ5dZ7gS0RGJMxo2qD9Irf2SbaTVEgtK4UyAiyTi0q9nJlxZ81sySyvCXYAdFDUqHOgW
SZVqpcIA34z2ISxWC8BUhxicKLsrtXWDXvKCfV92fYjfBJXh7JuCeaZ5c/fsjBo5BpVHp1R6wnR7
0EDhZ4vD7lX78H4yVkvvCdHwgt1c/+rVcjUKkEloKmZjk5WhHawW3rv+C0sb2d7eHTMO180Ze8XB
r24dCCep9OFeF6ghKDOpT+WzJ4OBUf+jNNHjUjBdasy3DWRUf5+IlQWi7FnGbLClcSY1xU2c5uzO
gdOKTa/n1dV77LQOImX0p5KjC5D/T4w9OuzrROQjJpzP0DakHebchOtHXiv2YMV8L3t3EBCg3rTV
dZMDEQDjr9itq0h1xJaUyuV8loGVmzzoj2Fhb+n41PCeYDKGN8f6bCwF0o5HAMqr/Eh/OmGKKboH
MYlWOfQlNvssOMz2eicWbpexf5IN63oHdYe0ts9bzPVvPMWGCzN+7ZMHn1Q670N8PRUXyE64v0yr
Wi/d2NNDGRrG43UGJL3LfK54r5cmrEWbGi8cb80NDIA2fPM75HrDyOFHzbVoDT6B2Z5QEtWwomok
zIhYS6vkEhpsjGbryt80l45opUiUhC1N9w2WNHXbTZyoYsCkn446W5Xv/Bq0iKnyj8px0oXkqKg8
U/qK1yFlGhbbkBElr6q7ajTyilgLBa1x4A+ses9LatweCtmRgzXLtAQXebtodhTSo2X2DtUgaDZ7
D1r3ZY9anzqUB4SH+T7ZTyP9ibtvwETvvLyErVdlgXwow84r38mGBbyyBgaGgaMuaRsv5MSwSocO
6zczkrVPlQylWbGvriPr9K0AXYTmWnG208IHR6PwmveUO/+Mmvriqb28RJ022eYuNdPBVylRb45M
oz3ioqgeHoVuAftweYiRV618SHLdfXJ2KxpwpU+9cbegEosDtG3joDgYwZUJwZ3+/lgvuF86X0v5
lBJYR6XC/j5xpL0orxXrKXYGMG+y05BmHm4ziE0H3PW7JSqED4rqosU3CneA0+Gt8ERKbDpK0ZVz
rRI+V77UgN0SV51cZpqKvZIpuzoSOj6+xqTzM0w2ati/3e4FZBR58yWKTm5H2ZG3AYfRdFo8QS32
XO9sRmwjykOUQhB5lr4ipOBOkyNhTjd0lEv+OqaduZpdzMvaOs/LMGu6D3x1AesoYbfzjYFrAFyc
To9tiAK9MWoYMuLesQ4tTeOVK0nB8jqeEM8wBaj5oASOTO8kFjiOM0QyUn/iFHERGLolpiWDeNZm
6r/CTZGuHJjC31KUCeanw+0lq2bK0rm3J9mU8Prrt++9ThGAqWkiIk5YaOpZMQo+LRd3xlfCZ7ma
pc+B5o4k74ZU3VRlTd0Wx+3U5ccwTnsCfA7o+wPmOVkpIRCqBxbVkWNEejvdMA6o7z+5Iy1th72T
Woj0WYlmDXCJ43sCxjGzE9y7D1uGAejaMIpDVzPSKYv9bVx9qgW0pD2XCAWW3AGuCvickiRQoQQE
sP1Bt4P7g7MWDDRJgfRXn3U/KWi8Y3rLZF+0cEQm6rWoc6T8u51JOVLvGM7FtQh2z/mQqW0sNlhh
hL7QPKyMerwrdS0ypOqBdsyVH9wmg9psjBnuN8GnsnktlfdT89+AzaHdFI4eiUUbDIWscyTz8Wtn
yPN4wrtLr6HRe/3srxd6wod7Vqmy9B5+7WfH0Vww6mNHo8JzRxfQBgFZWZR8hXW8zNIAW278jgVr
CRWlP0Yi3pfya9MEHCIvD97Hfy52iT/qkSwGQPhXr3h2WyPFQ283eajlOd9eh/sYTTKWgib7u03k
jnF0XR+ssA8sbw8Rv/R9IlQqzoC6n5qw7nlJ7KFX1zVfi+JcMVknA1rdDvFCK7TeNxqHpUoAq8Os
+F/858nfmwevK3wml0Bt1IhPk3zlUDO5GGKn43tc9fHPWZR7CztUWHjywFKFxR+AOVWO68QkMt1e
GbOT+opw9f+m7VzLulj0QqpkclkYtS8ukiE3RmS181j0o/j/I4vOHj/EAwk2DHbV/JtciedqjCWq
2MorKmlT5GaItBPpq9GvwqiHXr7I6iBLQwiI0JTAv0eEHIpkh7nuXJET8pNEp5aDcSE3Q31mn0/t
8s8C8FD94cZlm7B/JogX/Wc7bmiirXIR1nt2rQnBqGoF2hbF/NgO4usB4d/Nfxy3OHyQ+bSBinR2
yVVg6vy496KoYPyJQhUAWqvGMvA+HAZphOoMMJqemmgkrUdeGWDeYUdM49+9itZM0ptODU9ye60r
HlPAFa6XnTM7ULUlTujmhdJrAx5AhRkSBECROOsKHXNRJTM9ZvT/ULqhoGbIT4/BunhDlie3tCGW
AOYs6qMJVabUueUDwLGwpenhUDjd6D01SvsKkG2JqIc0C4F4/iPiDhvNqvWHBuFkeG0nJWI9WpwT
OX+yfPTi+eImObPkjOMV8i9hmQZiiRlT50ygA0Qej5QgkFoaoMuxUzHMkEjTDCSgKtbnChN5nrt3
njv+g1eHZL3R/lr+zLpbYJoNgANkBG9rCf6J7X+3+yLcBGKTUa4koEB637XA+uPuYF8qqlzFYSgb
EaBAn6NMu1mLZ4BJ4UW6NpJTwiVsc9b2rIZ1eCM295ygi4GDtNTtRvievIEJie7mPGG0mx/d7285
Y9R0D5AaISAdSO/yGGJ9G0lMBEgBoN5INx1IQ4w+GOErcJUWZ1D2DUzFlzasVKP2cVnsZthQwzDF
4VDUlOnXXK807Gb30Gxs5LtkQM0qgj/QZYwqaGJaEjk25j6GF8GPS1iXIhyOE8RhgCShb2eVvtID
CFkrwKfDnisSjCJmPqK7zg1ssMCNiIoN9z0kYxquBn7i2SGyYcjnEQ92ozajg2QzRkgbmRpzuXAv
HzEyOAdic1BL17ciHbugxFrCIWviC1fNqZAXi3DvMPzUojwerQAMuguR33lPpZ0fBUSb8czU3R3e
TJ2+A8ZNj28ZMSO0eicFEDZrrP6Whisel3tiJ78WaFx1XZxyJEZF7BSn50i3WBlSAieq/vZhFi/8
PIo5UMDDl/JRP5tOH4Br6Mae/S1Uuaopg8I8mu7U7mDKVjpfSItZzGK/oOZut+VNDWYsL3Iutjvk
3ElCR1LPui7QAOtd7mxCfwF2F8mBE6P180XpuFWVg8iFo7Pf6QkJYCOTOl4RbtRiQEDyw2LK7vWv
T7l6q9bdD976BKRkRuky7hJZIXPDKiRGG0vmOP/Ion0hltki5LDDVzAarUCqN9rn/rOH8W/3T8sM
71MSTSTXsnfYUfOleLrbTEqkFy2+K1XAlDwuS/bhfvu7F2HApN4FPD2bgWMziBc1Sdys0eGvwuUm
v1gEk+NzfqSxkX2+BIQ7B+XrIYa6AlW7zt+apLo7NalqX7LuFvEggxbSBI4uZofdU0HY8UEYtoRM
n4j0GMgcG2jQG4vR1yEJr4/rPzR8bn90MHMdkkgVrQ+ezwePdL7fyo1A8B+iQXCzTb+dWXq3WGir
KjdEYIs1kszbcd8uoe1+m+VLvExhBH7iuqNR1ntRqeb3uUDY6hO3r/5sHYju0C8Z8Qe1LHdNrXP3
yY6YknGwtVEF//Z15R4deo2y855CDwGq1/Kdw3Ug3XyP3TtBRRxZKBSQ4t8ycb+fKM2R9PyyW1dR
/BsYGCwbpGxV9YnMm8i4LJ9ePC2JfSE4GJO0PPYkGCYgU+JXsaYsZiNbp2LbF80X31U32qeweaVh
GXYRDxMOEH8p11V+186LlpSCp2Ew+w+LzAI22wtRK0Q5D1leY/AjkM2AlsP7IhaD3273JsCv4XCb
PGxlgmNueuMmOIBSoxVnnqd9YwWdgvP8dhimOBR/3zHzaQb/PnDSThdSGx4yQ09jMWq/vcUwGWYR
emLIsDM7mSrj8f3zN9Ij0KcY5NXTgj05Fcvq2UY9ORaKTSLmMweKYaASgMzWSmGN+g1NiLBT9v/S
WGgG08qxfdSodL8w2xKfSKgi9jBUC4rg6UBfE1V12jx5uhhpNQjW5QPkGHcszrKC+KCTb3goSiB2
Etlb+sRyWyjAlhP09kKiFBAR5IlgCeYZbIWlilB1gcaqRO2yDDCbH8fXK+BODxbcu4509nmHwQLC
XulBoKYRtCDSx/xjr2ScHfcVXAbrdzr68eFNuMXUtyrMdxZxm7SzDTSEJtHmBZ83qtUHa6CqZPjy
Rwo2GD0Nv/BjZ/fAa6e0aTkKTzBZhnuBPa+8FZ9i5cqpwt6bSPZCQ7hOi9PDLD1kv8ZljcfDKQ+g
k92PILWqbcZ1aIDJmoUVnvJaxMcfy4ZD5apIhliqzMkHTwzeI8DbOLNowHa6PTs3bT8wAwOOjzfE
Pa7iYszDLdG6LP3YxdxAiFBD9oTuei/7ImUzWOD7GLUMOSm0TIlUwkEtMCyRnFNVvpyqdPiXblYA
sQfCphJpcE/dwaEWWuQBOYgcKCFAAcixJFYH3qmQLfWctlO87X+b0kbwruixtKpTbzPKZBQWlqAo
JVcaV5hiORgRiFQ93cPlAlny4iieGk3cHuEwf2s5fRArQCkFT8R20D5/CAy/2un+PU1V+oMeg5fT
7e/eqvfAIIKvbblQ/3t2Tmnj3OluCkUHgSoJ2u8cuZZBJsqa/LHUV1WblUQqeEO0R4zK6fYj6ubv
GL9AbL2TMy4UYxvP2WMDtCA2PWsXQwkrWQQ1HFtBVkRZMBF0t+jAFthe3x3N9B9T+hucCvo5BNxa
ZnkGeCBiCjZiUvkUC8rlGKOrceDUEHHiduk8wpZD+5XbuVQwjY7q/jfXW6mAtykY/AOGasB3ipRK
rGrxwOYXfARqZuk4LWaeB3XTWa72lzhnzLk60EbejL6DJaFIe91Z6cfx2NNsOr+tBzd+vCBjmuMH
xGGTtOx06Z2ujIWTTLNPyqMod71YECvUUZP3sHgtLzzy8kHWbd3Uj/bUpVL6zRI1BvX4mN08XVEC
GcDVDS1K9SMyWYMrXt2DduSeC1yg8Y7E1r/as2DjBxfOZmrg81SYzn5O0GArWo1+mi6endUuDVyM
CM2L2L8uyywkS1LczSilfYJPj7eePFju80J/lViPzgj9vWZrQ6p6h81Yo85czz226/gXZ3BePVGx
4ov4RvJ4r2GdnWSZonsHIikDbb7Vjn6ofoXp6t8YZhNqcf2bjgyR0N4jwSHi2wcjbI/woVI9JChu
pkx8ZNjTDM2P0hbgZ2wG3La8p0ohj8eOQ3b6DQWOGhEjD1d1iBk5E8h1EYiUikewhbzOoIt7Nbs2
9Qq9FZV2mN6BUYYeRMQZZqACaiOCHC2ZNK0MmVEYNEp3IOyCVPDqxlg3nSjLYFukb3cubjeXqCcm
qtxNkeev/Mowl/AKI+NZ5J+SlxgL4tga2vnftsH5gjgnoliVJL26uBJapi2J60GfJMrgRYlit2Kw
uI2o04ivjmjK3OsNK7EGGiWEEabtkYRExwHm8g5zdIoV7keMZ8jXSbkLMAa8hJwU6FznfvMBSI4b
qKk6CsldNg851PIsriou1iu2X0lD5P8xKhmeMGXKau9NxebUjaALZHwpgMG7lGxTJv+SSV5LCeQc
llr2Va0G/2VDa9092MsPYufbDl0h9dWOEUK9WZ/rzzpXYUD2cRbY9qIkEUdE15NzwITIWhVg3r5F
Jvr3GillVwSQ+F2IIVVvHOJxsnR0TqLFrBdevXEMkpbC31sKpLg4OgWpx40UrkRxl/mOjjgkOj9K
GLyynW3etTdI2T5qvz+j15WiDsJYF/UISDFg3eX63eGCO6c7uGb1U6vVZ9DdceD5YCmPe19PUknN
ZAwk0J56qXrAZV16ValoyJb5PKSQ8c0kH6xTToSm5zdMZmtx7GnQ+Qp72RuOtvqoN2DghRJeiVit
83TRqPZQP08Z9hYfRdTgZ5TkdOJVj3smelLAdvrCEeGTfvlosa+33PT/cTYx3nVA9Pxcuz+sVA4m
Bj4CiLdPP5DG2WNo98D6KM+pWAtlQ8vCwSj+mYg4/aSKfuXsdAY3upz8P8e8K4qsyaAMUkdXJLRC
ex715Xl3i+WY06uam4tQCkkiPYDSGQDcOnipJ0+YCGlaseuNxlwo9QO+cO6m1VZzIi6iaMo3ctso
UpGZL1rZxwzMgqaqdTNo3jpsAxv3onQihJ/xaCj612V9mTP0uuDdXykbHFpPDlY5mxYzy0ygmFkI
g0apq2FtUKtGci8mxU0DQ9HmV2DxKbyn7gBlITJpg0kANPEqURo3LzS0jga+t1ZwrDspMm46epIb
j5o+VXx4c5vIQPudx83vKwUZrobd7oHXyq72xTaTW6F0wqDJ+P6B59CngCbeScD6lrawIQ0MNTCt
HfuIPKIS4V0kpTtWKESN0gM0qw9uctsr/tpYTMctVf9cUoOEY1F7yom6ZGos4nYCKjCBT50sx7DY
6+doql0VMfSFM/DiDnlKaf6Ns7FrZzfm+hJrRLRvU9/Nz4LMS5R5K7Q0a2Eb0+1agoCs7ovZiTgf
0qSvyJL0mtgjSKxU1WkZ4GZqdzHKirIhLkzZDtcfRNr3RlEuITYXIm/3lwhhHOlRFvPNi3nt31mq
JdZLI6rikRxfID4rc5/nYPkmiifFBr3wWMZh/WwfxynsDihPggY3994Pjuc7l+pTQeBq4nzCkYyz
wCESDFsk6Hr0IH1DrelWJx9gpb8WhART2+HsikfvtklDYB3fxP3MIs8U+hNwBoxym6/As/NIl0X4
yLXJdl+RdvY1Yx/bKZt1N7CXHzGFaJGsn3pqHdgUjdvutWRRhoM+UI4ViwlItKUdVwXtYSHi+lex
j7pC144djwi4EFINp421EFmH1kuaCFO3tO9gyNnz0lTnLwE/4j0mhQ8wR85d16jNLbyB/uoTiji/
6RMhA1LXT1kJNvP+2Vgl/9FoTkFIY5iTa3lBnpcLu2FC5ltdNvnhg16rf+Jt4CZUev9Vpy+/Y78Z
exDcz1+W49Z7NHT4ePXeBE9bTUqVRtJuBuNkPyY2kZ/w5693Q/muISE8+/r79gSTkl2t9TVGkG8w
wMFVxVLJvV+cr5kseqpUHLmh2rLrrVrQ5n05AQVmPox1x6QgnPgawsll3uVdsbchvCy1wzp/TpFB
eqpxQnP9iautGYeHdv4kOOPLIiEjZMJ9hkqMfd47ZIuhZoE8M1hoUKO/rliZiAM7mt+053+EUbVr
arorTIzbz2hi/AflXlrKdzH8GDj43YRCpoOGIySebCMSgYngJdlEBa2X6Qv3QTV63TUUKSbe4WPV
4YivC08S6Gkd5EzYt6h6MNAFvHHn1QAblheeLmOVW1PMOC4t+8utKmFv9Ca4uddStY8qr7qLom4K
BBAIJO/8gaEJLNu04S//n3TkVGG4BeqbucRDUfLSPm0CcrEBsaHVnzwD8KtB9n7rzBCGfBkUXoij
CmwiS/RqMomfwLxPMX1TqSFVisceqkFqJpSWhYKtOILQXcPer9x/bFnEi6zyF57FjVqj2fszty0v
3zeebotw0MsTjoSYlyRED7dWxRo1c72aRI33xG5L800I4IMobhd2f9ayjT5dAdB7/KFUgZMH0M8d
ddccc9wwJx7+/jjKK0PvWY3AihzlcqMHBNdA9vnjHESgQ4+0NhuAlbVS12tiqIMAtRV3rBYy8aWt
+fUUQGyO8VEILkGrt5tIZb3LZEW1W/LqhS3aFJRb4R3NoqtiiZFzEr+E8UbaiX6HHdz7rhZdhffp
fpKpGuYM77R8Xg3wP6eN/JEoQ17WoI5vGhHzZzIo/4jhxVi0eLlZHf+Cb/fuUM1vqBCvRq5sew6+
BObd0zTv/fSxDbrC/QQ5F0B1ze7L4nLRMNgKGN0lfJWaeucEOXYNlELZB4jKbhSVhdrbVr5HNQhc
zu+46QFu3UWzkJmXhGK/hsfzCYbNC4EYg72Tv2ztCmzjb/FGtSxYeRVReMpvDvaUfVDX32RuaakU
7lbm58ITt3B/KAhfOx7RdVv6CPSAk8ejaZTEvmSJxdDUcfAF3y/ikEzuL/wg6BwnenvogSrwJt5M
E8hFdVUh/D+DNb0s5Al/A3m6KepO9XdlUGMK4nn5L2eltm/IJ+JXUzorKSVR1/ttcHklxnkDysx2
PfJipd0FT0yLaGm/Hv/RjCZcNq/TII2WapCeWTU2gpS+NoDnTCk4a/DnebC1QEaUP2COSWNor9vJ
vZpdA3dJ3j6ouDn4FSotxvuuHSP5Z/CR6qG4wmK7Uacige/hMVC49/A3inI9vCNgRS1RpVogaZH3
HVkGEzqgsfgi2lofJYvOYqfFp0IQc2knRE0uPZdiTR8m8m9qaznJB4ChsliV++3yXES6Gjb8B1lV
jQdb+zqB+U+ORFgxDrEmnYxpb9czDQ19leIgpxcXY9i0IZGgALXVJNqUiQ7mULyCVqXQgP/ggoUe
I5B64Ne1ZBUq1sLzjIOPcpBtFL08z8xQCpBKVF68qaryH+8GbRTFQ2/ER3OvC+u2K8brHQBUcEo3
wrswTaM7oNObCQsZ0+PcvSTVz0+aSivz4l4vabDifkf18wI33GjIhw5OAqYp4giaAqk4EPKBh77e
dRr1ZTDJcegA4rbpwHUmirCjWtXJFap1h3o4y2UjFSKlcWBIoBqMQp81n2tTXF+9vupxG9FGY21l
llwuIsvSV2CxPLcwYgvKo7Sc/brZJqjh5aLDLRRf37DBK2PmA6Bh7CZgHMNHlTz6kAOBfbhvPGif
+A8NS6Qnh76KpyxMQ27jxUV99b+oNvzlan9BVM3i4iPTLl0cHX7m8GU2i32u+LiohQwAcGmeRiHV
e/qjQ5ldiZAlMTu+n2RogfDItAQ8JoPLSSKBXKSI9i/vjtJbHiAT+33y9eMejzXoAaU6qBjnDaH7
M6XGgzQm3yG3YZ5w3S1sE26OJAbYZipgSrDe6PhxZ6AMmQHYaJmNkHGgHUfuCGyX5qXC8SB7/J3+
0rm6c/V4Xg7YsbEXzRLarg1qrZ1+C5Mx1r2Tc2e2DFIphn5qrR4h7c9619GFiz332P4fENndAVCh
rh6JWdRyMEQYU2X6zVEH+zCeC6qY7t3N4fBCTtLXoyvnzSAZ4CxdENjef84vuleFoFjGgNkeVmgf
PlE6L7VxbjrG2qYKC79vg72yiOIeQJnT2GDwCOKkQP50SmNvdmH7zeR2XemlDC/iQPLBguVvBRJI
s3uehJ0VDeUex5DF9JtfabOs3B3fwlciEWiNnONAerUs8MavF0YPjCOeMEGFuXgvIWZgyrAy+87g
P3yy8TxBf4EqEUR9AO6Wov+75lmWjPL80VKacOdX8S03TjEDEdA2bcVxmUf60yhh1cWZn6fdD3J0
KVwnFoylBnazlnNMJ/sJLAPMlivmVQEX2YSMb/OjTLZFRNKRMf17M2Yg9+Inv0LUzi9VIL6DiHIU
R6zv5/9abvCywvEdzD5ps1V/rKJc68OP8c7zxPAj3dGwBSA9ivQxAlg5Z356ZDQpbmJkYjhLesP/
LdLPAdpooZHCkQ3khYmJBjVMXE9v1rEPxAFUl4ZtqsOt1Sf/ReXe735wvdz4l4CWjo3+HMSOYKp0
DQN5LAqtmy6OvX4gpSKOh9RfBFmdHVFARP79nLolorw5SpYjsAh6B5t+ffUIjFIFqn+aPsCMfok8
TQBafGGWMeEgzDyjnw4QI6jSC9oQ4jYRVYA7OgLmfIthofkoILdwLDvZ64iw6fziV/clLwBv/js9
iTYvRG7yK3J2Yb+y2evqTLFJGGw5/CcsUHZRH6GJN2TKX+EEZwzjuw/gzGWim8f3MDt+gCnNFXxP
N+6SQ6NTRJrFirSZiMZAced4rJZyupdRdrF00Ow18RUbnvPpZ3sTp/kiwDB9J5lhCKuCNjWmiDm0
hF9PpT2rq9/osra2/FrITWDk5JNLWrRsEsYvqfXr5FuPdtRoxRqRCkK+zdtyqfgGkXadpvBh2q4X
61C4KnkIBMKoKFXeHGoG70vtbC8zwujLGTG107E4qc2m6O9wxe9kN1i0T4K58DHx3P7AVgTX+cxv
0PQTxgBC/dSBaj6b3j+vKkLOcCfcM42z1oUe90lAY5nTWDbp2oYesbukP24sXHBEKLBDG7ii4AAS
d3E1YftMzpnudkQ+3nlbogPENZhlN1gk/p0OZ5qpcpQqTapPcBMXj9y2qYZ6YsLISLkf0N+VhOf3
mIMU6FGlPx6T1O37tlbtGqgfk3K372IQAZZiDN6KLRY5mI0iwMovwHi3E9Zkvx6FYmFdi92+Zci+
/cV+J8is9YsKMgx+T7DiikZyv5hrRbkHAOkDnbX4ID6/OZcuu1sWEJQTC73plShdXeCtiDOLHUp7
TS+0FQhykmj63KRNqtk/85xnZnyB7Za1p3ZHUjb//g1hU58q5Rw1M1FkpHDJREB6VCn7mcU8bt8e
uNHKo7F5wa9C/Uw1Umt/RYoPJKXSDtKXHioM9SKVG1nHLe0x3NcCQPlOfRGBAK5/K6LUuHiOW64L
Yd5CdYjGOuTtf5ZjsJMJPchLC79K3jm+T0DmoiLXQoLXsscvZcSnITUEUzY4YBO5ekrmNHnBRP5a
AtaXihLnFkPAm3WqYdZpxN57+MFOomQhbwpd4hXh57Yf65CszHVqy6KysDAWIYwlglZ4PFz/z/Z5
HYamSlvf2/ja40zX3/U+KjF2K9ApB/g9pPhdswj9+vNZIQwImAqH6s7AwaxxWHeaLRLn6kuCzz/t
OKvB6A810AS1HDWZo1xgFh7IjAYHhXjlug8KzIvSR6xdt6jt/ApJL4YGvkuXUwETjfogxWdmQxdA
4J+nhXQpK52TiAvikLUJXcLQYPDj7JtuY9uHW0ec33A14kGSQsozQtXpWEEqOUe1mZWqUGn87VRB
QRflLsqSZOVtImuYbRpszb1pS/Ew2FBTZC8QwTS7ERXq+Sktrjp/V44PSNY7QAHWivcfPPeT1aXe
rP6m1JdiUPwoGmo3fJnuF+9lYEJZGERaNWxo8d6RlROMbhvSvwgl1oj+59dvkn5kzq/FDneAzOjK
wiq1uIS89Zt8kajAtsgqcCdDVTrGh60a9vyURIA9meaiApzI0Z8SrAmP2r6OS2Dgfy1FCYCadb2Z
907MyBflARyJPMhm8/HHPYYN2v9fi5Tx9/pvyNiMnDBVW6Pl3pMvhSNQz80JiXryFtf9rsiyyP6k
aOxYVtthJyXZkCJKts10M9LFCtDagQadW1lLuYThQyfGXe3opmoZ7epusJhFQyNmCY/QXdIOoZXU
BXZMRk8/G6SnLFFyYuHmmXf3P/lr9aBhQCtwT7O2aHXUwasCB6jU60H/bQYaf1suPGkw0hJNwgYm
deBnWD1RDFYtdPtboGgVjmVVN1CKizeSWHSs2dQeK4gCxltEJVKN+/hz8v0waZzfnmw7vdZFNfUn
aKmYFGMKPVVOMSkJimrdP1x+pU6ao5o22OvKXAag0extE8Px3QX6X1Y2MXtGTudykVAGD5ocpeC3
nP1w9I5oo7b1g/DCpe6B3uJA2JMUg4vmfChHBH4j5OnA8vYeP53URsP81k+V0U7ZsbyyIS7vu3L1
fZBIPZ3mpPd3IPYaifdlIKtKIx3i6+tda1HpjtBoo+vgE4KzCbv2aIbiSoRwZNxf15VdhbEE6HUD
FFBPddEhwS9UMRx215VH+ZBFbdiAGiG4BDFk9qwelm6s8kBPPBoVR3x3CpRuJ+QgYkmAsnG7N8ff
5/5QgtyFVaPQrcN8g5gKlA4vSrCnGJJEyPHYpZEkDsLUIt5FM+zio7N3wQw0u7GLlJ1ZR9lGjhLA
k0I5PgdySyZVbR3Mjre+x+ItYBmt+rp2x6IhqoH8cOU8ymRYHZ/A+Q1/ys5+JQNb191L7JSBhK3l
c2NHDvSOTFBkulLyFQPVwEVRwILhbqMfjYVC6nutDIKWOjNhyzVtqfGJQ+vhZHZva32aBudchaKx
Iq1woSpmKtvGxTjksB9TLwf9hIaK9tnv/yvfwxDcRLxLo000389h0eADmp6SEiI1RJonxnF8S9BE
9BIHgarQdVWBI0eCiAyNEfm0+qoCZH5sfZ+wTVpQO9H1DVHjmlzRy7VadrlyKKLSKuYMwW6K0h+E
Ya3AYQ2FP+9dxW9hktPoKYkZQAlol3lvvI6Zx0ubW/OO5e36KeuoGDvG3g/KdBKsKuwYzqT7BjLR
06JAUJojmjRETgIY3t+TC4Yx8RVV64ZaJl0D06wE4kwig8rQkkahM8G1mqxLX0WiXKpULXc8hae+
p2FsU4QWgl8qcJvrtRqsPUlURBsxGRdEkoWMl/xBA2f6FAnMKFpgN7UVN4i7qUhGNkVfiqFtLkok
HA7QhSgItu34MwpTnRTA/4hpFcsKIr9gEunR2D+Ti9sYO0W3Aw7EEhC+w/kARbzZLDtR3EYdgkLk
rRPL9sBsAPv83iGezhzKZchQ9p8ueTO38OUBHZFf5bRUCPVTHz43WGYvqlmYPXBra2tXzHgO1cSn
/cNwXqAe+TJPS1394A1y9EkvItmMFPIl2QwaP+i40zRhKGmpyZsSmCMSoFAJAcP1//akXiSOHkV1
wrjk8YLFfwuoNUZjrTTkW8kSb9izgZNI6DYyRYa7TsuHngxi3RlrNnu+/F8EF8b8/gx+FBFFOTpT
lqR8WaerlAqW7Web/ulM9Lns4EgcFBGNWvm77+vcBmzQS9L2iPVvdHdv3gso42u1tM03ykss+xZo
qzClkNQWDPesrVGFZqBEafHILem0OFAWw0m8Wg2hPFmsKwzGLvpxxPRAfMIuQ+5AWQJTKgLtrmYJ
ApIHOYg7IyYDXaYIqOhyUWoVE9kWPoI8Va1mg3VXEAZPaf3OBW+OJ/W2cl2rnpDMa1VNL10VUgln
O38AU9vJ8qo4G2+ZCx+nuLx9NdGm+waREXne1+CGJ0ovK2ThJXuxZ9YpbT5m5TsBN7NeccehPh4u
NWWe2PQxS+PTVGtW2HRllwkripjwViiOC7TSXNaEsY5iCCn5B+yCFpdlRt1tmUKsDEF52sE7xYAz
fsxKnR35ttqbzz4a0if9VT3J64srAWFKMACTsrrnaQAddagZOZeIZwlgpcuUvr8NEkS4OlQ9bn0s
SC6Ejo5hZTvnqYh2cSwGfm2zDHr3b/R6NKS6LGsIhiYOYVEau4rFfHqpGLTfxjVbek7+ZsKOAMku
+tDHnpWTy7x0LudI9qy29wQuNllYDGbzeR9ag2XxnXtOpmphjiCGO11+1dPVZCjxmckg5jIyhk1J
m0K7jo+LAJa5AxDPrl6M/ddhZrzk+4lDacitPcfCxza8JDbDPLg8GoIjOB/gFNS9b7dGsIEghO7W
Cq9JGXc1Mkb6weWVY5u5xO4WxhGMk+eutDB7Fd+Pqa94OML6XXSMqjrRFkK4Bj9Z815+vCKqK64Y
Qagnyn0ZehXgC6ZqplYlf2yF8KBxQlXGC8PeIag4BFVsCHWk18OCs7EIZaPHqjYOHAipldRAUI0W
FN2MM7o/6O03sOw/rL0yOb4/EBUO3oEjEN/GCirgBbG2f4osKaNw0OYhpGCIdx1qtraHGHOfYXc6
TRlsmsFzl4Uf18YU7H/6Hjpn/708UgogehjBWPo6BaU8xiAa0EuWieZUPHEkwDYcZS63Bn6mfHgs
cLS/mNwV3sM7SNKytKoF5vzkGdeSAXPiUr9KfaUN+8WDv7nE0dnKUwjg9bAYIvdeuk/XA9VdBkVR
U3xs4DnnJgpd90PPOoUzJ93TZFH863FybS08NCd63eNt0QiWHMawJbeVI4gZO7/WL/P7A7DrYF9d
sxrS/Y3STra/gJW1lFcFD3tDmLw4XeR0+UI+83yG9Ts/iIXGDRr77IJ8S+XQj/Exh3YdxPhYLSc8
+v96XnVwCcjpdpPw/j8trkLg3LKgRq00ljjWIc3EHy/PF7gVQIXuPogdA1jRt5Mzcb/8oN/WMq3m
zU36J9JEOJ9nIQyeWItect1d5nIX2knrXjjsAZhZHlU4bteJh0ibnQhp5sqMJZNKK56Yh3tm7q93
p7pcQK7IpYA2ORMzjiV+npdlIMmPTmoBYKHKVhgIsHYHehtfx6/oGYSbu5uG35dWim7aD43zKEPD
EjU3GnuaMUpqOevK6bvlp8IcFtFQ0QfvjGgQmJ8RX9pucOrlKoXavEPlpvW0ubuR2kIMHbX5Ilub
CuJFWMfA4u2I8Gv1f1X3GubO1laO16MGNOTlLelCBW8IO66SALoQoFLPWIrXK1N1r1zKmvc+UzNf
fIupZwHsaU+RE8cKh+IPEBwkSNwfJ+bJ++tfb25Y4ThX/lDNLA+R761uNPnV6eQm9h5HLFnG9mAH
LeL37g5sfxyS4WcbTnX9wTEFmNDni42nPkjRSVwrBsuPYmFY4R7SPVbaOD8N3Abj1hpslcNLrz0x
U3fLNH+C3ZSeK5nn5jpbJeMBkd5cY/RNy0vpYGLazrsChlgSH2yHjFbtWlPIPZZjxwGCI6sHn6tt
aK+Go+UwhSOYQ2DX/kDF6ivaxvjxkfCdXV8h88hfg6kbs3Qeukov8eTtPf9bBjpCTF1F0wdw62gX
HJXkzW5YlXLOTGuXirRjsy3GSNUl8blNQN/aj82mgPf0uO4FYQkZj2dlAfmHNcw9aFfjtN84kfQo
iDlpCdvvhY+jCuq52Ri6bHRaSK+u3In3b67L+Lrx1Qa58IpqcrolQyLqX2KwyhjcXrrzMrXCfNcY
tbYCMc/tBoNjEQAZiuPpECQG1VMhl/gTXMs0aSu7oKFxDTVSpZTs0orHS9ExSYd31Hgv8jpvRhmx
BbnS+eVkvtKN/T+PmoD9i6aqUYTgFY1Zzo7gWG4G4zCjKSo+0FeHpYMcL0kV6Clu4IT6/YEwNxkC
QZVNwymFMZE0ATyeHwNiGwlCloqwlnIDAY1+r5RIoM6UUfXgPKm7UllEQRPQ/+3YD/846CWMNNxL
U8xMlrvfd+OWRkooaSHbDf0KGe8rc/Fe7egGPXUKktK1yfb00uU6W0/iBRQ0+zIsnneFcaeiWp2J
6mAJPWpIkqAM00E0E+QRtuNZRV87tNTT95NFijUu863cgzFOSQjOvzcvpShOQjtwM1Cp9vdK9rae
xGGfcT9eImu+d+sqO1hB2pli3p/myA9Ya3YtZpUG9zVxFrkFcAOJRYzEZ31oKDVYHUGQ6rfYzqBc
Rw5FWQwBHYjidax1L2zvrEbicvIsudv2Kb1VqFPGRj9YjzTuZ7CEKD9rDLAtgX1Ku4LxenCOBrOe
TxK+Fv95RkPJIW16rrptTPG2e7YC0UQuK89MwxxlHnDIefgqm8glaT4Gom4gOvlWXXRkt5Wq89yY
7xzYqooTb5vpZaqm0ZYcSFSvgt4Bs+XfcTBOScKY7P6uokJidm9zEWKT5kaMyCOxQj6q6fhwH1Z7
leBEbS9sDXNM7mH0lLm02sUNTzdoTLh8BfjE8zsZ2migeiLuep5yvK4VqFcA3azLD2h6NJLD96Hd
2S46saps/b4y6VwtXnXLVkEYd4nr3rp6qg0yk1EtRhdx+G9HzadIvPaxLYyfnTkYT30un/Xhp+8J
Zfv7czQnUITFSeJBYmfLji3nPYXSFuRJplKbRfM+49QZF6hRWyravdO3ARfuzQN2RylpFCk9D1RZ
vnzTzDtLegNdMhhjn8F7r73QcDdcHO6ZSABRrwgHvIzzS75fbN3oUxGLbfKH8MPbFHY3LefJ24b7
41SCeCOmfkmrDnySr52lWRVBYs3eTIceA8fc/CrsQg3aDgA1MqttJs49LGutpgYmVVRejAWWN4nM
6qvImd7ZYKMBY9OaJTipuiYRm7VQmKUHlgPwpoJFwYgbwFKu6eE2vMzwGgDo6zpTCKbkvsNEcCx3
9/0P8g1e6tLaimfZwOq7m6p16Eskp0kikzlKh5hjRjUyCJrXO91vTmr6CRhZoASJXJo6cFY9I7Yy
yCqlcYXxBTFfIfMIrYTD7t5jpC8y64tRNaybSjiaj9qiYw/n38vDTo+1eyZJnJTVs5rLGO59pib4
JByqg0dACtWPNj98g4coYB0uBF1I0P858GBUeQaiyMAoB2jGK/xU+G6X1SapmkjqFpQ/XqABFyB6
0vr0AZUk5mnLtRn2k6a2XZQJYoQy50vv/o4VvYR5JwGDcLF44dwvvhRMDJ/GNub2kNfLOLXK5ncO
dRZxKlreSb6OyKNTFK+Tkmx/K8knyxPhVoE7cAl+GB8q5gQHGHb4ws9iT9k8QPH3TXi4jM15K/Cy
e8TZulM08alyJ0aOHACIOr1SZQ4cqsJXH0vqtDX5D/UoO+7BI/ZaNV3RJxEFEV+xU+X64SxDXMNN
SB5qNR64omsL3Z/SCUOExpUFd5d/nGhP6xJAwq0NKW/rmzILi25beu+0eZ5by/3FjKkA+oA632BE
sQcBQTUfws5tbYzIGOAObvguxBx8OJbvB4Q5w3x5CuIc6i3L+/mV+g+6TxfvPcIQVm3eKwWm0DVG
USjonnsKyiONf4lcDneWbD7FGTbyTsexCQLh44u5XMMqPGjENclXcNAPVtsDUyPvVl8nVdJ/QTpG
61NR+JWO8Ae1rnnYqcWtQLb2DB8SkDrhwxS/2w2Lw4TL24zYAOBAJo1hZQM2LW6IAO9TTakPDHth
NANjtUHwK2nGQj4/iiugMvlHsjzSLnDxLIm/sGx8mbTnp6R6rbnmB9NS0JLr0aBqGNQwNJ/+nYfM
YBebNqGvZh9Ld+Ci40Q60f5C+TyjotHqy8kTO/Qrf//O7tYBoJbtvkl76fsdayQA+6Os3V/PPWAP
LSARJggQSTY6LlS0/KNHkqrVdXjJgXFdyGAlnKOUvm9lLqQqIkuMiR2hDxhpYyG6Hz38RKaiw4bR
V0giqw4Y2xk8nYmiUi/E0MVhqURC/MjRlIDbhQcUvlKb08jqIwnJY6Vpx4nC65WviVkLOVxJ2l5U
dujdOkjXXuxNgi0jcTuoG8E6XoyOGWJED1s6o/+Q5sVAJa15R3087KvYJiAuQcmh4pn5uYXDVh6e
FCBny/YdqlQfkRoncBeHTilUSe6m/7Dw9g5QL7vuCbxNe3ianmT/QnMa8DEm2TK4RcW2R9KUuen5
Gr0Gax98YvSJZXbE0hptK6NppSBZffyERNUUVfFgtcC0Y/b4DYWkIO5gXRixkbfHjy0hqvNkFM2U
vSyvwojgE+yz9jK4KH4lDn+bx+kwuOLIQmJcXulw1A8NcAqxlGArbvYe+4C9QFc/25R4Lr5Wzp4R
jLPsuuO+yVgvXrUyk3L2EoeowYF12mqh+YgML6wm8h3yewePqEBaApIekvtSVmA7wopRzR+ufcbl
4uRTEh3Q02cq/3dnfKt37ZM0z7bg2UII3iSm3sbXfnCBlGQYOlp8caGZzQsmq56T9u/B7gySKgMK
7MeUNW+wst6S56bW5bq214aU34DZq2AT5HJAVxJUe76Xzg50WpJH9n0IL34nxL6chUqVs0ZfW50z
k+/00beHktrzcBhXv1r2tgRwVZ1TmBaPpbEe2k33fSYVaLioHtiJYUDtJKnaUjK6zgjgrWvKVAXd
Ae5bLc3RZ5eljNUDQMVc50pVqzmMMLahaHx9n9C8uBmUMCI76lj6qIpHqsGr8aU0hMD6H1OAnjSe
cOXaP5qWhKoWkxiNif4qr4iqaFh4/mhRSSsZ9Q0Dtn4n1ymP5xxnY2xeDqItfQtwgEnIFLnt7b7t
KY9igR2Tvh35N8DWCSK/iA1hEIv+5qKMoieiFslpMADFcHtuYZKKN5hU/Zcxln/bFbbYMqO6kQ6U
XeKLlDlThB99/dxbjV09v1DgJL/hjHW00W4KGXqC03dzSYDdiG6zch5W6d4RQuNCQzQKlWjO6AHU
XJGLwQNVXzgFoO5QBGjfO9hM2yQw1Utynm/tBodATagGDHpVNDnhyb+h4Wrv69YfrRXE5KylQvsF
cSnk8qU9zneQMiFAHUFu3FORACgp50DXN4YTzhrBKOn/Zv2fvI5WV7NUE6hCKInTvz4UYNcBW3Rh
hKiFcNPHqO/5kluXAQi7uG6tFZ44ZXwTLpXECu6Qwo/8vpCxxs1JEB5qDl8bsGs8VznWioOx3RvQ
ke/e/o2I4ZREWBOMu90F/9iHrQX6UCtWnNzKKI1CZpD5+6uSRj6dJWOltmun0DSXb2srXObo+feO
EkIXp68G0NYXnFBgL0ucKi8AFkLJvRlop6PAUmByxlbjrdTE6eEY5BOAcp/u1LvQBTaHkHnT54dq
Z6YDLJ0AXejEMr1hZpt94xJAKYMxemAxGuZZfDNb8DNkGI1nM9oz4D8lcSBw9B/EU4GwxiRLgkSp
iAIYFCV5NqHwywHa5hgXK04lXM+L9juFcgGRqoAT4aZh8sfYYE5gs8A/q0r9C+vlNgWeYd8mzmF8
iLLwRxMDeuvZUwk6v4DAMZmTfo0BP0+abHobq/5rBUESUuwkOvtif0o0hlh2x5wTfo83QrwQcQcW
YTvb97HPt23JH/lLACTlUUt8hSn7E9mBVGzFYht0/IylhcFGTzu5H+gz735+SQf+MxBVfatQ9owG
09COVKSL+t8uwkmDri4zzsTJFGEQgDhjeS/t0vL+UlPavMKbj1nfDiq5JRdBj9PEZFFJZ6cG7D2C
oxRqjUy+dpGkL4jkNi+Rpmf9J0rN7u2Us2ngYsvf7UTaOKM7zlo8qBKihRTY8g45DKVg+2UTBxP9
w1eKMVVWwSgTygnfdIrVN56js2Cu4XXLAz33NBTTl6J3NEOWch2FN0skpyPrD5X7IlQXcgZlADvs
R5n70N8zzKriB5b7JKJX1k7KUkWp9bBceEqkBFSFq8Zo6Ot1y7jNLDCxmeym4kqIyLXNXvy4jpwx
6XJVJWMhJVSM0SLMSHCq15GWpPHiVMrqA1rtC/z3WWL+4jN00lSPbLaMP7HuX7VbH01TVMWa1BVA
5UnAy/twFnkTYSNq+51I0l7gDM6ba4zmD1E7GdPmTK8Z/vATxxxSohvQdDNIqCu6YGb3sHndpzBd
QywQVDrw+/rnaS7d/TCRFeyshyfo3c1GLI4kYFyHdtQzWMM+0JBZJFharvPUSxOA1zXzgOVfB2Uo
2NgQnskobb1jhdr/XCZPASE3WFegExGshjYNBx76lPXxV2CAcF59/Ow4yxuh3NF9oyd0H9CyIfkN
qmP62JVdliBEWBt4pIvNKsu9c30Tg7UE7a6xm2PZAKygkv6YWvJI5rbnjFN7Z4iRvHNX67W1luU1
Np4a73zYtTynIfoEiDZP5Z0nAuAvWFGlNfxLHfdQ6jKEgzzMkVL2aaavk04Npbu0URdRUIggx3pO
SoONj/Z1IuNsWJ3fxIV/QZTMWzr7+HkBsHEPBDfXSaMo4TpKNliGQWNPeRDeuLtbYk6BEPJLucDw
4fTrjHMSuqB8FEwElhQoQshdrGRUrehOan2QdXmTjPd7Sc6/hzZ0oyYj68b6nOgMlD8Vng0P8JLx
g49uHwtp2QlLsDbq3Fny8ng/YWjYgw8NrnQFeHdnqMBmgUFNinDYYDm7xRFazo1H9OOxKn/A3qfx
nMQFj5gCRbtc7481Pg0WYpci2Oie/CygyO7BwykxU0hZ4zybTo9pYIjPFQTTpEXXWyO/6jTrj2fh
BAZF0QA07c1YLJk8Qbrx6M+K9hMFt9KZEsKIxwDqelCpIaH/PqZt2Hk4K51IsyJ8TH+2l4vs7jqt
dlqCTZ4w9uTMXezxIGFvFLpt7W2faq3S8MNLyrqQAF68oUWnruOdE82yOJfQCQnGz+uaAIDzogP8
stqSbvX4TS4QE2Hk3r5dBC0syiyRodET+e7o0cmJLaoL0vP6S9kAL5hYeKmjLNDEMD8Bc7H/xTzR
6UxtsltAcBgEc+HYXb/Y4xO5qaecLoU1VWM4JqzXZG6XaK/Pjxzat1E0LFeTQDPtq0rZr68snInh
PJsdSafTir1j/zZ2eSshA6doxW884NAhZF2+rFPqYRldLDr+bnsUOSxIyZnU5tQLf5LHNplASXoB
/4POLYagz6a3k+ZnUIKH2AuXZFZauHYMV4iF8x9WlK3CZjFUOVMWbrn8C2f2b3DHAJD6w2aB2khw
8Wq1BhmDhB6gz/tJfQPQ36rewDIcJhACbpxI0NVIBJI7cl6GgN3Up+ZdEXqcoCU8cl9RnQG6q1kI
XN0DbRP9ve7stj8Ui+DjUJ1VsZBESxK+R/x82e8DF8ZGRyozsGKuDDqGcP0iH+n8WmGxsYf6C66K
dPiW9246O5o1tUimG6haTZ5ZD3J2QQQYZOqStaEj+lvnQn+t8CkyaPXPW/WKvBMO4TfrhzQIX6FL
QhU8Nkv7quBFMhwC9IyLyKIIk+Dmhh2AKhXTjbOg5RwDgbvaERT34B9q8Vi456EieZygtVVPP2p3
F96gmmxRY1cuhEeupfJUgbHkhLc9z95kRpPJHiO5p0yoBQMPFxZPOXqcGkNeLHINDYpmI222TVrE
OnHcSw0v38rOJNSD74sWbVAzmXFRhmy3+bQ1w/UWh8mX0uTRPHjtSgnL7WFxeN06UmTu/vNiRIG1
hpxGkiGBvGtfCBdB7IsKGZz9Hv1Jhe1X0dz4DhYlu6YpdzPfJc3/vlzMRQgKQhciUnO3B/1uAjoJ
+J+Os4uPTo0/jyUpc2FJx1VnMFY6GZ+4XRPj5Yc6Y/21+PEjSBTzIc8C+sVCHFiXm86BZm8O5Avr
+hICXvztjsJrhaJffWu4QH9NRW4zcIqtPmpwx5716g+li6Rcdg+698TJjd4kMm/4LKrI3WiDxy7q
0zUFRINKAE+oiXXJGdP6YZf8Xhv2RHDwB3J9IOrglHqLu2bN7+N9Sp3bsgSYOUDjSzO/DGK/XDqG
d3td4E/D5aeTq/L7IA/C2gyBgSR7rnTJJllRh1HKIztdmLhBLH9mtg0nkw6m4nA9zxrhcFOeacYb
AqdYjaKtXTnz9M++kmFoaUMPzWtGqunifu4l+O2kADFNqMHRftPMxYcgeN3JPOWjQmXE6GNiG+3n
MdxSfoTA4EzasNSwZwC+fIToyWxu23UJ9w1K1vBTOQKBifGYtbf1FmKzGzVegEOUgSg466GU5nqC
ViK4EVSP4TiBqDfdBW9Mv50GJDBdY5r8z+EfCGkE/eR4iNJD6QUEZj43VFQ7HCOpNfw3HPG0Mv1r
LHOnM7++RzEP24r78S7oHZv39+nXYiOCzgbwVcXjp8tqRdBV+tZ7yD+rvdLFNSzG/ntExzCakE8D
hEWNIOD6Sgn5e1TjZ/cCNKkVSuR2mbfUCz1foTeZ+GV/XCWr+7rZNSXt4bwpsbtNgTxfMaDrLvGi
RoVKUUOXQZWyg6CE3bsskeXwPaFSKC84mI8BBXXLFi9MOoRdDZ/cddUGxwV9MXk4f78o7KiJi8Wa
VomrWjqKsw46hy2S9NtjSuJ3LJ1VxyhaP9KhjwYjNMMf5Sdm/GTmPUm+VNgZ84rlfebNVuUhKyBw
F7dGJrZwpnbHAKkCPONj204W6fkxyu+l+vQJSFolAX2woiRqzVCrNj+LQvyN93awWLamUU1soNjq
rd3ZJ/J3Z3xLJ+4ppjsaK2+lB8pQOqRc5z6S4iYQdonSnL5hTmV9enU/yybQZ2lqzvGD2snmB5Wt
LfV3y/s+Jl1Ifaup/C//VGQW0wahgAoqNxwAGe183q3aQiG3tlehOx7MqDhzG1m+R4aWpCq50iXv
bJZhMTmDS4l4//DhT35CMmc9X0z6mEy1R9eDenZ7rYnhPhFRw9cGKr3tGGtRfM0LthboSwm3HURi
pmcbKIv0yWjS9yL+93GvQp0g/wAOOsO4y8Vqq70Pn/v5Wo/+Cnn9Gns7Q3G31ZSIt1oR1nsQdO/v
rRtHPFmZ8E6qOj6lf91mTnjkRhZn+ku8+NrULdn0Q7NQkaIxxsM8LHO/DxlJxOIAAr+Bp6qqDjGz
+nw3r6Cg/yyYngYnZ1tZeIog3Ooiz2zlVY+ElXukhdTk2pSzpxe/REqmE275/fPvAw8VertdBfxB
qBm2vf27jr5opP8FZeBKE4HWCcglt70mn3fPTTU0lht1i/a904woW13TnD2z02ljX5xYwuwRA7qY
7JUyJxvtANBEjrXvvHtsRCgm7OP69lh7GjyTIPyWqx8hn5pUCvS7+BSSjcY49LR8RWfTUs68OPRz
Mif/TxV/y7aHsOV5Jid17ldi4JL4RUOh1WyKttl5jcxms7vuJZM6xRwoaK3MRlPwPLikBxQdVxXZ
iqyjS7F23e4ISXwa+zfkqsg2cRStKseyvu/mdNY2SFIWsP6D8BjEhQ//Fudps51EjLZ70aEBPP33
vSaXLWG0L3JakvdiuO9/lmtLZIdd80drcef+PrlnUF3p42jIpsTcQlkUbqIWYgxxSpxKanRzhEZa
IRrnUiKmZeBO6DGpAGBTNPpGnBvWFxQKNdIstWNOO1uD2gFOPmVQimQrc9qVzQpGURHirweEXpPE
tBcdYiRPdLTW00tDZ+zr9QC8RfMt+5KnPNoHtyXMyWrIqxpmiXq9Rj/3MQKCV4w6Qt/qxVqJaV4W
r1H0CDvnaOLJUp9mzp959VmDR3tptO4U5TyszqHRzCAvgbuLRsx9ZY3BF0yC5wLwYaucB36wTRYb
XCc76BNL1J4YKN0gTCNLKmbnpB/XIqmPR6ck9p1HD34tsznVbYJ77qVabS/QfrNBxB+uIM1XtuvJ
Eu8kbomSWv11RHF4PFjnaI+GmnQaGVcFHCpJ3UpeISDb5MKY+gwWNljtyo0iRsxUDrosi/hACTbZ
CAaSKj3rz45IJdLh4KEV442vT8sK0hBw05dbg/uEcWCiWX1mAnEkGjWPFh6hYLwc+NY30PsNa/c1
XeyJpVB/K27HWhzdnvaiSEPp0ev/DgTlsGWXPPpUrjAqNrMNeEk6SCOleNZJ9D0l0g2iZjJJ476N
gucVRlKfaBMf7ZvWrT5bC+HrHI+t+OIzj4y6c3LoCl8HvcSrQKrDUbKSx3Fy/aHbLA+7mkl00Wxe
cBLzMHIWo91tiI/SpRZsG0z2qa8lV1BfZKMjq+/5YqmhYk8lh7aiqavU1bVlG1ve16LZCUS02g6F
PCKTkI70L1tBwSxiu8JD+uBywPx4Jc2TqTXdON97BYHaYky14hKETgk4D4J4yNutMq52dEaKeYAW
QMxwfl75W2ydaZ1P6QjJr1CbAHt5Aopz5CvbtkYY3D0ZNakWVxw7J9devam8GzvRZ5lxkDwj3++L
yXY6Kbp1k/O/O48SHrL8uhHjBcpg/O6PxWN/cTOnoM0lajH90ekSJGzRvClV+5307nYalD9opVP7
XK7LrCn85cLGBSOTtoSszn2i9GP5H2hoTJYHvoNUrWprFzlM5fI5jdn03Zf0u+FbRBjKx0GJnCSt
viW8m9BzcABYZaIw8XEW96CNqcZUW2HDAzEeOw5kgEpjFdxB5tgrB36MdNNIVYhbaWqM2P9N4IJc
zayM1RXfAsP7l8SbQJzpKlqUAlz+Gvsuzm55Og4UGxxRP7Y6VS0S+Lgzy8b9RbteMenkPY6DWM4S
EQF0WlnFON9mqO2DXbNMSY34mLV/IQNom6BhHBoE7pfsaYGvVQ4WnHqK6Ixn1npRlwqqUbKtqHju
nfrGcx13aPgzLqVfuOQ52ggNiPmkLcJF28xN8rYRY2oVIcof7L9ucVetqFu339BEN4Jg6pYJHPgB
pgYYl608goKCaz4cCWZylGtG3MihV76ZA/fZFDut013ji50x87PT0lcSMNbDtSUrKSO4rfEEk1ZY
RAXYRi85RcJ8TaXK0N05QrXd4mAulsn6JgQsuo1Yw/GswmhHTq5BZcCw/4khmHlbZSIdQ51oex9I
RRimxTx8l/3IwiXMDjYMmk9RmnpB4kjjxOwMObqrhvs/49ffEiKWU8feG1E7SDotWDP5sEfPwkbi
COkDKrkSeL9/DNvQQLKGKP1fwLlNCRSQgPYV8O6JF3D3hApZU5p4Cb4hkhovTjh8bPwHxAELLXUA
3I3rJIoe6AGMG6YCO+MqRD7v3XNac5ZCrB6QXh4a+Y+9WC2b7HN+gv26yerRDQ6PaEo7YgTmpCBc
Iv8axkhGX5ozJfuw58ci0iCYkTSAfv68cO6Rev544/rSjHAA0fyjuAgY9epI/P7ol6B/fuzVm4u3
ehxFpYP/dr6vHHe12jhnoCCHsr2U5sjgpkhhi3COnzhZJybi/CBvqnxPAb5xWNLuDJ4+zpJoGPe7
nTUJbIRfdXAyPhZ8XwfBxCQC6ZIryqrcCIIa7wjP3XqRqvh4rslK8pzu9kfs5WfESNdEZ4mRNghe
zyUiAnfkyjSo7kCYFkDxWVJDA9DZfwj6r5n9d1bTdb1IPSAnxymxePGXCAnOOe8fA+jgu78TXNbw
9Pe3/mCYclmS5u2yd6cAF8qY9WHxRgiNSU2AHsDaF9WU/pp0aJGsYtuWDvviZqYN+myy/opU3jnK
fFMrWOgbOUMxIAMz17ZBjvy5ZCbyZMagEV0ztL+MA+XMLlN82us5dy9+GdzDfsBDJRV/Gu5KfEer
EJrW6oMASEVDeUeyxWrW3LbAk3Lw1rPt6Uo+2SM0slKNT2hMQsmCaHM7fnq4Zgkm+GAo1iKzr4xC
IzGMWRlhLAUXRC0tC0ekyvHp3ZC3d8Cwk6bagSAnXbvkyshELmj2cBZHlCDcLJbny8boKjTcC67j
b/QaGgO4HAiSFs2i+PFvv6V3SYUriFEdxAvUBBp4XRDiab3FY+eD1JNfGanA5PjwYdxqOnrSD1WN
11b9h1qSK8zsGirBD4bzTV886vY4wy29puLYM+s5ue2Bf6mjvSkdzZlAhLbNnD++ZElAg30Mjlfe
1f7+FXt3lmm1vgvdROyGgBXj31w1lHmXtoaxmjzr58PK4uUN3uxmR6oABc+yod5c1TmA59rN9kC6
ydRkad+4uOSOvTpht4zkqgQ4k0NQ0PG+Sk+15u7foJOD/ZHRPvDY6AH+2cfLmUW7wKHklSYQjZl/
JJMDeh3fbWuYRp/Uh6FoFbimVZvAGqL2TYgm2BQh8uJ39HIZ0j0PfBZmtYAi1D/ppkbQWfSOZcG3
4sUQzNMuxP8w5ehTMu+kwJ6Z5ZjHNDH8fI63WCCCGwmhadeOu5Q4Fl/7uQfEMvzHDbg/S2uM5Udb
M14apqTkmMnSqaZUd4EHVwTKYKWLXS7mSnhtFyYtNIfZVGxqc7TTK+Wq5gqa0o/RO2fFMZW8WuC1
ccLHKBOgM4z+p+xuHRQv1gvyBcxzw+UCg+AkF2iqpdMOAJxkPSxZe4sRnBezXnUlJPdqp4UNf97k
739Whq4zhlRfPkq3l6aR9q7GCRyvhsj5vmY4/VGQgeVyE2uXpeQi+8ta3GISui+MjRy4XVkze4JV
WCxdy3UyQHVfjICfKGym0u6Y1wUYlJXe0gVTHH0j11XhHH+/EySOvCn8hHcjkbxkwJhropkiW0QP
8VPiLKWijd54yTlBiSXVmeiu/IeLCyOCCJcTAEEFM5A6VQOXWxR0qeQLAkgn/bt6no+P1QOb/S/n
pP0HQOBSSCHR8u9BC9LCXb1dqy8y+1+B0cmvqB4WCwNZi8OGK/4gxWcejVWK33s/0w9ka2CZbqCQ
oXxCobLYPST0tibsD2LTOhOwNmJTwS6tLFoqnX3VTTVaYS/YcIRHd/I13KJ3NsrL7v3NtPvOX6hr
qUsHNY1J2e54qAXjaPsCF7vebrZ0DLUxHL7sMeayVxbvL3Z19sr66K6X/ZGuc8VqYDn0xbpVaXe/
T3hdg22o/k+bJBaybe7/qaJQ+Iw2ilieN84T4NRX+D23quzGty4D0vTZjg90LhlD7/T3/4hofL8O
cTQzbCKVvEX4xLGiRrEq3O0FiGlBQbDx/myRQCAYQWVrXSJqcFuU2dbjvrznsW4mprv82HAxku7I
yAtcnxWu8T9cQg8ZM8uTcm53IsiRPFLVPWXDubKmW7p/qf+sG/K00T0zlcCN+sANzRnwhSZ4KQPK
Iyt/utFs0niMLJ99K6IIC9sbxEZbTdXN6P6IgrIvoti9ZIacJJeVGZ6NrtpXYVzIwUCG7arMi8L+
xZB6IWMTXPgt8lAkOnfkoPvvUJ0qxxUYLVQ45IXUZs6+8q5Yq2C8Z2iNxIC6lfB8t6juMK5su1qr
ZiIsxSTh7EoAVkwSGFH/GLKm1wNTZkXk05LRF31OAqlkJpA7HvYL8MCMCgQOBe9kFIqJF0qMWJ5E
HWIyB3T0Dc5TaKGMWk0Kiofgb1Hn6PRLqjQ7FDym5aaB3jjCb8Zmd95Fa/JmVU5OorUUxbJGVnsb
WL0TrHh69yuasnc8qENbBMvyvWT54r1wu3468B4LLA71/n1gI6CY5r3ZIiHcnSZO65Ydb7S7OYgu
XsS30Fn/8nc6O9f9lBYaBIiycwMZfBCC1wTe7KuYt6yaQcCwyNf4MZEEDbCGewBkJkjGnkq+QSds
Gsz52JXzBWYqye/kqrwlPStXFhLXeZUaOP9V/pCOm+H52Lfi8EsvIZszw+C9myXyIp1WhxZTGR+6
nsmqrioH+sCasvdOUP1m0pXr8iUuliBGREprJk4gl0DRO3pK3QLQFZCX0DiqlNzcBH51wpK/VSVy
MvUaez8+xp2zcWTQyqX2ny5g7kh7Xi9xy4Za4NAUgRYd/dwX9kIIrZppntET0+D03CtNjtWpBpjO
L+ReO8QTUjMdWNDZQyS6b/hKSFfr7B+9AC/gdG2dXQpl1e0RV4axMmBrDh3YipXjSn0D0+zA51QD
HMWzcq9Gs0q5G0edIoAiPKqQ7AWVSr1imTt9YcqDMuGMz2uHNUafVJY93WxPHA1LLk1eXfTa2vEh
adW00V8ar+TPS223qI9IYJYYv8PFo2tkxZCOpAXf7q+25j1i2kkWTNC4G04ER4PEYPdx3dHB5jWh
okVGZm20DiUHcQaH8j4AcOiqU1G+slS3zYgwCWiNjYWMmoMHAGQLGqnlLbRx0aotqTgpdUUfrb3x
7rdLvxFbEjCY6MlDTHsqRuoSZjCv2EBIwa4PMyxvWaCG4xFaYwEP7+vvj7yYiL5r/dBIuVpKyrzZ
Pk9GvywkIxC8MFo5c84LZGsIGuAw2kfyWdf5i8sY/SRPhEf8mRvwi0D1B3WNHB1sGUr0HPQdrHx7
9ZGs+ef3tID0dIlvTaAgocq/xFulI9nB4i9OpxdF9bBhxqM6uaGLKiaHU4w6nCVAFvc8PThlffpN
jK13n3OZ4Hc7fMNXtmCQMPzzYt7oroa01avuYqJKTEj257/TxsgYudgef3lXJUZOGycYhO0V+rLz
acz3QvY8fec7KMConzoMhovs5+/h8Ghj9LWJ/nLNmGgUchAJibNGW07CnnrwcNGmBhfIAgHBsNM6
t/ov6YpHbRQoG0jBquudsOi1Qmo0Iz9JSPRNnlEOW9DWVMuu2V76VhyMCguzKHSR9wdJGlg+DqZA
Z5JybJrtEts0cudB0Q7o7nXfWr51q/pSl6NGWjOi9TGWro7xI/6PMx1ZvSsoXSm9qcM+g07nXelK
MqjrrDnOoQoFvZDjb5WHaetMG99lCzydtdP6UVeJstp6Yf/drjkJPNFPWrnJf/LUoCyM3MzFoXEU
e3CtZMEOr+8KKuSY4ZTvlG/HKdT6Rmr7clYLwPSCxK/2WCFCL9nB0q04F0aAw8E5mxGNQxLXCYS2
jOM0WHL4HZfm31zIu6xX3Uk68KlmSEYsm8fvGOFK4sDd9Msnupmm3udDyGs7gKRxAGGWL7WCwO5i
0pFQF2P7s9GISv4A76z9OD48hCVJzdWql/eBLEZecoNfagusA0Ho2my+eh0xYF3UMYb25tpGteY2
df2GjKGr+4P/wDubDKHmf3M8jJDykCTYkeUPu4Zd7/boW210+B8XFdpbsx+alJmq9iYFLpuJ2Skg
pjJ7jq0bwUMu4nQ2sFGxijErIYw+mu4ZarfUBSpPUH8O2swL3kqKWodyRAjRto2DpcI69DnnJt/l
RXqoufuiSlQ37VCPKgpEpF4FumYvRbLx9estmAESXI5r2nLWYT/uZjLA1B5NFIxnVO9dnd+52Yty
6IbKaS2I6YLGqg+5Z/yZ1ljZMNjH0Pbu0Ia26FShbj12pTb/j69TyB4rwJrfjnNXXyei6ToJfzGA
JbdJYJJMOipLF1ASYD15WVa4WuI9QixftugaEed4+fTK6c66uRcgZRhMLIx5deoQFJwbxhPagTL+
2tBtXPBgRqPMyylgbDmiEU7qDqoiwEbYJpOoaWQVoEZaWPkcJ8fRPwvMQ9iCBUNKHhR1pBEglqPf
iYU38WHI1jFfgAvtjVvaTUQYUF/tWLviRxlg4e3GVowdQEaxWmTTEedwkhvrMrPQgJXE30FWkoV3
snHuBRrMVHlwZUmIDuQ7SYUbts2aXs8ux+PsMCFcvPmn2qwVOpE48GRhqh0+i3C5otME0n/zl7WU
mmPBCR1tXOXNlf/pEj8KzArq/36V7uoBI1VnEfhwMupvozcxrWvy/tFCp5GNlDacvClvRN4RDM2V
dub6d7i0VywAm1+yPxNTeCWO33qUblYSp8D14WQ45RHJcuna5/LphuG2neNGGwGiWk9LGo5G5RDG
M8FGmjzTixcnTkC0yobGMQJ9VJe4VGeetRIiBX4nmiRORVvjfuw0uDGLNt52s4u0O8YvajPBjsiM
EGuah9e7rCbFZHLUkPPAkYx8KDb5+gmG9+WfJf7flN9YLZIw2Dh0ay1fTy0p7+9HsBwqznzOuqON
JojJnyQZeUxUDYK7fO+RAsE5D0lhQXg17NbYkSu/9nzGuc1AvAEhoaH7hEFGHxmD7AEsKAEvIHkR
Cu/XJuhAlzkGvHsBK9RJl4U2cuVtxV6K2k1DQFVnvwcTnuXCaF3bUbjhpveWbSEpf0oNj/q6F2Ry
qAhtSsSD71g8kmMoh66+jahcxamf895iiJ174mwYtbZL4ENX2yxGhMrWhAOlav3gBk4KyjYIQSDI
PJ/4k2wZsCV8hCHvSpZvOopek+RP1VXMB797Q2WTPsvTLaDX5Dfj66aPJfWUHn0lFZzpegfhJa4Z
o9D7AasB98nW3Q9JpyPKOvRZXiCBLdEKRi4QyySmPg3k0VS7ucPGGr5BQ12fVg5RkObWoCGho4do
bY6nNrRtH6GEFToSC5geFViJOe0EMiAHZpsIbeiRrw4QFJOSWjDO2eVKaWEWsaostSxLcDnaN35Q
CBbt+duZW8behjua2EWoOKfsty++PjqISxiEdvOSPLtgiKQZPhBo1l/reOaWj87v/zcQFOZVHSeV
7Cm2xjj0xcBKatPjlD0Z5fNwEz6i7WmwsuiKVIAwDyyW8SvdlnuUJyIidgEqzSb76JJvj0qlsfzm
UZUJAc+2+JRQAewKRtGHF9palvp6UTBKvm2avFQ33yPyW6YKFly5C4/0SxMWJrjop4V1qhrWYZwy
1VUX3+kqrHljfE7KD/1TndMM2xbId2UK8VipG1JnEDx4BWiMqHiReZh+fFvZMF/cSqHvmhKoEAMg
6uZNqk3LNvucBphHOe4cGwHlV5/rSk5as72PE0sBI/ufN0sM95IwKzwOauDqYNSJC85K0bLm9BsT
DD4XE8eoYSO10/fy5I/78KCXP5GiUoXsMJ9OrwXKF6If5ksU37BE3NZrn+XryVueR7GqR86pJNgO
0U/GewzprEyn+qZYMgkCR6+1qGYunxQob7qgCvojwDoM2491XbTkb0vtf7YNC0pNei1XW2rjnY4w
TVPEZS5QPuvHIzmyenlg6aKe5r55Zp8y4bCxecyEikdQPImVdGvp0EG+tUa7tukme8P9mPw7gk1Y
WTuw784FPECGB+zkvC2SGC7WqcmPIULSqtN10erxhGgO22qOVL6w6QL2KJiPEJVszPPN2jrkiIBG
LSytWloyiqqhOLWH5gtc6jL5daWjwNLTay+7Z+24eN6YPScM3ZuJgkACGew/WUyiU9PBrbE6EnLk
FO1PJyhZ7DLP4KbqBjHX9fYHKRbJIj7tibmm3fHe8DeMWjw/KtsY9HZdb+/YGN8ndo6yE6OZmiaz
BDlyjaklJCafN4poz5NVNcxmU7lqGOBMtDnYov3rw2Xii/dKu263uI1lc9GbP9PEXstG65LxSU1m
9uFvjKDHqZ7ebdWgpFsd1J+gejgomezHujcJEqFK+N4IPQUFzx89aBny3OfX51GcfBC1AP6/1AMK
wlIwZYZYEkU/Q93KTDUNEwtUu56tsfeRIUThOiq/iQhw/pcsPihqLFdFg+J/C54ccWW+PxFdKEDL
KUwd6zcfywUI+cfUaRrTahpfTNBFYSSSfET2WKBKMXSztLprnciGxB90yxzr6yNnWfe750cyckdF
5g2HeS+9gR1PXDyDNctZvMHpA81DHJiZ0PViw/ihZsVdJzhFfxmirdRvR0SAoRKDC2qFCPchFtQD
wEGZyIRkPRgTsdCaI6D2fwrJT4i2SO6JQ2DlLez0/WQn2qtO2wdiXSIGyL/z8YizbjWBY7ksKgJE
Fjxa4vD6qaw43oNYROU+VSov8fuxDUXyANeGo+72akce90J80URdhoiZv7GbxQn/SngIqjP86PcP
Cqkbz6fI3W9jyc9ptyO29cA83B9cPBn/b6KPsU+Midfm4mIMRHbGIxX5nF8m+4ts8jNuedTa/O03
2Yg7GDGchyIaH8L5WRoJrnzlSEwUBFezKFhAfxS50xG1DhJlynXRRN79p19rI8s314TOOB32l1/I
gkC7RNB0x1Bujq+izIqvZRsJ29sWXuaUTM3sJzyu3Noubis/tkv3FL/2PL3/yhcWKIT3PoHHeLUx
7UycmIZ49AXDZI+IubaBqyXVybnKsS/rOaUU6Nz3iPVZgWcCRbriDvHJtnPhpoGHvh0+ztZ75jJv
Thp5HZGsFJaTm8csqC8ovHPaUXNS3oKO0tTXTgeUhkUeyK6CwdtDxE5rr++avzGLwhWX5BllcI8l
AWIALm6Mg9RGc9FivwjGYwd9IwVqA2Ma/OvM2oSTXu0MK+6XOzsCfSGyiA7acwd11cVIAyYUvA5P
HJ69HIW+6opbGGl5Y0D5/uphOZqLR0Z2UAuzrkIcH3457u9ubL2QVVDehmXEVF5Vf4iVpGw3TV8V
TGfavIgNApy/ERF7p7/vsZHbfR4YmweV8P2/mIJvo10yzPqcovAt92GiM6J4ahIxx767Cmt2x5jZ
Y5ySvsrqiow+LBJl0fTg/SYMlxnv9gQLY4TgpTyWxP/r4z5FueVHV2szlc0DPqVYysmkK8l7Nza8
Vk+MBPjeVvEWZRXSps2hkNcLPX9AKG3/DAYiFikkmG3HlJ3awK2/rCaRY5I03m7MEhT8WmNyBl52
vkMAnEkMLbUFdGor1MvOyVcLUKG7XfJt2RX1gSERBgfY2xuUX4D/pbxTl2eotabhxrzcUC0LhMkZ
/oxW6Y4tjZzTTj7xrOo6uddBOJ9x3gWpKNNVfXA0R3Ek52zu35XohlkHc/R4kxBGYEIw+XpqP8pj
Vy0ZINt7vy5k4gEZ7nonAw75iPHqY5md2QhCeGcdRthi1xvm0CNDLANQFIQ8dCAKHN4rSjYH7wZ3
eklWmgPwngdo1UMdGbX7nHQ8HAAjvoC5VpOKsbrtDD2Pi7NpGrTs1cmNaXgFCXON2uaoCRKEWw4i
HYRxpreWR14vTEJlsX24se8LVzsZg+k8Q1CHSRc1ZMKseyp/vQ4IoE9wwNa9rf+eJMTJHXy4sWEJ
57jA6LJ/zhP9bdam39YIatgfUvd4/IIAlmWPi1/rbiqIJuDxu+s5hKj3jY7M6vSg0EvqdHJBgsRw
LyKm3va1ab36hbTpXRYnRr4OAx08PFcRO2BWa22wXAK0XMw6MCHPqjuwie07P0qFvvrHCaqeRc8d
7GfmoEchPE3s5HJt4vhOGx+Py8iG4wfGmbOV4djyyKbgx7NoxlSMSXZkhGZMhM2Dd0/j5sOLCRtW
ZOQB6CA2j2UZAwUjTyiVdCOE/NEFuMbbBhSiXRnZ3ieZKsA509B+BaEE2NxCIUDRHtxL45gK532W
g3GZRfDaOvsspA1RHQLNOWjcEGP99e81mBlKN9gVroipLjanASNpsfBW4NRc/jQ8s3NQzwijunvb
8ffsW4xWlLcjm9CgMRD9pKxmTS2EiVWgEBjUSlOoLjS89pux2yHVXRc65+QzgcB+Cheqqir/voKs
hPJTbBNFiU4892lioozzYOS29bo0WiNJJKkZLsSct1JLCAFh3l3YdfI+TOY3FjCtWgTyK/TnSxO8
idUaFW1Z0k3VlFC4HlQLuECZ5RvEHwyYZEXn2m1H7hAixk70TYmMAvO2oqwdgBEF+TqwlgU/ZlAl
uDSfg9lBe70A4KMq0mO/kw5UVDJwkx1uSdfVPJWphDXoLz1yyhZHVxIJSKBpzO9udhpkHZl3lUbG
7Z2B8lVeXk07+3SI5e55dln+MkhPp+ogYyWGzPBHXO9LzeITi3GI9eBN+k5CShsa02Vk2EigDtTt
a6dM/tESGI85gcSIJPFj44xiOhZe+dLlv32LXHldA7BI9/wRyljmuZobfD+OUnnaRo4/84ctm6Y+
bhxg5tyEiy63jOCxRBcI1boql9RZr6ZDrt4WUqnD6JQJRUeGrVSgDZU8NaeSntipvMSlkfftDklr
/oJOZk91SmDzG+U5YpPAJFSoTSrPPGtkCYE6HnQSUautKtRrwLNMSffw9UkCCg/DDXVNFzLA/bgp
Od08QcJAanVVqvC0npT+AnmoMUhMUXZ6NOdU0UFUzu2DxAg4QZUdabowW99DeSd5JXmFgRIKyF2t
KXy/ERASMr1uq8c9TJK3CVIpo8yVbTYk5qxGMhJM2lGQ+TxfcrjjDyOI4hkOoHdtJjCbJ07PuL6d
9nRMAVtDMtHEdezAcx3y4mdPfMVEiTco335J9yVcYKeQXaR2m+4X/glofTUTV88XQy4SzUACvbLp
q+AdvWeUy9HwxMyxz4kT2xWg4/MYbong0mbFdBUj/+TKsKfnYgLxU61dhzPCO7242KzVEbjhcdvP
oJEkuP4/HCL9rFHo6Mrg6q7GRJQJrIax9qpKvIkAwM3qAJkwQHZXxh+1uprzihMJI0RErJbE4lFB
RMre29bnVHnap2l03ydi/srvck8D8vVAmYHPPAIBa5h1qno2fetHVv+OjxDrRifdAD2F4dUo30Zu
to8the3R3Bs75Wp5wY8FTDjeqZ7xPmuilp5eb9oUbzYYl3YZymnvUqmcyghsV9BFsDUgM6cZUddH
sZ5nSGqQVvOglfkiq/GDxhPpDrovL+a80TPfTr/Nk77OuBdNQ3UCjR0IAkC6Ag0RI/4VQONxw+RM
fiW75162DqTM5L1auaIN4vnpGxwpZLX4/8v12ozC1GbPs7MMvSpBVIvLiX3EOhvz9kG/f07ec2qg
h0kHO6kve7R1fi+0oplBpdP0ISmlbz4KWnn026R4oaVUjRNyUwRSbaNn2uHhxNRfGVofry/KDy6w
giljdfnfs7BetamFNIDTtg+W6tTGz3W4O+n+mvAS3Gj4uhKMOH4Y5om3xHUXOxHp+N5WG+eCGEYx
TDrhfttpzvwgbklmUYfs+qoxsRyjnN4gK3++fQstfPQDK6kG0BYLH6uDml51d/KiDUtUlECn5EQk
9TMyMohLz/k6CddOod3klKNFM/x1xpuMp5GGKvdQdP3rHLxWWjpKchraNH9vChKKkEtEEgpRyso7
woGYA6XRQg+yCrDk6fP9ohCMDh/kVVj9Eu5e+h9fcXmHex9yVbCS9YlyPWGIUGxtqyouNgZdPHpZ
cl8wrp5iJPB4/CC8s3nW4rWC1RiKE/kOtHoiZ3aHJg/WzXHEOuGqWOdu8JSKfxTbxnKybhR2p3FD
QJOZvWqZwwawQWEnLq/UVHuJx7T8mb8Z24hznHyVVMaxltEcNx5Wrjt453R2hxI/AwR381F+ONuI
h5zcwlg5/GuBO8adsR5XZyh9h53ZONUlo58ndARvyWPrSanzK+WPaAEo8K/iJAzU6+VHZrjnrrJ2
Twtt5bGWigRE+a2zeaukTBIdq8sPDo2ORQOaKu7o6tcodzOAnPGa4vLv+44b3r1sg/ClR+cU0hn1
I4JVi/ZOK2D/5Tzdh7IRVKnTH69DNFR6D3LSyGzXUrTP7y14r/IS5AUMHWILkqwPJw5K7BOO1v8v
R/q0rwh/hbtdchcMVXvusAwaW4443EkvfNs+4jDvljAG7moRJ4w1RyU4176+N9qsFlmEDTiln8lr
nGVQac9osWcLaA2MWKSWc6eUOGV3WWexAQs/bhaYPxjw9KleFIX+wBgdgXfy6VndahtMNxy9ZwCc
m04PQA6x8O+DEZ058Hv6eRUAZRFZT47XAlRhmxnvb+V4NLiTvOrTY2r2xzpRHfbcPCovZNV4yngv
YKzpxhQ35nEfAa+gbEYz2P0xXlvxWaq2fXJwviajv3UiiOYXkGCv9xfTJbazC0OYewNpN+IlvWg9
IFlrmStydOx+WJa3onXVcFaEQck4tVk0wODkGl0CeSX0US1Qf5v1O4RPuL2I9JFrqLBe6QintXfu
cnhm117ig7P2LcqkxckhRIyCoi56Yj+iD6qDtZDq8TtT2NEBd9ilS1dw42IattqiH2kpCpfbPjxt
+H2tv2W/wojGEPUKxkCEVAOAmhqFfb1Z8kuM1wPXsA/aWNCzjH/3wdFwSpiP9vThkM0F+G1dVJ17
HzVemwab2vjcQfvm+MFALiCFdBX1olVmntVf3OXeayda1SpzwP3MEqIuQ+s0YHuVV2OWVTjGWVm9
Sdi0EEpFsGic0h0LJYIzOLbxUVS6n73aaguSKRQVlO4ORRjLuDKnukYCwZExUflReqHxsAJSrRjE
817QD5XtUkIgJ2UGibq24cDQFQOjuPGb9fJHzWKLN9Qmzn/J3Js/ROerItoqvUDrEt3ngeBNjHW7
Rz6HQu4j0iYEUfvsh1ls1S+B/TfhgjA5BowO7ccUC5kf0WxawV8jghYOcfHfnMz+ud8eKQE91SJH
DJ3772pgV/JzE14r5K6CA8E9E6+dZDFEY4xxageswyEc24llU9vTikZmATULsOLVRGLJRa6Xd1Xy
0RvLZMsDDxfW86hBj92W9iTr3+Tnr4VoI+vyVqhxu0rgNblCRTl/s5BCw4xgpOrm9G+z4GmVhCow
Dw1e8BLlB3x7y7wf1KT4cUZLp3wlWXfe9UdAEobC/TtclWBCRZJWUL1b0L7VZNDxteudcqXLuzR3
N1vOyIaCC9IDCIhDKFh6TXGB956ki4X0LykgYj6gmTAZit6U3b3f3VRh+Ry4OEux0jrTSH317X7F
XCUx7pHDjpDBEZwHkLY6sbcwjKfXmiIIv5Wwcw7tVwceRl+gZoNjCnDHbewMRa2aLASOC+QB0NUy
Vc4w9yHFHH/HFVh42bso5OQvAgQCYFUbPAUpugabT26xy5VDbT0ezHfgE8oM+nSeDEKyS+yKSH1z
THcZ2HmKdY3kIINH21fUlT59ZjY6rC/uNmlL21TzptQNKEGhfxIBe2yXqc8Aoq1XoqGR+f+dCFa2
byWXuSgH8Uc89sLl3m+1X9UVglrJb8WvnyIo9Pd+DD30dDw8Ai33Om4ZtTbngrG84ldkowEnZ62t
RGQ31y8W1YUbPdeY/i6QQpYlOlB5b6RaTZA7PX/sjB5bkwsi8B4UPnLunW74xDG+5KyvYT95U9Pt
Mrs8hnWZWkPM4y6Qc3/wnO6vSCW0f41uKYmXcecdD9U2gpR9qibAURmEC4mzhTddfzMdUpSSmlPc
pRQnoYv1UsbetGvJUmwYKx1zAXOy/M2Zyh3itSnjjjVmmJlPfmZTa3EieFCG4BeVf23dsuCV2Si/
EyewI1ubYcAjhdYHIsypwZX+hJvsTNPSwSPB/RYy+PrxPKNf/2if/xCDcmVFgzi36KGczQfgDnc4
YzYlWhI7Md2AZhSVLcudOAPBsO1v9YHlMM9cGIaWb5NmDkfUEfPV12V4KzR3d8sU4ljiILhW0ktI
DQD6szsW2FiL8jIV1y+xy/r8TAUIVxebRa8eVcGJz+IDc5d8jv3yR8H9Drxq2r2/5ccC2kA9jNk5
w9L4RvFKVlq/RBBi15lD66bXuwxVoq4iwYf9sj+FEhsn/gg7qa2FDzbVCoI0B0uvzOHhYAisGL+Z
08E5x6oYalltk8exfoRxJxUdAZS6VdUTzu1Lyj5cs4S05WBd4qNGOM5Pi5++1iy9b63H6nI0QP87
hNcR13X1MMwZHtCezAovioxRVJgVSx+CnAH7iJs804/zySsoWIWFWW0g/KPk2WbVR25brwz9q6qu
ch0svSJlGzBxWMcTn1GrJe25jqKHI/jVj/KzxxOPFMr2S277wS020AFGeQyn/mhNxg7uDYwljMMY
IvgtxCTDoXBCLExsW1aifodEDbIhwB/KD609gTGsB0dB/E1hAVYxEnitVK40hUpUVVJkZKFxNfXt
QKYD63V59A9mt9g+XlMIf9/oMzCteqWWN2Pd1AUJgFW6PPNurYVDNGCXCFTayZJz+5aQmPmW0KL9
amJG+xxY9aqod9TWd8e71knNaWygwsfV6UFgbtmvZx/8/B+o+X2b19CvoqgG/JObAHz3DL5htLjo
6rLkq+aCKmCH4a7lWZ5t1/9ZEmNkqFmReHgbb/2QycbWmqpBkU7FojyF62XAgsRI5NV4cfSxrkBZ
/BnZfpJxP3adxGJMLR0OPcdrZPl5yweelg6+9+rLr38Fp8Nhe1J/wNaTw7otLsoULL/4CGnjF3mQ
NM0wMDzZ9wEGLN61KASQ8qhmtd2Pob6vlOKeyhCChBeeCuy8ExhHxh+X58Kyv3rsek7y/l0RlTTN
Ag9PDfDPUTqFjVV2orMR7P56gwFuQXG0R7lHFYuPeMOGu30vXscgrCTTT8LoMrrGHqTkBNxyOekA
P3U9fA3xVknA6lNPItArEBtmfOHtRvGpAAoUqCWqfcCNC+iIrd8fNp+EJN3s/hk+j9YjAh4++Znm
/yjSNXDZLh9SIcpBTvZeINRo4E46/jjZyKUXRI7vCyQztmW03ZlaHydueg25TaDbU7azDikOtny7
BPuooGL34E9Q6qv/X6cW+Jl9032enkVOSuvKodBppNoShSrw00mbuoF++9Wpq6SAGilETCnFtam7
sS+hwH4wKCHLxDxH55vITIoNpr9qvRrFd97hCh9mzK+eyIZzwO8UlR4Z0fBRP70X46HqSa9CpjBv
PUpWVQ9zgJdHiaWlcAmOGqfcNebg3s9vtbsSVojyvNBfL0ponE6N4FYDMdSbH00g76ks4vtKg2Zr
ukW6uJ2yntwhJ50DLjM+V3b2C6Y6nIZhMIT7HDp1HExhMuR83UjXxYvwthYb5V8pGqoDRomjvIRQ
Rjm1F64QKUc+SPJdTj1XMS26Lnfub9cm2Rx4ZckfQymPzs3GlQLPIMFQg8HkD0HSO/+JZkY545yR
+ho0sWlENkb+uBqvY7fcznq2KHtewRv7pu0UzHdMpaS6zuC8bLsg3+gukC4Gy4wFfYsrAHVtW9di
xAjxTXl7h4403/qRd4KsFwERjQWiOasN4SdXygAQM1UWpVVE9WUPuGNjgBOk/no4I4OkdTapcWyF
rJM5BSwvTxcf5BtS/uAvzV6uvLdffVTV0XXlJjEDinvJETaZCg80bUtFg3fpqc9YwqmsSweLfMfZ
jcwEPUFgEUyTADGQ9giQYg1YXYQJ5M8zIDW7VOBiiinH0j9y4yCnW2r705RgTbYw9msZ4Idk407f
dG4yLH+C5cUyF384+SC28vDJc35ZLZllVOjszuqiWx/XP7RNZT2jjxX4sltH0LGhwTsceSOpGKu/
g/R1iqYchsVO68nHhPTP1e/TRA4SXIwc9G55MuHQy5vg0rdQislbYoB3mKb8PmUl74C59/anLqjm
34lpbueOWkHNeQIfqz7de0mVwas29O0EGoV/DKN1bExv+Q5XKKB1Qo+wpWuUYlbsxgRMa3WYIFEK
XLlbA/0+nEE5xPWGSzqZvkdtcyHCcZtEdbD8hqKIG7yNqmitPUPL8dzvZCKhf7CuLdvPLre4OQe5
MXYzbeOU2w3hAEy1abGzXHz3fXeXZdxNCriXgJzlHXEwkUgMa4jj6DB9SXXgnMFohLWJrrx2BqsL
aN6vZzzNugEie3nhGxbpvGoy5P4hSgOSovFWNyd09+GPxUSm9DZRubUQ0OX5Le3iicA2GpULIeXn
0aBJsha+SemCMm6U5kVbocgUclMBdHBMQZI9+vnjaxK+8c/MnWV/eBizEUs2+IQ5AYHGRYjPqZg8
vMux56LSnwiMYG7QzFanZBER484dDSLoOkS8DkABI2OCWViNQE+m+jrmNQxtYXabtNj/Jwj/H8N6
G7VMtpDLDiKcaLyLpboOxSk/iOpnukEObF+SEkWsMkpYRl87E9vUkpUrwPGw3wZJlE6cG4y88teB
1H7txa6RIjNJ8JmESgyf4W3pdfreUe2woKm0DuEr8wZ1Yh8+T4GMZ1bl5pvYobSvpjiaY1KVJsdL
XMS4Ag7U+5dWhA7wG34bKqxOmljPSh9pQFz6UX+KcpocSv38N6pfQXhaQ8LJwiOAOgJtTmAP3cRi
XZcA26cWLyKD16KlNpeiz0cxT0VWVlpvgfklscdouOb6+p0hnhxYDiAp6/uD/PSSwf+CZ9Lepayz
P2C7C49x7iKVbYWom/BKh7zq8coDPUqaBPZtAhp4CO8H345dRMaTLQPjsl8ayh19iSP9l8V8rU6b
7GZ/5XACxgiZ5pb7/LdR5rWlp26wKST4rA7u9ERF8mG14LRiq1nBlDgmxqW6QgefftZAZB7/yN9R
04yRemZWh+sAwq69iFq9eWS4Lu95pICgq0NDZJNkM4Z9vuzfWltn525rFzhlR/9OlwN5jyErMLUf
dpfMbLR3Quw9wN0nkiD16NmT98j4fE/CZyhrLpABzufz91SdoExqi5XS92coT471KD2whIRohKTA
uROHCxWlH4n9B2enftmxOIph730Qq2//yXREM5jp4/73CTV/7LQLguX8qD6gprkU9r1R1rqoRG1S
XFIc5Zua0rHUOG4TFMrzqpi9RIlw+IDYUW+LTP5wv0SUEvZLfyRbfTtRKj6g9NTC5ymJUMgYzip0
HNNnUqJMqtLuZzbKr+oy/zrAps+MZd5RHvybxXRNSTIvXFNaMJ8dKBzqk8FiMT7QR5Z1xvowTJoo
STZUPUC7Wp20eI2jwDyh8/kMDNBiUReaW09e6don+ZxdXNIgCAA8FH8i8X9zO0H0zT91pEoSkVqS
21ougGTVy1mRRb5NYUMYLHerzJ2MHlVlUXVNuM6xUtFCJCykLxy2PUKMp9KMETycT+U+CJ8Zlwsb
ZpqtOu34cklO9ZV/N7EawQwLSh6q4cotPIZNzamYCPsvy+bo4vI60Xby4xw+tlzyIyD5AZq4j7Q4
WP1l6zs0AfGXUZ/Fs6MfljCXtSbQBDEGmeApEBwq3R/aaHHBJ7hLrDJMwQZPIHVvSxcOtPuNhErf
ZpE1PE3seM2CFMurPzev3aPgbZ6rhzoW3o+gteMoJSvedh/goVMEJita8D8hiDH7B8QcY1uMC02M
JBIN5zWkeFaV9LrVL22cTHk40hw6bPvrodkFcO85FrZEYQ9RuZY3oZOrH0QIvmUwWvAcknmNTPUN
WCjtm0y8iDtdGAsOQi/JBrBo8ZHcpPczYUDYuQ/jwpQOOET8vSf6VuQjD9Brc+AsGwdjdpQ63BzR
+MTKnttgPgY5mpUJ/IKSQaXG8XiSvNfgXT3wt9ZWrHRZBpkyE05C5cQSGsGa39NGa3y2xcKoCISp
Ul+F44c21bqh5V6EU/xMr6PaaZTBIto+7Cdpf4t7h2aCm68fVH4VIIJxsqw3Eq55qzE9YU0e7ajR
qTpVXbljagbVrkLXCsjki3addc4MQHBAuudvhRFAcTR9vFK/LZQlHf/RU6lxyR8/hIRyTHKsOKR0
nmUcXslt28AHpFF7H+3A61sUeRLyLmWHKirJYtRzM6n8Ljwbky5JM10srHq9nPo8KGm5Ms8j+Cwo
JoudHfhfFL+XF6MAn/MaSfyY0U2qsDqCPu2zNshaX7d+KHOxnlPkerIrd/q0eVmaYz7QIpZTTxB7
+sF/2GMNKVYnOskDf6sUkTOfcakPwo3xlpZlhtnwQgWoc8qgGoqsaLGVJtcN03X1Zt6CzlWViYZ3
BT0X7tXdQyM3IQIo9frHqgOGd+ZKwdGEXIakRncFwlbkWMwf+OYdJkHWLK2YRAgk9Kl4dciwymQ5
DacvdvFHu7+DyTXUeTHUOxza0LqrD5AKco/SGV65cHu5jcmxJV6HZGBZ2YzAh7WEOroQxhGaRjdH
S9sghrA1e04rDRmMdlE09rxDa4Z8JhJEsfOnUy7NvhA+C5uWrAaZEItlhKoWGiPRbEXLWrve6AEx
vP0L3X31gAXqZMgBCACsmbmbu8VAl0A1RVNxRsGuDZzCOjDmuMXt8dB0jSmmk0HicVBj/bs5Upfe
xBI6MHbQKHXGDP8uYlG8DDcqAHr2DHL4OT8sp7OSQ4n+f1W9MHAssmIgoRHzL1FFGOr8FdOfJLFr
obUuc1Gefpz4rhZVDyvBFV8gHvmZ+tJRkga0lBzc9G9xaWBctFwwZ2gRoGT0jgoNTDzujnxFowWc
ipHhx//S+pxCLEY7p3yHonjUfG/V+Sk3203cbjX4s2L7/SyE4brX0zr0hF+0GG0vtP6Fji3bPd0D
ZaGv9o/PwyrwYa2mMkNWbwxRmF4hPmbLWLzJ5CjB2OpdZO2quuCpYgWmftQNRh6FwXT6kO6kZ1tk
JiJjdLcTI5dPXEhUrNN1ByPAd5jmi/3NOIiUNIzkTBLtwtgc84Zrt3uBP79VJIBQWfnzC0HjKBtK
dR4zikplmjFUcLkJe3VRcn0zr1SpdpbO8UFHLbI6RlSstfClcTiUsxwy2RhvREp5mjafaHpUJaxq
AnJqip3Q42NstWXLxLq3iGO1CKbNTzXC1AuDvs57PDLCqRKnxJSvQj3zAq1zGMFb4dL4xTofWRa3
zcnFjI16gU/rmCbChzOt1nhiaT4M916vxipI1fQd/yMdMtFD5KQpkt0LIoigpm6F70F8d6HcIob8
7clOc3O1CvD1u7nYNv4cuSXkVyiaHXSNQZgvgrAUwGp5THBv1nva660ksxS/T/+xEYGCH18cj2Es
wKuM1jtkz3NMFv01D4VQiXaGIyu2sT6sna8aLQNm3HFs+p4XFRNlr2WC6J0mLpO9e31jAmv4OYFv
DMagc8xAOYrCqQYreEidk7zaPrtU4FX7b43aOYXdHlxszzFPAF0KxppV3eyG5dypYsaSYGqCrQ8q
dl2cECi6dMd++HmBADaFuY8PIhgs95GJWqD2p+3aVsh2/Eesh0A43FPUbyTbMz+N6PwuJ1SHcv3g
AYJUfiP7itqMzvbnL0ydj+4I/lYgg0nsiOwCJhQ+TU3VDJgSWOD7yPaic7fdj4DMrI7qOwhh/fAY
r6L6dLTYvHS1gwtka1F9kxyo9dyRDze3CQfnlarnGS9+pwDifHSf/38jTYUPDFgqHY3KtRoycfv4
l3TJ5BG1xLnA+nZzYVrF/yinPUDr06iizuLAvqA3K6YjJ3iuKjVlGGI+jn8fX5naQ+IV/izNswWI
DEdvazRC7WRguvtlxfeRwEDUP3k+YZ2ei9Lc6NoEnQz2E7Jll7E3+Rj7wKQAY6HKRo+1j97lvxg8
Z7rAe+36h8A2w1tOM2WjozNx+rVXY1yf7UeH03n+Ur7cchb7j8M8r22SKHDwh5VBRcJ7uoVHVflj
hlTSa8p7+cDPoiNw1AtNyNV82Dc5Ho0jevTnlQqgm2qoyLv3hwsZvRr4ZKeA0ojTJ+VZBGsZCXaC
QUcPGHhxMN+X/nspgFSieO5+Pe5bzPPqmTdmVL28AB4y9eEsulzfr8Dq+sktt2B/k9CIzT7IPtZh
j7EUN0bulk2mKxn1cckFx/LPQFJCfAiDr8iEwfWpxXi5iQPM8gT8rw2UfSmJSSEbvZZq+PJYOmHq
7KqIJj63Ud3aeqWMlVPT0nTvHicWKLFjcdEXGmuzEOP1gBb0rC49OUK6BgqT6c6DkabOXGe+myoZ
Rooc1uKfOQUJ8uYZD+s0Jr7hIIaLG3Sdc5nHkVEXR3gEjFYk/f7yRr7cPobDprYfno9qZzARfxkt
D4qdAxGBLkRhC9DrPL44Vdspkc2kJclD+Es/Ve9auVjdWBScBWhyMZSMKWjAStOIER2Y1YXpj7xG
oInyjqzy926qxIMD2zgbTeiciOcFwz0ZXIkxTUUHtEbTFPOkh/WbtJUxw9ACQsdY+8fc2iwLolhS
0p3xPBNhDTdRv5kY+3cSOfVARK1vYvPJSidzCjPgi2hiXoLLDquhi4cl1lPIJyBqlyCKawirx6M0
op82u2wJUfsP0TmmX5YdGXGJSbz3Eq0M8Kz33p/ukVe7Sot1QDUWt+IMEmsc7qHPAbMm3CzlO0XE
bYsVwD3C0/nJsnYuhfZkk2+4ZEOHb5QZKU6xUou+4M1YtTOOSlXwpVH+mO2JjWsBR8N6NfHtYpun
K+escMvjqELG0fQBf4RoGk0vAaH+P846aXHbC8l2IoDAOGruv23JJbAfPbD92OSMIIUw5LFGK6t7
hEXsurQZZOXwYd9b2XG2T7qEgYpCgpGUD/PXO12HFtNjHW2XW55nJ2lgkNO/prgMtpf7pphEwuEK
1LZcByYmPlNO8FtG1xfheeGAycKuTH56QMJZvSJPLiEhDmb/kQvDbsJ4/AdjX33MEp3IhXwDHSAV
5k2ergL5GAQXcSw4zuyyEUTlmiQTQCllf8Lu1rPA4xBJXcw+XcBvF7VxhvQRhWQB19Dp11X56FfV
Ju5pAs+DxbeweA5VpnFuu58LRbJWAU9hRckY3tDbVDq8/e6hhBTU+NZGJK5vRKnggEDVojG2c7ZT
WPmlqnRF8KNjaRfhMJjWwtq0DF6EivPZ+IFiuj9VSO9+d6lUneRGwQaA6TB0MmIY+7unGvK/gbAf
ezA1b8xvC2LrLIBwUb8D7DZK9XAeVxkXU8gZHdy98OvC0oAyIxacTomhAB/QWyzBMzbqEg26xWN0
j0Ay5gm16a+lejupC5Wg5/ipEEybLcbrqKIMu8PkrSBTpfGH/xJfbvB4c3Ttffcz2TWVodKfH1Rg
ngu5jgMWYEFtCpSIEzEXgOjEyc+v5+ZmuM6Q+hWBiNBE23sCPckHqwi0/OjLUO7AXjSNv7YLSB76
cGDr/BebXmoYTjwCJvvuuk7JIPolJThYN/mab2sis0uJAk0Qy6tC7SzjCW/Uuz4l82vlFOWIB9HK
s78Xe8DiaBNqmLVmd5fyQXgJgr3kx04BuPgYup1AjlitElZcnqbvztrkdZ9ldtU3LpN1zs0Tq4xB
GDehxCN95HCR6M8vP8LwIgny9VkZl3NQuTbOTpqWku2oNwDQQ6B/tvcHwfe+1qZ9ffs+MVB/54n1
F2F7LcX/KssGxr0Hur+Kj3cQyq1Ad0uTX1FWde3/jqRfiLh1IsPI6SvXMfQ/KLG5PbI72Ixi+aid
ZSY22i4Gw7Xc78AjaZmiLhYRUf5qrykszNM0OjeppEdUFm5XviZvfcMWU909H1apRL5xvCYbRaf+
vhfNPKYzIqpT/BmJZ01Gts81wCUXw8iZVzM66nb6cZ+Hvj1BPE63Jh3bzXo0z9x9+JQCismBGSi8
V0EblHcmJA7i+82Zg9EjSHqj6Epod6k1gbFG8X3vSr2f0eEb9YNM2R7nsqKf4iOe4CnxmitVcH0K
kkiEaM1cxYrkJNlm8IIfZEsS5cuEIYLRlbeaeezvEZHQJ38yIQyQ3qTmf/H8E0y1b8QwAnfThKGx
8ZT+F4nyxQ02n+WXlG3Xh2rBdEP2I2+Nsg9oiM1LW3gDGUYvFHVkRWBqxDUMdxeA899yi80u2hya
UrWZolkKa4ED3sF27aQhefYQsxqi6VZkeVDbJ9POI+qI/dWg8xCNOQF7NHsj3l5Fzh7OWczK4AQJ
hEERps0DwnzXJvRwwUyl7iKkrmmpdc0xA0U8N/xRPK3XmtG3urDW3U7cg+EkRcAAJs81LwoMRG7A
gTxATnLW3nATeFs/rT2TWPS5ZHxIf4QECrxhs6rIO+QzrvAVV0kW2SskDbodKxnGXFur5564UzsC
SGMHsoWxFJYOHk1A/UKypOQU89YaUED3Vm1FJX9o81obqMJ2mQ2fZFFaaJ5ZIBKK842FHQ1N6YaT
AuZ3uiOC7bR0kF2vGjIVVPnfwRKZQPDJFeEHGbePxKTy/R5h1rDonwzfBbrUmWWH6Ioop7xO9MZa
Bvl2wNN7uP75r2OlPolfjBjVxzFDI2lwZX+/7Xdo8TnjLk+l5xVf22BwcHUJcEGsDViXm/Xt34Qh
LEBMZvMEBXtVqqeD3JpuSlZC8B1yhtAQXAPJ6d0WgaZym3GfuvAIQwsTy4+aWE7tdFahhu2+4exQ
vrEqsQudti81wJUDYQi5nnok7GnpK9j4ZyxdBOfZ7O13AzyC2i+lqcGjcZo4ogg8MCmEwvMdF4+V
MMHlBcnNLpIr+h+gjJxSgbjqfgBTZbWp6PsQ+wMaawFYS74qtO+wejZEC9450+YsTmbXnQEg4aAU
wkZ0jW2ipeOnaQ+JLC9/bB4FQIo85arjQQOD7fmz0aXwOuYin1EzMvPZLaL4MN3iuMgWTlUP+3v/
WAgCRGgdMHCkuoJmYTnb702B4gQYi/2vluLn6FN8fAnYNw+OJ7bJ8xOhSRvo6MUiAjqWL2SL1z/p
ueiny1W30k+3krUat42Uowte8mRuCswxtDicXL5L/0aprMs4BGAmSRZ6C0PQM8LZg72zKeJLExia
J+ccffLxVzZCHDog1WJYeFYHcB84Y7JT+VJnmYv9cE6dU/pukLH6/L4+4aHSTXHf7ThrReUyVSjk
r7s/UrQTbjf8pmObXy2FB4SF5ffSCrZdsE+c3/fpgjdCjeKMARPRMvF5jYOdZImZsYuRfu+jw2PM
6P+ms/aNUUJH82PRn69RovUc525ZzYgKCOUvl+uGB4CrraNTRC7le8QGtXAyQlXO0JYDkev45pUb
OoNrpIcxTqHR+GEUUCe8f75ZKTnDvLdLkDIuLsx71HIVXkwT8+g2chXlx4ewfVnQhnoG53uNhEiN
5WFFpKweo9xlQOU4nR8yhvm2hxtv5isP2DICaa/FfULk/Rdd+hHa+uxPkyhU4lAKXxRrrzMfIgm5
CGYjumc3Urip+bklMn9QIlFTeHU7UABh7G8/yWV7dV3I58vJd8EK7YRPSEQVjWnLO/7+26ZlxdiY
zyINbSMp1iQi4mOVqP79x5atOndj2gKBa6tLidX6oL668v+0X+01WpOf7DdbQcfO8HRk8R2gDTdp
RxzJHSYlC0UuLD2tZuI6Zto6TcDe0DQpoO4o5UT+xV0Xqa6OM88xLICvfYRxG5b5CGy+AnZDGlrq
qJaWl9EA+IAeQQ5Av8pStja0Sg3wfC1fxn7GaU+c0SlyTUZ8y14nClioY8ICtc/uGiQ+dZRdEC2f
J51HstvQgm6jvs8K/6HlclX8GLL09E974DwoXpvWy9iAby4qjqEGStoqOkyQ7VoDGoRgRU1bXvSa
UiQGUOi1y9ZtZfYdvZakRuH4RThDfwkO23RDFwcojD/YMYkspoiy1dcCmdctMNZTVj5Rv5h62CU4
zlsuwE6MKdeGPVnc3GIWaIo/Bt1GupK/ppVej2Nr+7qmJeLz0V+o6OX0WQxn2/t41wtJna7C5RdP
rdOSO4mTuKUbjaPoCllBJuvZTLZ0vFfsXE5j+3urQ51gfTs3stg522oRn19X0bYRlHImU+nhJcPO
hFw/MZu44XDk0XQ5ylK8JQtwNAosHhXWearNgaiekUlxsCdgKFSYCPnd9bIfKjQzj5eFQnaVGQeY
l+FLZrVSDUZ5Xv0U+bx4q4kHkPdVOCK3W6JKsAvMSefZd+jh5MN1qMz0SfKU6iNdFTGtCU5caCWX
TKKtOmgNGm4Bce4A9B/E87Idgj9Bqbv8jMI1GeVpSRh3ZUXB5BF2Ps3bWSoCt4hUOHLvE0uox4mI
OW5d7nPSEP90j9db4Q7eDg7jMC2c3lu0ZZgfjT4Vsu3JkL14e5p8wcdr4OPckGqnibzq27ND3usj
ZGxBABUdOQPALaboMaUkYsuLeerpB7uLN6ao+dQ5dX9Go1fw5y8cu7k2QOnBUAZ77fA9trqHlQyV
c9GqbmBwvaDeijsQh55xytGewHnF6QVYm7ZuaiOsC/ozHaBn4d0P10cQPjXrO9xu054Zq1PJo9yw
KkiEwmw298VOxcjvEZsrkA4LqnYKbobn4jVG4U4YL1HD/hb2u7C3GLrFQ4si/inzUQZZ9EZ7U06B
KInOALheH1BqRhrnu34R7I2RDTncVDxBISQcitH2gqrkNh8BXxKJ4qIzj7pTsFgvdPDcRUsmNV72
cmZjcDIyAOKTR6FEw0qe2spbjNMLr/ConsQsrfO+vTmWxfA6unnT1i8YAcDHWu1MUV+r4KEiVTsY
2j1VLif6tMnE0rea5aL/D9QZhELm0tQ48/+RS/p7uW71nmzUoxGS6URI7ZleSqVv4fiT5SWlfspq
qhWJihPUnie45gAf5TYcavHR75rCxS96OY3iXYIrnYGdqdj3fyy409hsV5LZPG5Z1kyBC2pMn1ip
NPLyeD970YqKPOF3mmGc/86w4h350YvYSqAmCJjOooZZcYpI8jEThCyAUmdXbDvf1lgnl8P/mMEV
AKy8zYuEQ0gnea/NIjTmMDPPNSrzYwVf2lcBZKHNcRT+wGVYSh8CR9LJg+HMNPMUXU0YmkHShyez
1YiD/vPrEYxuIHq3exnuf042DiDWC2J1yENAZNjIq0EMApR6UWTxeJ0a60JwLwdk13GX9PwFUGGS
ZEVuhKEJ2YWiVkXcZ50gZwdzuTa+bFnmWcXdzn7QCaG60Lqa53sJQobNYNekerxbBOAlNVqd6RsJ
ZzVhG94wzCtUfRMZUb23EFEyNq9wRfCa/sPinBlj3j5kFCfM15bCZeLIVDdTdy1jsIKD6LU+i8ru
sH9ZMlxR2I2H6KMNkQ/KN0Pxo9Dn6kY0t0Jxws4hQpwYduu6pPhzBHxCdmBw4r2PqWuU4sm9AggP
PWkTImMpujFLFgyMjNlOgZ7hhYcUhJMKovLEGBydEMRNKv87nxsV5qDvVvxkntDccStWgQ+skI9r
9/EeSsE1VcagrRQmUF8oiQ9rsaWf6kpFISAXCAYdXrhK4/i+rTWELJ02oFRPQBSmbdni318OUy7A
kIveuwLTDNNpnIhchMV1W8zPqMGU/8nCfOsSyZv0ls8rZx6Ho8Y630AOt32ND4s51r1XE8JRAz93
nmG9vh9xM0ESgAziEQaBoN5IHMbfB/21/Od7mld2S4RP8pWztoLv8GBq44Pcek6oAbAE3FLwwnYq
qexawT8j2IxD7DA4x+HVoVFGq8UUWPVPFGHJrxMc2+1azUNipiz/+nYQ407j52xVxK7QgWfsZFjT
y4quee/huCEnEKSjxPvHcHbDsZb0FRwIGMDXMT4amE/sZfxdir33K68bSMVHbqvbdxE/k5E4Fmi2
lmGh/H4eq4M5xOwZB7zN0gQ9iCkEpVhy1Ou5Dug5yORbvarz+FbX85JdaFcWAcJr2ZFtTwThMIxr
jHrq0ZjbAVSXTtlSyt9V84YE0ZYYlNNL4O29NAOJwGqa4gjFo6KMnn/W4XZiQB61zqiaTvxozN+E
jyFaStHo0QUuRYQXvGXJC/bSNuWBBBmvBb7Bb9i1iVsPZ8GZpghErjzLN7jOqWJ513Y/sGaYwTYK
Vlf1UA3lOxN8NyGl9tgWdJp8+UW9qB6B5BU8XT2h6X6xqu47kubmc1c97qqjewYrYNtpYw9BTU0x
YvQaQxz/fni1F7ZAE/zxSheWMa2InYMXtWM31qejF4zDCIJPv4+uw1gK1Vx0SzZDSps3Gvq3S1z8
bLvgZnGoha2k5L8oFSYqEO2RtteTqPDupiz0WfLeYMdpYSlLlfCXuqBJnT1rs0mqtGu1yM1NZWeI
CoCr9YII80NmFnqA0iWG3CinNk0SxqCOdRc5Ux+s4XgyJvAioNztVZvcmCC6Oa3f42q48om3DCSw
ZQ2dslFn19tZuSPOL8eZ7vRIQ1NVFF9mNdhccv20VtQF/tVwb2cPGBGy3LrwGfbWyn/mIAw2IVWo
Dxx78qmrd61ppg8Kan4zaBuWLMb32L+lvFvN1aX+hNyP34XpM/DUzDXd+9qWCsklz2FngsjzrD/W
BoQHoXrxWf8UmEjTZxAlP5TJFkDfuZWbwEoSPBj0xJaSLoD3u7qhEscdDdnfYZn3p8ce2y994Iai
t+uXCvU7/40a+z5XiygqoLCZ33tnATe9XATm1NtxLjQM+YNFBZ8mJV0AlsuNSddm9K2rOESM6MF6
roz26S7DFizC3ADnB594CJQESgVt12iPp17QFlZBLbg9Aw2Kw+9IrZn6Rw7mGqzLKJxMTODY3zBT
KR6/L69Wk/jOE55ErRnbjEM3SxAlJ55mAFm6rfrJT2tc7cu/U7H221Z2O0L+wxfapab76MWTKqsH
MoD6ufRsHofYffQ70kh0bJXb5CmtImIBILDmsEFOkmu/+3b+LHlCfhXOEGyGjvWfFvZkfx5Eqw1c
40v5Yd5/xWWBijgDCVvN7RHkD1qpwDOUPfHUPj24uodzPQ8rZhMnI0kllHVGI7gDH+oopxqaruI0
DObJ1TFjYmG6Wi4sPJ3pdGAJhpl/E6XWASe624gJn1oBh+yLFtLoWxUG+Mxi4cXHPEFB507P4Hb0
1CT/HJGlqPyGQpoCBNpWF0UfU4n+oVz9VyvZpFWxQfJfyiIQJVAcmGe1ob+AX+V2aqjPvVJIJL8a
YkFi9JbwgceVYS2x+satl8+7shkkrFEDlWjXIScDIAOF52JtnVDMJ7cbPRRERw+ZLLzNQzTeZItL
PCDDd6Wk2d4ddDQys780auKW8VJU/fu2tMtoDnccQHpLKjooset/rq1UQmekIADGfYGj9clHHoti
u7SWFpF75qL7XeVuNLG8d3+JX4dS2N/4+5S8zY4PBwj+avAOJqpWnJn/G3tiX5A61RveksVo+udu
sPW37lTBWumQktbOT+/eje50O0hB4rABIferhVZIR1pXn/7Yn2UUj+aAtSoW/KdqRUlVYZCogeRT
r7yivS0w1m0VZZnIEfVOS4NlHzV+FeGtyyhklYmLMupra3RmEqlWAanlrYzSEOTV21HBBNGXUa57
dOsid6vXFbgOQFKiyNBUsPKScg80RqU35YmL3eud4/n+hT7p8VnbUi5k2KLvV3Aq+odXXa1OQS4V
6MlS6O5kF8WXZ0dpUyxwXWtWd5rb/94XYGPcOt1b8f7do6M1U1Qdm5uYxgcSLNFPE3bPPNfgdGe0
3kmuFRwWl3SYFKUj4MIfDaU6KEqbmduBSxYI9xFx6Q6fkfPcw2bkdnqpS5n4xkDIJ26uyY3GFoxD
UjA9s/tUkLu7iUKqMaw0IgSXu9idNQweyeNmRUQPhmeHKBfRg8AEUd5+N/8JeYjhyOQUwZjVahXq
iqYoKt3OTP0P3phKBJbekIOM5beAj+u1pl2t4tAXvHlQmsW5edBPrv/nwXynnU7tg0HtSoDeNBVl
2cytx1KGvKx/YdrILb8XhO0oHypXpYQ2iNbWkrsuSfChy4YFX38/3TQsCLh0/EuRg0uXCCiBjT/7
ZZjEZw9UqX9yD1O4+4fVaep0Hzd4gkCrwnWEditmTQO82IZ+CP0yfRHsB9ahgZCyubraiKC1LNFz
bACH+eHluFA56pZJvT+GwDuPrn5eSd5nwAw9UV3UJQVWJBBoohKQTTvyDbQhnqbOU0zzYM0UjtHV
IMzxXzDG6E25ic6/BnEOKxOlgLsOAaqhPxjMqMmxKrpFNALqcotV99H/PpSxD51mN8QMzh+iPyXL
47AGcHULzfd59SRFAgFbCGoFnEP/XP1qReSJ1qBtlapxn1oWl1c/aEAtpEumxnNyRybDdkbhYNhM
4X5sjwSpvE4wdEJXMbkg1+cbkpmKnIrK394S13f25XFPrMOKnoK8nJwWTpCkowgP1bZgWQwmK2pB
z4qhJ5lFOwHaUS3zHWLnJ+F2KSn++G0gnU5oboq22HHL4xkSXPFgrKpEPyd0xYWO5TZZUEfoToN9
SMMTxqIqPT/8v4Fe3SS+jjYB0e4b+apQf/EX+lq9IJEZtFpDhye8u6xM54LppQ4yZVMA5FGObPmC
UJDpJUc4uy1Uvp12JbkBfK5PDSDtFl5qyyW3FGhfunYeMp+s60pUU6PVY8dG7eah7whWtcOhGKer
9XxptIRr+XQDDU7P5XhOh38iMJLgw473PPxvQTPruxSFH8ML3oKeyvf5nhEwDqqSj9l/5ayqwN7X
XSjZeSAkARAmWJvMcERvm/vFJG65A2Dmf519l1PKE0K1JWQESThBigY5jR/pGZXQIS3GC20OC69d
kP9zuM8g/D27dmKHo7VujFwMvktozUvdSLqvH06ZPnpFVNvoMBgWUMU0HBpTIK5SWwyRxxUPlfmp
7LXpZF9IaeamLWmSEapVGm5xZFqBQdGKUfVESElvvrJ8cMix8BHajk56Q+zTd7sYCSkgy9JCigBw
3YWKJ9iTHBla70YbDYEpVaCauQ/nVlYlcJxNQBA6jUoAZpzvwDxzqi0uprSQvckpzgRAvLymN7V6
am17fpiW2a12nl0lUXzDaym8LKs3iq2I6v/BPHTErkyjt1ktTqTSBAIPZ7MSb6UA/tkVRzVrZK5e
wpn4LrFRstShoTnDteRl/BX6+prPhsFxmvIL5GTZokQyUH0sKVLBS5AizH0ZXhd9pBTQsXrr5TNJ
pawRCn9EJNJb1rJ+i00CSWZJfMGKrfakE0IDp026zA8a86zIhWu4VRslR0JtACqUAeUNykg4GSLf
hWSRVcrf3+cZPq+ZZ0yS99Q+R29JmG4RbeQvcQVgJ9o1PFhHgcg1XBl22dKly5pWsiAEc2PVEsYs
YPV4/ysDCUTqrH2TIn35codWMYEs8tzURrvoORnTI4U/fHJFCqWpkzq5De2J+4bHBg6egBA9KsGI
Y5FhAVE0VaL4gxwU77SUec0wrTVE6csusR4dVaqK4cUQdeK6ZL2vIxyeY+pGQ1b33ZxJE406lR4U
wXT7QEr2xgoBF3OMSbmCFqUW2yoiv5cwGiURqAUIELCeoeVQhCMwfNe+ceiPayP9Z1g86WdIsYo4
oSQQeElUm63sI/AiYAPsmZ4Kzw0WroR/Ua28fRzp1ZuBY1sQt/i7weVotVuHCaNjqHkY34GM7b5F
SKt50EwpH9haf8Ge8DhdTjLFWKpXZRav+GD0GtFoSXeS8b/Mm1/nwL1xSlGwheniTBT2Y7hgE0C/
es7uwbpalOsPF9pdPybUO9MZ4ZRSfOKRcsNIrRvF90ak0bW/4o5l9h4ro6D7LO6TQ5XtTd7GcHys
vl428bZmiT3bww18Qvp99cV5iZGRCwSgbvtWTKhUQBKmlZVx0WDyjJpjC0/CbBUkWEIP2RUfykMu
hXec6QscJWuv2/Z17q0pB6LrTgmVdapMpLtgOeVQzksgaI4bUUbnjElthtcwEt/ipIeLklKQwGeK
7beUPr6f2aX+s9T+B+O9IM9N3zTWAeoJVkWqMTzNrKXKnG3J0D9VCn/HK1mWMk0MFXulYIlPzQ+8
U7XzB8UdZ2SpuhrJAGKyocoRRA/DiecXV1ra/oBbiW+OFWf93hS7mJ5/2jSxCRFgikh1hCSgLoN6
RshXBEcnXjpaBEqsbI4Gn27vrodUYmWnb+H32R/WFRUFdX+LZUfCCFqoLArlh/QNjGfrBp55MGGw
80XHMYzOph719gf02DYCKIW+VvCEmlDNyJkBx178Mhya5+NVdpSyGADbLCkjGhtNpIvSAC+fXQXy
yCe1x3dbZBw1NdVzbWUBCfAo5SG1oDqDi5YO431peeIguubdsMZpzXEtgb0NivptXHGyDQonskkT
1+sN/87PoQIGg5G4nl9qgIKouaVlDcYmf0wZK8JsCoC1yMXUz2JFzdaLSB+KS9Q+wVkIppYAeg+C
0fPHYUyoNgNSHcY9jbWyZDX+oPia5S+mXgDWvIrjLfKQXpCa6oMxWxosKlsgx5jm5ubnTTOoHeSZ
ScqB2rN4+/pagngqtgs7sTbaO7eSaoz4hqi4dRNkMZnQx0svgOkpXBUSyVPW2IkhrYu2qM3j6J/9
A75oLGoa35K0xa0QLuxgJlYmwjFHEBGAjXpPEMAS40sJspJhYMUZ7kaWurjXaYnTganPGbkP67Ba
hUVyyMtqiHYRiP0gaa9+gl+5noAp0pQ1K97EowSp+YQYJljmHnoe7JCNv0TjtunQ+2F7SByOcf+r
WEkqoagb0NUlowd0rSSsPlpyAZZhdZmIjg5epAAL9MoFujWhIXaYICf/5RG1KOM3mQ4n8iBUffXq
oTwS997DuhvR9Q84GtgeKxZYaOO7aMyeAQsVJxA3sgpMGycwPMFYDW25hJeawyVzse0bP+163xcG
ktzazhY3gNVXHT4DSLnAUDjHKWUeRQxpHVSe3NKuoPdpwziE9Pivdh7tQhkghEcWNCwAgsA6MKfR
MdgyAmEWc+RIcy6vtrOgQyEHZ1Rdg3iriBypgI0meoFAqjUz3nliDt8+LI4zEKvevKIRfyUiM2kn
PAiKW/PvkBMnUH3HcXEsAiKiviVdiBRBHjjvH4cVtxR+Px+heVGfNF4h/DaHNQK0xKxKxuqd7P6v
VXnY5d3aAi+r2BPAUaFb+YcNvNJAg9J1bZuytVRGiXi97S/xu7rS8GptCeSkLYKnKDXVBT0Jj7ri
aFIIj4mRKbw6i/3mnIcd3J2SylVENw3G4RM/+nujA0AqjOq27vWEHaPO82RYpbgrpBlYYooCJGcr
Igzxi5u/jISAKPl1kNdL8DArOCv+xfqVMH74oo9BJGBu7n/2Nrlno8OqMhUid77KiUCFgsRUkYM3
Z/gqb1txPYdl1Jk6gAA8eoarNJAvevX8wk9G0clFMZPl0ON7ci45CnMiuZdlscv6zVO1nhaLrI0g
+YInvxWZPNk8I8jocQl/1139d1rMIU1DaSxDn3hSDqxOrAqVjgK/ELNs6IIfWW6mcIBTrw8IthhO
g5HghOwVhpAsiQ2K/pJ+EgTzN0gxFIdAax1aN2WPXijNRXGR/ECl7BLmg5tNnSglvXwlojtB0q22
Wv39waIEQ83DRhRe75qIkzoYXBp98Sq4Q1u8XEBqNotoaQhiq+ONAPCHmJ1bvbPIMcesEr9QAhd0
SAKsiNjZ1y0h2p8Jhj5I6rji6fr7yll1CBMKDLINmeXG/4VwrWFLKRRI71/QBBflzvpiW7yAYNcm
iFwD+5Vz4xYhwOjcD6ft/TdNkK9M6YiGxDMNsqoYsYCt/IWOy6mrg9ZUtcm70gxARR8jZh4dm9Bg
ooI+uHnnX7XsTxZLsfJigcqYSta+YgIVdrUl9YY4wyiOuBdZKDxgoeUD2Jhk4+UdJYcrwagIWjvq
634DUEkHN3VVOsiwt4xLSe4kp2pboQuX3xtRkiItd0QDpzYg+y/jHY9y3v4YV55PRw/WDsqXI5fB
z/+ejCOPvd+3QDilEKdBWh+nHq4hydbrt9cddnuMexUzvqnNFPQzcPWGI/oqMaV6GCP6dGXZ79um
sXKemILhdAEJq7yAs3erUw3vtjck4sRQNTox9kQmoH+ngaFtmQApElm/z6C7DFOep5srYdDeJ6cs
BIt9iB0BJZQkI/E7itpc3K7r8RBgu2ppZJQwtSsSX2nfQWYdUEWqxa/YgQnV5kGEYc7olX9Wl3KC
ZCGaN6TBJiqXZS34V7W8yaUbxQPHP8s6Gd22siaTAPIhsOkcP1KkydpH/9dTzcl780OnlA8sWL4P
uHe7zHa1QboCU44hMwU4MAYng5GiQha7hMAa/yOCIgqCW+DiuoRK+gPlfHka5+hl5OLPhSmvTORs
v48/NqP2HAEl5zZ7aaUmXh5fyuS37up2ubH+Cd42wx5II9xw9++IkZG9VYFfb6nYgHfOiKA3+mGU
NhlwdUJtA4Z4lnjQMPaGnmhvlWvQCJItJgfbwrF8G27hpLXOSVml7adJfUIxSmDLsX4e4ZtK9er5
ujdbPS+fb4dbH9i/vrP9v0sj5VONFxK7HuLRvH8BcOzWBTgC/mw1MNm3kR1eA/oZF91wTzjatbnD
ZgiGJV4uNSpQWTZzV9BHxj4o+ZuETKXNViwbfh4UiKFfBSQXFl0Au3TVZb8yBHswf6xsPqGjBYWo
mrG3OElCtVPJ8PQrwf9TGnduVivKCmcEs9v9SVEHlq1MrTJj1lVZadoG0AnnaKApHdOzhG2RfJFM
euDJ3N/aU7oh8gvuQUBSLfElO1V8Uij06KK6PuUXm0O2TBCAisk8Lb+nzkVtDdADIwNF3qCmoUzu
7PjHPaICGTmPG//Kkg43EgYIEtMjyUe5808QXGnSxg6GkTZjxy5CBbCR5Uqe13LGu2CIyadZFUFz
oqlXnb3CJpirWL/mHrVbS/7qJnqiAOn+x8mLdKuT5fB2pKg3PwtAlt0/9Ynrvah/u/Xbpvi+sEis
/DOMrfqNBN3X1/zzaTGacKyZsj559CDLe0ENz+k4Q3o9wACwrOrQOxIz/8wBKiLTIOJGIib+6R0D
wsINp2otbzzVLL2Wdzr5UvG1a5C08HaM7+A7VzJaK7glnGknfk1Bk9baNH2jUdWrCjqODQESprIn
JkOhBVscvfXpffPHkTFUq/5JTpDc3uOyol8ZodO3nD8ksmWc4aEkrLfvOVlbPqBsZ07eLFk5ooy9
mbn14uqdkuXR2dFBdWz038RzfiMRwO7pY86RTl/zGym1XG3CjDtdkjXepp/69GrELGYBBJrGN6Nr
cJfUHAjTb9EJr1ItKL+EaNdnag1azoX4mysFF1DN7ONdzIqhK5TaQtotgn/0Qml4+VEJu5w5VhL4
xOBLTP5pEgw4GUbe/GFB+yzCz6i9+P82a/jN1U85tTekl9QOI994kF/AORd0Zz6L9fTQ2AQhW4sY
PWIDJOEYEK0go1wictaCFrJWVW1VnYXImtY4Eo6v2XS637mu9QsOQwplRilnrZeoAJSkf/BgChqm
J8wvA2jNqzBfzSk/H/vq0bmvbm04viHcdUAvBR17uhzAmH+AGv2wCOnjCxHu4jC7jhNjO2ycT9Ma
nhdBPEWTpuBmLIs++7MGXARYKlqnvc7jgmK255WQPSIyKl0iIEAKXdSEL2rrVaL4jBP+v3Chu48k
ISfapDqm+9me7d8KmXFdZKqQmJ7eoxJKIo0KLzoxtJsjCowOjgpB9etlrSxx7wqbTa9SJgLVpjzv
yqz8fb35nFKotI1XTOZ19B7vGLAWIjcYOnz6rc5DOKiI85j5/lb2DerzJABkBG5zfwsKez9dvDog
UYzxOsTV11XbzE4U3Le9FfT9xhbhdFX/AVXTqiIWGVJdpmczN70uVX6/z1z6al5fOz5PiYtN2JpW
SDqDoYiSdJXiHhkPFaOD1koBI8v0F+Yyd9vxBwKEX+bco1tNFW6JMpk1hOc8QDbmnIQrJhH+uo2D
LYfE+qNnEyNW4GZFqc1Mv4m5jTUdq0m7kuuq2hwCmZrBUjRZ1tcHKqh2r46G15h1Mkqudb76WplK
4BYDshif0wee3FNq7+Hb25ui4j2g8UbF9Uo47fgwYRShLOUqGmidJumjsCJqLe3WCWZouW+WWEef
d6AduNmFr4OygJ0xIPK7gqzLpmTnXLr4mFYaUygnti70R2kCFVUOCbhCDWfb9g0jDdrdyt9aBn7/
hzcVXlJIHofIlmJisl4drTHMWLydNXzb8rVob1PyFqH+kitkfHTPWRO62/WiQ5ICAVk/c9tcOLFt
HdGcvephw4LRtqzEI3qHXyuHyaCWG7kEhO/FEywOZXb55aM5V5SB8snrrNeamZ87kOP05uFwigLb
fOrUilW7mVwdEj8pgVp1X5uLQzjd0Ut0h1nDQGX2bcS65gki+9nZtDd207+6zpRV/l6SOi3IROxr
Sd22eOpAWOMULSiXKfnU+9PZSDH2SLeQ5lvL+4IbQO5Xf748dqSokgFArfWJm0Bzw2VJlvOX/afK
j1EHcWkpouDl8x+rn4aqJ+24SWX6ysZKZGh8Fbqrh0bZO9VDg/Hnf/Lm5M6n4Q6TphBlL7LlGaR1
6bmcB8ju3abtQihT/tUawvUY77JAALlF2cAZDx5kWLHPuXBhlvappJV2xMdJy5mDeYAn9DnfXc4g
gjt1WQtXe88hY1NiYiuiHbVSnL5F3w0JihTOUV55c6m2cvywvp4pkhY5j+m19JDeKLNxWzb/ROFc
qQMZzvrifoh23OpGft+fk4kqPbMhqyTinyjba3z5ajj268M5vVUz34RXG6CZ+L1aFXZL7gkQtzrH
7Ro2WuKv6uF0KXEBYHZIQcqBba4Xjyw7Qgs2gnXBF07A+NOFpo+qfF9MwzlyupLCpM0EcUSUPRqr
9S4EnLtJrfrqND5vwZzUqpCSSD2yruTSzt3ZvL3YoeedRAZZd77LpHJU/jnwfykkuI4CpLVjAfI6
cMqqBn1PPtewlbn1GajRzLsgTAgmjOBtDK3RlFauXYIyhbZ7zAe2zWnixs3MUu/27DijSZO5Wufd
eYA8fsrkW5KpBxRMZZdDkCCAxUNKSSYiRidcun0QtrnmGzsIyHPYgtpBMxA36sGmZhjo1grddrQw
hQ0UoWUG1cYRBLj/WY9eLD/aYvASdfG50weKp+Ipqrx+wWaN/E9ebM3trzSHNMIzHrzMsATNvnTE
8WOl1q/IE7kZ6/XJzJzlZ+8MCuGkrz4wJmrS8UBNGc8orvW4daVIhLYjgxY/sZYYPE8vHTeLQ3nn
6iB69v/H0cmXWndC/VbT56IDjWvsuoQwAoYz+mBXko3UjbqlTboU1DP2MNuLAq2KS6HnUmkR6lNo
IoME6+dD8E4bU2Aydvk/mwymDvwzyVS/c16TGPUyWSZZOI1R92Z1BFIg4gsuVMr2IL/roJUfIUBa
Kh0JnstoPNMXPqYUlq1P7FgI63CIPWiL1ydKZRj76fnTVWDoHKUQHPje7yMYfLvPAd7hFZTt+5OX
4jQb3DsTzctpqul5Fb92cD/oNBdDT/a1sTEtU7iUmSMjPJkReDfkmYBISNZyffUN61YJBNggXDib
/bvC28DjVK+YgBqDOPscByO6wM/O3nlstq0OcqmoW41GFSPYk6JfOM09SYvauIcI32QE9Xv5gndx
9/+0phLaim8lyscGjwuEWHXqgrv4s7vZYwyMLmL9PSgYNMpIM41j8FWBinZqcXO/BQSNSxHK6y2Y
XzwB231hl9MT5iwB+WRkNer61YJsy4V5k0IhWObrTXwakCtNom54QSuGrYsvV0csp2cRttDCvCFd
0z0YfWjZYNPbkJqdAzKsVhQWdnnlo+lI+RNyTDa+Elz6i0g53dR5d0/HEL6pddKMCnZtw02e3c+X
Aq5rFeqtClIRsVDohRxpGgUEf7t0GG0B8BEwnbkFSgRLjz343kbU7YJfS7kl7qUHaenReS80BkpO
RDDWFlHtu78qGrzdaoEDw8vq5z5j8MOsDfShjEbIQus+DGRlBD+uBcZHAzkp7sCHhD8JpdzcKWE0
JrFkPApAsQ83n3ZqYGuVY52POgYta+dbXIR6bONzTSGN2UQ2OkthVmoMYSMurOHPhA4RXj21izuo
FJ0+LyL5ohzrzDXAm9OgLY5Wb2O4atXb6mrvzOb19iLvKCq6Ll2C24frnO8C5XeS4P0rQR+JJJ7V
lWb8m8HZHKPgULrQbTAIX1/Mt1TGimrNi/i8d+4EgOoMu6HgwchUvEO1P9/pj8qtZXSaWpkV+W+q
DeUaJGPnCmazBPiNpLdPrPRTVO9bQ3UTIyQJiPiFn0rwEUMaKpWlPZAmXMQMwm4Uz/xbQDo0IliD
s2jKSmcxjTuqz/Rh11b6fudmw6KWXnpcnCTYPIvp8hCQ0i44/IKRc0iitElV2rn1N4vFuQAmOTH2
dbznwpteNc0RzQAvwMSqda+HeTlsvofDK42fXnK1tfl8OWut0/nacsMxxgLXyCa34DfA3xuXfefk
VCNBoLUQb8jhB9zpRh+eCTlg6aWpEf4Edmysrz4c1lIffL9XbvbtXxauXQzdY6hqbrqeY19t+oxP
tS4cDSpMWPnzrKbgp99ifwu3J9A5PIGgNMrihTV+TPW8r54RmEDTi3hiTRC4JTMIrLS4proiYQuO
wmWfUo+7yW56roSOIOGBol+jOvkxaURLXicazobFe9IualGrpOX7nuVF8oMmTLbeB7DQbDTaE+/5
cTXs7DJtfGRLrf453uTNO9V1Tyn2qxAXynnOjhG5bZwh1UTv7ewEBFZHm2fndVC53B2mq4vfUv/d
KZ36y33ibk943gY0GICMJX6X7ZLL2s+Td7W92CzRZeFOFPeEV08HssrljDjXVzZBYmyJS9q0GWUS
D2zuPxUXMDkBqbCCjegEvThaVPo4/QNU+sD6SN+DBkmzA6m5bjAGKL6aqK+A1seC6aGJqndzBMU2
meJmIvUhvkw65HYdzcAeEofW7jdj0rbut5B2JMS9FH0VQxDXhD4yQVv/DJzu7iAcYRYyDylta74S
+BPEIeF4A28Fdx0i7V82qVE+NbCGt8Ui02vudboB2CxyePRGRDWFX+16GLbdfyBbtR7VNe9UYR8C
YoD8d828Up434WyuRmSbHIu0lLY0ka1XGxWu8l55Omd5z5gUavoeZ89oww++XriEj2kkbKKZ0pzC
IZx4IzKPcrcOKpUSLW0ZKYvMz64+jzXB2C0wqvf0S3Kk4fcTk/uVpDXnFW61I+Q5tc5i7DhwzckG
L9mJn48qvUStXKei0fhCeOkI22GmlOu4MjUdZXLyYoYfhoettTvL8kG8ZvyZJp8fdLdSwSdkl4Vf
EN8Pbpg+tkxkArDXDQAF4cck18bYqCTQPPR4GQ18zydxsSlFS8LKGeJI7sH9qDDuParzq7s+0UAQ
s6p7bYtMYA8Lx6xm8Vzepouv4wiVdqvPoJ4YWHOPhIltkES13DKXtLMIL+OJh00iMXioPEbQ3A8J
ZiMOJQ3f4cH/44gveMP1yzE5yUTAJtq5sd/Sq4YAubuT7TJP2j+PTM4LIVhc71jbngzosSCwC8sp
nAJhTItyzty9zCRTM2gepay7xaIQXJDMNNPzywrBPF4A6GKdXM1Wqcqc0hMeMOBoxLAWyP+rdtU9
IGVWfBFB5qQOWP3fO5TQcpgzq24Hz9cB6z17RITXwKZx7qaJRvw/vCHHazQtYYMpWhjM0FSD6LWZ
bVQXn4fBY+tkbt6aNTWIcR06lEDO1j8rkiHAJ+GgEV9UaaCinOL+z3A8PVuT4DhvJHpN70y4DoGE
oor3nc2WslHafgL2ucDj4brgVmtBxvk9QhicQac083Gaj/2okI5v6CLCdi7D9TqV2F9Q/4703Gj9
RfbEAEOJ8/MjPGjRWU4hZP1nQM0Bo04UCXjVFA+spT/4Y4VJG3vCDdY9HxxCTV++EbkazA3I5NpH
YRojpdbektLdck45j/dCswkwSojNe7Lxuz5aj9NldChmKF9agaAD5yJHDvmmzIZsN5NNbnDLQ7zQ
YQbe39HDsSf+4146r6jeIPVAk4WaAss6uItRw4SFbujPI6YF3P19I7GXYQwa89/eOVPK1z1NzlP2
NGrDuliuI58/0Nx5PzH033gdQpwUiaU97ADxIXzGA3v6Xb2Ey1lOr2+FBMrnzW6+rqWsJREhZjZt
jeN7qTzOOGmFT7kkooMa2kfMDDSVfHqqDcq11RimAkkjZ6XKlmXh6+VEgyi+KluyXFNEga7E5B86
ljrFe6z7JqcYBxUXlbET7sFGG6JRgmW+nMd46NHNkYg1Udisf7BaI3IKKCyLJYeKK2bADhMxel9B
MicnsXzxR0G7YfFVQCc+PnZFBiDKuTinfGmSSFSVGaxtehsYzYBZxrlkzdFmPwtsFzlQ1CXi7U5L
oFMBvsA8pbb7dcKylwolPAElPefDQcZ6i71Oe6jqvXLQIbLogMcsJf1YM2eMtSJKc3eDmhWe4LUp
eG6LFFCR91aIt25VPFlZG7HMYHjnp6IvTZfdN+19dy7ys8J48I/M9N3o8qP5BbEEu6gWPNxPLg2Y
KBuqO1hmR5rJOrUvCvGv+r/a8UiXYPEKc1rs0RcHvuO2pWXoLqysM/hyjoauB3Azi52qgIZ/DmPf
v9NUddsFDghv8ag8gOGkNTOq44jUwcnrCzO1XnW+9XVDfQA5xBhzVns8LLPgb1RywkyUuphtCYeH
hI6FalYbj/B06KaAO3FPVVZxS1Bc1ljZ/rn37hg/NAj/ylp1epoqPw5FXQ/Vf7Rn0wARymFx6Jow
X98Ky//WIPGeKbxMH+jd0IfZGMFYE/Zqq3t6gMltnpj9eVAAlYUQYjNK8MGbxLbAgS7BOriEArpp
5zw3x1/djOK0/hFBMvhHIoK8JD2N0Dg2vj8XQGk3WLyQivMkJb5j5eQ9XwljIjTyZHXbRfGtlQyC
5oRQcBGbYOcxXS1jt/1cb0pRmBiNzoSvp46zweXE65MITmO0ZLH28asmXLgBRuz1oj5Wv5ojDAC0
c3jKwDHtmoqcl6xBEVo1D8reXel+1z2DbDVKEgvwal9JNV5af6C0K0NyEpGCXQ8fuQDt0t3bMz0n
NnRtuzatPBS0P0ffe8kCacXmQ6HSLITqNPZaZ6aT9FPlYQJ7Dw41+CZfrg6GgU31Pe5wcCw3p3+S
L0jrnxe77/xN4jjkdtMN0wet+nK6jhZ5/6bKJjtnOZWx4YGn0n8XMEK9bVrc9g6hG6z1g0KvgaWj
3k4NZQbWfwVVzz5XzJ4mr7qOr52ZdfHfUhw1QavEWoWzDbpO7XPKMH0KL/Si54QzZYmKDMEI4ng/
c2biy0FC51YSJYadSFCPscV8SjGt/A5EH7WVnjGQdJZI4kw3TKCrG/IgEc/By/mjV/o8N0SmserK
ZMiRuAQthQaF2AxbJ/f6ho3SNHwgvURjNV0IzjDo1GZUthsHUjyFjObMErhTyGjMmgNi9HLh7/q4
ubTzBa9Vo3So6/v2LbEJN4NB/pBBCePuSruIlTuslo61/rr8FYQ2z4fqxnuUTIaWRADdS3yNUdak
hGokaHxPL5hUgZoMvl/xJ34oQBtiCSoG33RYpEcUc+K2cbhJq13JCEgKdof71kfptJ+7c5bovYgL
k+0wlVcMpcN6L/yq+x44Ijlcav0vugObeiA93g0vdEmmgEbbb+kRf3lFXyLLxBczyp9FkEbiyJqY
zFg5x5H+8WGI6n1+MSK5c+iAouEAVRwSfgBxhojZQ7Px4ScE3AcvLPLtrACAG6Vhwh6SHZWxLDTX
1RaXOVEfHGZVqCbOaGWAcuJHQ2Ad5xy15kEr+/fYjjbQxAkzLSW8WXOhTAH6zBDgeraNTBaXIcvB
9n4K2PfeKquI8p8yrM+hxAZbtANrx9VnbbU4mBVIwV0yDFCj4fQDo4nSJNLon7+toit4D03sSeuY
vRynSt6AthPG4FGei6QdRpDfx0k+fNsnO62MbJ39XvTPIn30+jpBnqL8HiKe5X+W/BbVHjqgFLEy
sRBSe2Ay4g3mAgszrH/rVTCfpavHK43w4omGbX3Gra6ah2EAgvQxJAJm3T3vaJm3YNSqgdReDEK5
UkKgWueGauUQB1ZFgcEM59L3fqFh6PJfh9F7Q3J/XMfmLO6bu4PW2QDVOFLXxHA7nZmoJicK8pJw
I2nXZ0gIkVDTIimPqGksnLw7vm2wcLFrYblBWEC/uunCPXXaBUIJ7ezWxXiqHMamNJVJcSP5GZ2b
xfW0VhxQxhdtxCPSAZQOonmOLOkB7Qu5WFpvx2Xc6nnETY3RzBPLeOh1Xlst84A3TBY26C233dYI
LEC/MkS+gSL+DgrurbvoMdXTXRDoSCMK6M0qnCQCePeYv/bci691Nj8m05M9y2rMvJHdG6Pv0hkf
1YmoKe8mvWcnd6zqjDAQCw+1cN5uzJRZsgeTzpkL+RnHsqqIsAXHfg3WeTF5inXjnf8NjRuDzHwj
8HVJM1S5x9eLsj+ys+oY5GNESRaWsnuP+byoofGsBl5f802SUwBEfoo5fRFaiw7I2B9yrE87Hrdn
fMh1Ks6/ISQ6MefmBdxxZPEAGtDqhpDE9Fdzl5v4WZGpsgAEj4KK2eDq4goEKX7zyPI7FV7qlC6I
Y22Nn5ftOWUb4gSKD67T+2hj6IZHr0CJm8pgwmfa6XWZ4oJPzQuodAQCKekAOq8ifR9BG3xRbqAS
oHGj11qLW2ceF+AoGHuqghmJ3TuDyeC8l6jY3peT8Jk4WuQgWDpmaSbtanQrowIKvrl3SCHDTVq+
toeEru3oFsfTHWoRQEiHX2xPLYFZwfGO1e6vJmjBC2ZCuBTtMBFhAC092u+EvYPJYW5jDk7cuHG+
RzpsTRCXqjUpwnqHIO2wYP/EEX2nT0AtpR2A10PJTYv7k36nEPCGpRtEjSVcdTUZl3UNYXZ0oUEU
2ywCJ80k1KxmsEz+NkxmcPh6/rxvIMEKDzdg5FLb8aQRZgO2DIl9/Z1vQHuDYc37Xtw9Da8szszR
iMpkUs5J5S+ceA2kAQpszE8xAUiw3aBzoJ+ofRI0vNdceS7KCSs7wESrAeBf0uqoDe08oxdoEtTZ
fIbK8p/UUwvFYgNHgk+0ENjNvtEC4qwPXamA2PGCXSSPnyZQpRs+yppTd5s6JDqw13FPf4/gVUni
TphbQki5APvuw5VUrRoGVVydnGMDrxWEDNhjL5Ngpelnjy+Y7vrzFw/9D+79swmrdweetNrpkeG1
oLa+ekHIj8biOwGafWkXLiu0Xu4PCG+swei5DLGiIewkKgFryNESV9E4XyVnAe3U2XFGAb1gNrAK
tIYJjrxmCjMtwGn/MoX+jN2mnl9Hne8clO8ENzInYXOckpLn3fXIys3EAIe8MQ/xEH3s2gmwZ85V
nHq46DSxBkzwXCGLjfntWuIkyQCZGbArh+X73KpPxHMwuu9H4sUvDYExOe9AeYrE1LMELwhYr1Us
3xdtprA3C3Wc0/EI4HMb+Vq7JCC606VPn8vLEtwbpg+BrgBu70eWYUDv2wbeHHK6IRkPwbPMQCUd
Cb89J1qU6F20/FSBdYAC88VROB+kFNxiyxvo95B9U+3T4qLa5qEB2cv+N+y0B1JXZ8R3DEO0Ihuz
YsSj4lnGumIATciqpoeYPe5iAyGrG9VCCQdCrB957xAL5dTR5Ir/XTAbfWX0UpLlnaXn0SgHyODJ
M02yj8ha0YhqvbGt7rq0ODJGUuM6pkyJ1Di0rx11IryldkMkhhG/tndbSvCcDAhqzafy+eKgzWxc
EotCHRMwQ72ov7pQ0yHuXD+xfbEnS4yQ4CJX5TcdI3QbVf/w/sm9sxocQiFDJWM+qEwegDaruQNh
9Tnkm09Wu3Vkcgp/nTP+LVpBRL+8LjifKFpwhFoD0CAH3Ijzub9YKqNbgJAIgw4ijjh0ZiVX0XCN
T6sZ0jZ58mIL5fml5HMJIoKbU+rG915skiTGtt+crNFvh4fFhpLgf7s7VBnJrag1fbsiHIf3Enuh
255IGSP09yxb20MTQl5alLMFSAGBNVvKedaSJwK9XL1kJdYTBeJ0dG4nX+8I7pCbJXAQQ4IVh8a4
VbcOQx2KUtxdUCUrRFHjxzoA6F4R/6qdQPrEAn4lQ5WvMBIT4DzM+m6YiHRjT5FfXufXNWlFfJZ/
p+uI3tX0OI3ZJGPXdbdksi/h7l3g7CvAINQkwcgZM4K/Wamx/IRfd5DUqVCxI7nhN73jeQW4UAvI
7PFKSKBitvKxS3wyHoQZPy3vM6NdgCHnUbFUXv20VFPLGx/wzjiyPZWiRI6HgcWVOIx1vYTTdZG4
sYeQ24GNjbAUm7jCr04oiXKFMGuZsiA+O/CDT5Xcr686dfbgU/PuAd3Y8Dr5GASQW1vsmkgV19k6
02WpxiUpKi7A6PXGc+V5mFZcrqyLj+9qW3zmABF8jy31UfSa/F2/AQA9AbCTH7/NH4NVBOIqCqYV
hBAvUq+V7MV9cZgkOxwYvUtQm0z3pakV1dTjjblAJSduCxEHu/xHxqAqFnf6hGUv5r3154WpNE24
m0gLL0jkxVdd3IXxVkjc7789NsNtlPNUvzuruU6WyNXe8Y6yEE1Q0Amlam5lldmK00BT+sAUbeYO
gB0z/Z1B9xFC5xzOcoGzVUobSwJ2vcO4Qh1qTcb8vo0gHMuIwBIrO2eYRc5tjqWTezoK15+H7Ocy
nqxMygCDfO2+yGqYp/OKH4i7Nq2QXpEryA7HQK/9lqCrsi8pwarpUwM7Z582NYm1F3qYvxwqVdQ3
QbijBFw2Ji28B8fcpPtqi2xsHRyb7HuSn+rval5yn+7O2rwhIBMXFzz6QbaECs9K1J419yKGFOCu
aHwABSlov634hYAUzY0pNe1osZD+vtdGcnh8E4zUdgUQ/oMrQk20rgEdezVEXCVrE1QM8g8kzInV
sRwYiU3R0kakQL8jRnvKYEmd2/+7IVVQTAtCxcFsISrQVEp9XH8IkhcgEPK/L+SwYdlARv13wg/H
QBg0pkkrHhx/xNmjO+2PQ0uWQY86xwBZJg0oE5y1nET5NegFmmX9FYlHgJ5E/F1ETApvh0KZDsOJ
NJyR0qFeyV8SyWOL20rjy+i1QWkBI/LVVFd78kFv19X1z+8NvgdiDM/TbMzRTHHV+hjLPG2a90Uz
gz1CdR0/DdeV0H6ywZabAl9VbFkE3QW+v1iO1m8QKP/LKb31QSTta2KwTKyoQznhl0wqiQcIcBiM
6JPTyHyXQMX6EZ/6BI10qMiAYCRy3IRmwlmdPNO0wcwp0doPvhdQ+SM6DBJ4/yxL4EpfxHoLLp74
tExff4UxWGYODnl+LY7iOqpZGBJQDIETqo3efvSTn3/n3Q71dc/AMRVnNpTI6Qj6CeAsgmZqoIHn
wZc7MHatTA72k50nM7hBY5/B4pOn/3Jvyg1p/th1sNqxINPYxgXMBQg8D1VczalwjzxxNwbFEA3m
F/1rXVwLb35mf9FcojRFuRMl62OQHerNFDqTbVONaQpt/1v7ypRLqH+2+Vn477jCiJZ54uthL+Ah
x7BVC5kUoR2M2nAw7lNXGmPrSPKg9RNfLXlQFVH3sMxNbKRyo/ww3omXs90kO84jTP7HV+Gzj2FE
bPPTkQmXsMRRO5dZBNeO58EuBhDsPuUh0mtKTwHrYMTT2idNAZZW2lMWt15XHfS52BfTmR4Nnu2T
I5fbysdX0ldGn5GUjGje9Mr5qKnA/r5AotS4ZK9Xolfsz9RnT3F2yiiiC9RqlQNcozZmw4v8m5i8
OBvpr3llZ3c5bKKGR/ZjTz2RmExoL/7+fHnF0k6ZmK5MaKyBnML9ovGa/nsyhuKiDvQyhngIohUW
hs8WF54K3Zv/LLIAqcmDnW3WPQHkCZkee+LRWbaPcwOJPHgv3FhzspIBHKdeLaC5XDLUPam7xo+4
B/DievqlbaBqjyH5LnHYIExlFpjahQ1PAdhW1Aizvtl3911EGyn/8z1xucjAM/E/fP4u/jsayBPT
4TJfoc5F8LXGcr+PYnFlmTyRFkQKFmcva1eVx00XATwPGnECwnVTjK0PUY7fPT3H4aW6BYhCRy+Y
nJ8OVyNM9dSCuI8/59nCKsPRLhRWxhyP7fNmnXvixlfWaKIhy/oBqLqAQxZJS4cUVok6M+5s9y6i
4IkZkqMvTPR1hOJJac12FLIdIf669qRjsBMkMHggMlH4yEhfrw7fJsmoY5b01Jt/KHUWsUjcHkEK
Na7i1s0RRFXOIa5LdU+c3OtF/epQr4/lpkWzUui0J3xKluccdJGIoqf5mJUY86oOUzKGPJvqKOjB
gDbZ/7ItOFQmv3gGg2VjxsY/GZ3VSM1bqTR9t3c8MaNO9x9+pm6qByyloyZp0mENORSMmMKvGshN
i/eHCjP/fwoAVYeX3IVDYED4f9ePoLzEb0whkWtxY7ox9wni5swECc8bSHdkgAMSmjUFmjl9bOjn
X3X6AyC8N66FQ5zcPdkUDa6efgp+K7Czkm1y8Pc7E1p4CrLbZ3wHHcvMI6aLsVET3FyBZBPezCKG
iOaCzD24ep+SwHrxkoUHVQTcoBCCIoDnpiGAfHsbFioFnpCpCnscH0gtQMplHebn/AlxJv2DRlzU
q8kH3uJwcOfxifg58C0w1vpoMODJU+DSVoxWqCiA6n/4+eBGuFKD/Ae5N3iw8CTpSgb+pYPFq5gK
SIil3Z0MIAqe7f13MP57EUpAXSpCMi15oz4QdlF0WRcMoUaNMiKmLeVoJLfFRBdbWpVqXI5kiIRH
mDf9vFpXERkAOlS17UD1Mmp/dPPrDHyuygSTszEZmetpmKvvWzKyZM+qrrOI8d6pNjmTA3xvYkE9
XvNebZLIamE1uwjJwxybT4JQ2OwkApZXdNrcYfzGNhs42bczW3sc4VmWhc6mydyr+8gGCo3+ZQW9
fAf0+W+sZsgJF31TFMqLsPDEf43kQsAZXGFPrjX/zwSInO+cfuQDNCZ468KcbWOOH47gVIL5h3Ow
o8o1b5/ix5jhs5+Gj8gE5WbhKM/7OItp6HTZ7uvUnbMoud6pnhEYgOVK2v+Jcuz8iHYZiqH3wcLH
kpHSFOgYe6Rs1r+W4WF+otxteyjIu/sIm6RH4dtGipceAIJJwNzFOll/cNI+vTWtvAA1HYUxiLK6
HCwm9uwKpvRmeR/E+ry4Cq0FtZvNKwp7j8l/SIW+lVstQXSVT7sfraWAZ7ITsDBSaomsp/Zy3fkQ
NSEEKxKML5OogpFbY182pBBvzgjXAP2zvyLaAE9GGKytocNnvCHFPEcSWgP8GrYkcMCgOaB6F6F3
zwmpi2guQU3YVtvG5S1j6t33OnXJZbkgqLQ1A1nOJt9yUugZDddk8Rms5+idYynl5qaXrDlgqv5M
lB73BCdz0uCJceN25DeDgUWVfU/ha5fZ8/I3KZFuEn7o8e5L0TycV5QolL3O6bVJx4qYpgDacFWK
33XqgEXx39pufpEm4dSz2XLS/E0VG/bsPyh+fXIlK1MB5cHB8OBYqEvNQOlHULrHe4c+8BYSNLX1
Aq8NL5k9APtdhIb/y0zyB4cIl+EyxW+zUWxSfLjwc7gUY+92L2GAweoegiqvJ8hLzxIvykHquqe8
xF9rzA23vqiTgvTKq2oiHlyhhGL9xtGzddEwpq+yFNT09pDPkzzA3EN8QOMmcNBm+MN+ja7yzSkh
5UQAujDwOubeT6VvEsBoK58bgnSUOL5lKepwZH/GGsrMYI1H3VZuWS3KSxD05ttPcjTqVfEHGV/d
ol5o28R2RAoCYgmk+KAgrVZ+bojG2u5k1F3X6U95T2y08tL75xZ0aZa82Zk7JEd+8EsypcvD4iGK
5tjUDUyroCslzw2KCUMEGISV77Q9EOUnIKDiQNyql9C+QXmw0ncQ9ShdUCujvw82549wj8poza1W
lrZ267Mek5mrViIqmqetFHqBXLOvTDrsvABNhVQFvHR2qgttEqQPZ333EAfCL5EwqgXkj1tbq0ds
ffsbk84DlCK6pVul8Bqf7lSh/oGmgHIMo5JXGYxDTBuphnPFhshUarck0zQ8vsuwRzisdklPX4zh
WGPxLwAmJVhyKBuQ95e5Gmnmzdpd08r+p4/UDSnzJOVKDBV0Vb3qoj5lFpIxCp/5mk8HdunaeACW
y2gLBQNXGmOAG+IKujvbsKDszQ/pCq0jMBXBrRw3HCx/KeqTugBYIam2wjYaJ6KutybYqK7GMIwv
lSbHH0Aarjw6HoQYZnHfXdmvCDp3VEtZg112ffh2HHBI6BG+wwBzD2PtYM1P6joUJlJTgV2fyle3
hdOeHVRYULZsN5JA2ri0XcpjPoYUekd1IOi6fAVJBes/S8tIsfNxQj4jUVy3abBTHCRln3shDUSZ
7bu7uvA4cyDemj8bSyfMWr1UGgmWwdPnCzncxv6h3KN3ejrCq05RFPIUOABDUNHl00+bujjEQuEA
LFc//PkLvv0oGeq3Gne7KIcQUxiOwDzfOhC1zRiwlNJ9B6ML+glVZVxM3UefBfx7Al/YkkexLnLN
WiibFpPkk+bfAARsqS29KvRXlEmSaj7AK2YrfHQfv8qY3wsqmZu5717eNXFMt+eaj7pHnIBAEYaN
SLBpBooecZTw8a7TGSeB9cBHUqD0L8y4x9+BRhfSqwC6QHoOz3FPjdxqZMYU/GnI+lZ/cDnIzdqi
/O46Swuze2WXgtWc7sjO27BUFns7Xj5Ibwut0uhLEycIwbCV286cAHIKduCGXThuqirYv5nSzDNV
SrQkd1jtfDUWNDZ+9wdjUxtvm2ld1tdK2gEVUY+fpzzL21ClAHPSXQIl95coauAVXwX/DPlsPJif
0h5gT2CHCChby41x0cJi19J6rE4Y5Vx9ZGaq7Av8RjbHnjcKhj2CG+WXVH9k94JxG1lw9tVLlc4Y
LYd8kQQsQoKS3uQLM+/1k0SQLGo0O+RFWX0b3tIQbWDxtz5YTZ57RKHGA0wsQhavew5STEcgbdav
f5nAktc13W/CEQvL5WVbPekKitJ8sCZwsT9Yb1Narc4YjCTwbZVNwJ4FxUa3mmAEa2Kjwa3gaJ2r
Q5XKDntE+rP+w3G5B8ED/M8tSwVGiAHLglX/5mQR4J2tA7wXJPi/KvNuJiZIzghk2iCn/OsSgB0Y
/iK5V/dNHZ1Zq4baWL4d7Jb2pCRzGn9cWHbb9i3Xws/RQkfCIrQ6jggPWwVqqSsQlxVsXVhkv4ui
ADCrdnHQQrDHnj4olX4MNMEwTZuPYXcjNITaIAkcuQBLfO+YDX/5KbVUdVNTDTQ94999HizZlOhr
j7cwgtpbgyLsSH85++chV7viGJzk7UtyCGfMpcHM/iTlmj0OCjQ3acihdif32O8yXRy1Mr2w0Lxt
8C87pI6TrBXeilVnbgfisXtHOsdbU7jfWEGeQW2nv76zNtRO75z5v0KDZtEQS0RjzuQGH5OId6uK
o6Ki1jCiwjLkBuG4c824TCsqTufgZCYx/JJekZRWgzFUfkp4NDnmscmyJn+CPEu4y2tdiIQ0Z0UN
jAqKZG6YMFFlfPC1el6JLRjc8+SCJfcyXejSrW6vjd2/cWLqQhjuSLVQ4e/VdXrSu3XJyAmUk2lf
j64+8k16ucgUO6xdQ+g2Z9NgIKNzoouILFGTuX0K/veT3inuv8elYzDdPK4hCu24Wcg7Cv9heRk0
zYgl8D1eJ7vcoSOlPvwj7pEay3ZqFS60rohpDezbsYQtMSCx0Skqo/+gMUrXyDtQlkkldZzVwzwn
WFOS+abFH/FpP9vPooWv5W3fDY/gFWCY5uv0hRku7D+wrjvk9kdNfIzziqTqMtdO5hnGUZ66Z1u/
RBMTO3HbSARDHgCnGPk9gPSQYnQsIjUq7eXIcPn7krb7Y+6LJudEnOCwvxKSVGuQ2+7wGX2GXP+W
5CmDGDXqVinyuxdpBh8dFvqewvRsb04Ni65nYgtxZIGA3hUI3SqEBE+LJmpSKmPfvWrbVdLoWGw7
j63Hl08lwj3WUtbGZJRkdgRlYsVtaZ7o90YbfJQdd9kkppJhEh+MHx3MwXpXZ9vX8AnwnYTeKsPI
cQEWBJilRa/2sFvwJvYjN7m9ICjWMHBKgovm3PZxvZawzyOeYw3G6vDhGZNgNNQ6VsksX7g6cwUl
/tmVrKr1hFaBMY2nknLouWF1FaCkwMHwJof3HcfayWj5T4zVbqB8zWh4RznEwn79VtNN+UI1tLxa
szk3wJgsapbiAqM/79jXoDFDis5Ts1hn423l44VC+hfJOkIeOsx/6FfrMgLuRll0v1iPLtlh8Hwc
C3rXpiwwSJhcbponc/cJWJlawgjRIWmKYdlhoyjj628cU4/+rG9v0fiPwKOcA31Zv7hZTrHpFWsC
HmWnQgyDDCW5oKRJytRGiX9Rb/E1ABLMBncZzFuL6w/TNsPjp/WAWDbiiufvFbc+KW6w/UKRHrkU
GOyOZuEKd/tLqbtCe3Q+kmeaGyckVpDd1IsjrDVVyMzomQxvujyBsW7w1r9fLySWsRve9oVuQNP1
tDV9T7yQVWiGbNtEnZhw1Iy0SaNKudpxoaq7gZZ3dXTUSVeffWo/gBywsSwO5kt1WcyTuC+fBqD0
uU0UhVpXyiM7gHqNDCrVwhOqh1QdNNha6/xcVFIueMZ4M79OeNco1lBtB9cSo5DMXGmXWy57mSeB
eciy/yWAaUfxnKnjjbWzEXl96NquiekTmcAxEp9S6RyRgKCsavVOh5ufCljtlCMgfqPW9mMgzPxF
flhAi+kBf0pzMGBX7x/lfIg36tt5l+Ve3RmefChn6ycnNiwGi7GmOczINY02jCxg0Obx9P7yhcXv
U7kjMsNDZSbhV7IWVhf9e8kaduz1HsupSJjPBnxjCc80sWL1k5fAkzbp93b1vVZqoxiuMssTJ6+U
r7U8cxc6xsIgZ0EjBQK1HkJJZzofYqUl1gRIkrKyIuAtBu6+AtZYve/R9evok2p9QAKldmtwLUMP
KJR4i4Fg75Gw0ihvfFMZa5e5VTFf4tQ9IecFJw8wH3hNmeSONq6/12Numwn7GWvXwVgn/MQKtC5B
d846DKlQHNNk+EBDSEbnIMVE/DeylERhJLHQi0PxPf4e6RpS7m4HlrUXwckM9MhxRGv3GY0peXTW
Ph7fsZ07zwEE1vbNTE0OHZSQZsVDdlXx3IsmTu4oHNyOrB7W9quFS6gHMKVWq3xbdy925ZO8DZTc
PWXsxAUrwGIshgbd1psMbu7MCLYwRiGGZUIZCt99k1SLSyoCFkznwbjyhRJ6CU1Tiylk2Kvwl0/A
9yk0j2RWl+jM7BDehbiMd6fo4QOwGwoo/eTihI/ZD8MYshGzMV+Ysg0hKhKTQ+vQPk/Vh3czZfQa
MxXcPwIxHhzMQn3ohBveLGUjyRVuQ2xkaIFMUqznaEB4M720Ohi5nD4phLQNgsS7R3QqGroLLW3u
vtUGHg6FAqdAZAhha2wZDId9LLQWCjhvPgUxLEf7jrqXSjg7Ztu2JnGCiAAkDTOwXDvYpGeA7gXl
4lJE0IOdWj/iQBkAv0NYEje2exeSzhNFdriWhXI1kjXoGIKO0BxTTaNrLfWreLJ4zwMKWg37PWzh
I7BA99B8ZwGokpQ1nSflStP++MaZealw0zOzehet+QxFLwanE2+MNYQPY97rm3PLyebvmI3PYFkl
0uuHQdDEiU1ml1Ia1cXKiSmXlS71ZqBKmNy1/leIkpUD3HjpEkIdf55SMkho6dS5PoKqxAxsHZUo
miW8NR9mFF6fV3yzvDq8dCw/c0YDdesxU8E3EGZciWfosd/KGd0F/IbFKLag0U3WzHKXGHMJsCdb
uX+1oc0s2mnZOW6So+7TTsKbApaQ5nuuK0TdM9LKoNV19h7P9IL51sqJoNY/kUHJgABWvfnQzZ5C
PI/8eFB30gM88VSvSXwxz+hLGAxua6ZmyfiwIjEAPwB7eMw6/DepzypyHnNEsDMqhcCZ30Fa25OK
/O6F8zgwlH/TX0p8bn2/Pm9pDhL/MICL89ZY2Rl6nIWG7cQFQ79xR31GmzjrZw2R7MXK6dpHBCa5
vJZd5HrIIVhud5zXlftxmINTA/8DwffAiHT01Xt0A0HV8C3FuC6+RQQ8+eqeRgw3tTsEtvGAR+Oz
kNpWB08QJbkobzpf+Di+NmQ4p9rbgnFGysXeknezGxStLwkGlBb54n2EfJ9C/hvXJkMRUeKciWs8
QAsQankWLMnwHXHjwj3inbm5LGVaRPWAnxmfQw2K5NG6NVGuoj5m5aSmL/XKExrB7ANBboP2EPL3
Igo1z7wrE4C7zlSHgpXfSiWh040M+HiBCRxLbs6x5D9bCG6x6ND5rAmSTPRcQuYz1MLlzJTBhiYt
Cx1uWqyEnHQa35P4gSEPtr9lUqU8/oQH2xk5iQeRPT6JIvPg3sEfrbi0pxW/veUEHavI4V3pQ00r
q0+s+uYndeOpNUtOJ7pMseIvK+N3ddpE2ZlTwEICovFIb0WbKNlnZY/pkCBJu1XYSyPCgEIIjz7O
QV45U8pprmq3sO83q+lGNocZIuWhvR9ZpcQnxwaDJ5zw/5ieg10oPTrWLDNV8hLsG8qjpm3Ciu9B
ngQ844ncfQG8O23Mg9kE7JSLOB6LNsIbLQkJk6fysyg/dak73x3S3eOjdWs0aG+n9qI+pijD6hV7
p0ar8XSflTAvKesumGNs4tLlDjwbtQeTwukd/gHUGa2dcStlcv2QcAHjkSZtOhC+oOrsV1jwqPTg
B2bX0ijSEuPeAWE54JMYnwa7POsANJjVX6YKsXLWQm4Ob60gMYq5ovq1LbjWkq2S+YUGqTztgBXr
yA6pzfvRiqIXTb8XrvS6TU2Qwk4c0Lb2l+BvfATCSLzBFM2UwKew1BNP2ZzhNmZqKm7gEk1mqu3N
8q1qYRgvFJESA0/cvs7vMRkHKxraVTwIB/97+iWbphTn1bpKaw78STjuvSgRTl+Hpo0C1l8gPHDa
yhazorZL095qebQz8118nYkhl6RuhY5wxGcTMVxeVnmYO8xZB02W4VZG4nmDe5qf1s/B65vc0pw7
8zm+jDBn810NykXrTh7M+VpFSit2amCjsI3j8YkRaUGD1h6gu48qriCE2T7xPq45K0oIScuKOUzd
flNmbc0RRIT/aRuP9QFaUv6S62gYVTYpXWaYkUGBfvu93MHhROssdpQ/OSTbxjqOIcW/HF4FHeo3
iVQGk0oPoMAEi37HmfFVk0OC+XUNzr4sdstffQBxEhv+sszARcIrK1Ca7wYkWznqMdUs/iVWZJJ2
77lEmHwM6gG/mrUMQKsNJtx2hbJCzCTsmAmonuI5NPnSyzU2BoY0RnDS0Iiz/BXMlf+kZ0xKQkIU
7XtvirF7/gVNgl5BMWqmtARDUdsd4rZgylytJ2uW2x480ETwJny1y9oiy+SceNa/nn7zZVMLG34q
uHRAbjBCLHNTJ7cPBDCPya3CtdvS88VSxEaSWpzEaryvVoTEOSMD8m7mPsKzl7vQtCjE2z9ehjvZ
GlDxVeZwJLH5IyHL8tw+UyvYvnpTXxzcNbKNkGBZjSz5sxKQEmO/wQ1eACybusyB1MSPfxtxcXRd
nyKH3iVc4m4eEPZdnqFmhqVgsBttsSwg4nzPG8oNert1uNrUIVqWCq1FeeACjPjy9QvIJ/uzsxF5
NcxAq5ByYuOtqtwB5o8A+5jblFwW1q49Oth3asV84JsHwee1pgfiJzHc4iFPDSO36bjHuG3l2i7/
1eFL8uW1IdFK4ZGDmDsM5kayeRasWZJrWGbmmdDzGks5cW6vR7cS3tixrOtOz0aT0szb3P3VsI+k
UqbTgkYnbkushb1hV8xfhCGD6rtYc3UQZQ0GctO3Hx3AFqP6MAPx8PVE7Km5PMhwCdfYe5xhZhLJ
w0W9+NnxCboMVYmyqTm6uYlnk0Tf7M7Llf7F7BXLQmqc/TNIGc55y2R543k46+EWhkiXprM19yUW
7Zij3sE9eaAhDBMWtJqTaau3iSBZ4rZ9T7etWhkVnu6jzs/8sCOqvB/WFaErjZKDlDpwkABLvvEo
lo0s01pYDOYW6IDoZVFDc6oDsVkcp2H3YAAkJRaR8bacPPIITVClDR8oS2GBrWn2D+4hL5ASzeCc
oF9E4afHHD57jD/ES5znNrHnCfIBwG8Ur0MSTKmhz8qo/B5JoYTx7YKVA9Y9P9lwhiImo9erjrPN
k5DboKnbYWbHWJAMcOC4tBjLJlQ3M4dFF4yDPtecTM+zbqdpGl35WZB5meghUkHcw+v2xaUlrwW7
UyCeDNPNp/vc0XWwGr8IpBkXs2gucS0hYpie+9B48O47Kl2ZKmiorWfx6SLIAoY+cJmY/xrR767d
ULOXD3Et+84iQGHATDCqGV7ZtkfBQOEKhffm4CJ0j1Td9u+csrXxnrROGlPGbWM+1mejGeeaAq4O
/Xvdgs1+RjqskWAKvwwTtk3+oJgMTOCNMLbVlLqjj9z9tme4Gx5tsQDBC8SBcbfnsy3t2sm3Wecv
r9lwxLwe5DzDAe9KHpj5Xu34mvpEo2ZHPkB7XrwuFlU4TBK7mqfmg/FjMtIeqN4Q/Vcyxl/0Nub3
vjrUAmW5HSwXRGovOojUhiHgZcOJB8Koyl71gSqLS5XCvC4pYoHiHKJI2L6+2Sl2xPkRLk5lABiC
Vdgg7tvAJMQuzyqN8XCI/AAxtR/kA/iCUgsxzcrAuP0HZCRsT6nQ6qbzt/3mIL0F+mS8YtP1QqN8
4vPf7le1FbcpzsWflXkuHyisLCGyfLPjot2awKiOkOQrh5MhxbsJ94VHQaePqkwPh4rOu04MLMgh
R8Gko/maLL0noZ3yIGl9k2GZDs261afHp/CIaFLBFyVoXFF5cKuKeVPsgn8xMbZcKvLG1JPTs6zj
36V2lrScoIs8jrwduaN/juJ7Bc33PRenp6xKUtK3u6rIE78Ubm8sQqjWLhGavJqK1ctLTSZAuWQZ
18yuD2BDysyQEXNza3SIymwlTU9CJreZ+UyMTuFJ3/2QiEsJ6BRFUll7NSYLlfcZy8ecgZycxTib
FjZ5oFPEXFHXlapqKy+vSbFi/5RpEiuMtIWh/p+jjxpzJZwU1sl32pE43gD1iFjjfjlDxDJtmEU6
5zVZ2an/tV7f83W/BOWpCNSS+hxH3/4cZfCnXznIVndKqUFyZUBXBcG3BqzHVN2e43EaEEvKvoPk
xsjeHAAW15IIZiIoIZvOgsHj987p/RADLK+h3E+zkvi1Ct5tWhCu5L3qCpNLQ+6cD7f9RnfjpC1B
7RhSSdqh+TXQte8s2kydBvrik1p/iy6tdKJ2CHO4VYbfkCQoKGGuNWsVfO5B1jHBey29UrXKD0L3
kPmJQZSN91+p6Vlxh4hySqAU76bDo6iDc2k+L5nnFamyL+sEX9t7I4JvbTFibQNPHMh8RvH7BgxK
JQAikJT+IK3JSo/TQ8QsiP3h6NoRHlIIYWZkom3hNBLEy+ITh1MJ3zf3WqRj2D86m55JPFVukxwQ
anM3jMeRnpf9tqZSscHYB5f28CpTwIRNh4R3MrOcVz5vDZ41GpBkuZmKazHcjd5ILLqgLSAl+oEo
4PvfzhZZSlr7GKgBpkUCe1kL9/Aplk9ki8aioJ8i7ttIuOSAYqbOprtsHdWil7iXFQAC5iHqlFGH
eyDBeDyCZvN6o7zcq3rMerp+USbIdf3r8Ao3hiV9mBxQEjbBknZpsBRkuy87URMuMHUTAqA6r884
/mOB7u9EyGq5ckKJJYc3j05J5sjEzhQHzvGIJRCs9G57IJiHpF5Qe1I23LVM/dZLtY7v4YSphCK+
TL1Lc+wOZnlyT/JOG1A+m8N0s8jVj8jg7ZkMmLmyItkKjmZmlaXDwv7o8ISqQSD6eDIHqZ4xcshq
jd2vAcsdcrWN3wsh84mRpT/XBpPTK5hokRmTQxOgnx42RzmHmQrVEgdYsse0638VCD6YlRxqDEKn
kb9zE7TP+GwewW/M4pnanhIsElPYvTZXvoBzqx7HL6FLe8RGay5LNvRkxXQrJFXdX3zmq0P0S7SO
Imu3liBpBXFPc6yJis2tgAF8FB1g51u70+spBevpgwxeR7ReQ0fk/JBwGj+1hScMFM+kL4OIz3xf
S85qglP30mXpJ9LiPasVdMMNbeMhuJY/Yo3d0rUPUA8IeI2rNUXX9lW2TecE1aRhrd3siDBbKaKW
i223xFewt2bzVn1eIdLqezUwafWfUBE3a2TAqZqC16aOotEkgDyumu2eiN6/69c+a8zBhWOWZUB/
A90xbYS7Fjj0wuMjtgw3KXjBhFuDn+DFKo87Ruw37WKZP50fWDU84MSXvI+IIRb36yOZwkWKPhYm
5j7QL8v3zzL0vRmz7bVzu4eVEj5b5JoPOwmvJvLigtiL6Eu13Ja4QdS9LbasvTKj3dp/d2vi3+S2
+B7LLIyDxhf4hqV5SCf751e2wtThHZ/HZtZNFVvh3BIt4yGoiUL0Kj4kZj+syfDGjEBBYw1m+xNF
S8EtZUvbOvfZ/m5K1rbefJcrrlP13CB1FgryxLKOD/JQA7L23cbSd7wvNngmtxZRG85KbtomvNNq
fSP7o+MdR1EfIgCS3rHJS6z3nXQxOtdg8obJpJh1tpJmquHDdySFzG6ZC74XfFEKN7iSZYZwOD/9
W2Ml2rfM3RCbNbSDo52ZDsr4Tlh0qop+rAb2La/0sHjV3A21tHPkDkdDb0qXWHOBUH7tiyaRxu9h
fFkZEWdRWXWAcbEdJdQYJWEzsqbNYAetFgEauFOdn27hB2NFRbskBv3SqcyDAja/HxHuuZOmgP4q
J730Ml9leed2cYWGkcpHNSa/10RL3bqO2X5pAp1/No2ghC5RO3oGMBQiURe0+jb8t0hkqFb3LcsA
2Zj6MphV3wDAHzl1VG/W8eAqufZNVZlwc9pu48hRYF1SE+lWynxBw4XmHvHmSdmshVhaJMIQy+2E
sgbwx75XwJbM7PEOpySn5wRbXG+xQQAT2f8qz9o8VjgtZJCw98xjYWbBb16ZCUspkDz4jPU/jolh
4h12aV7bPYsPN8d/ohCUnMnKHZH4qgCiWDjOLib49R8tyrOjfU9/BK/zQX3uvgAPQrRbaOPu0wEO
CfUBkvI1Bvlq22cB9DV8Y9aZgxwxTa1xjGeX/AzMLQRUpitNqPQZfSdSrb4QhWXlXzQtPopIGWBg
ItFMCHfbmNEp8PaQ397dZXfFoXyNvjF6k8pIqovZ+14JBSunt1oXliijF72LPx+30pCGh/SP5+/Z
Fcw6YBS3nhRGpaNj1pZ2dBfaxVQT4osZv+2QYlzGOlKMDvJpk7Lfw/1sLLVKZIKbvd4EUbXhqopy
nFvC0Vedq2WM26UbxwHJDFT5WT7fVPLPBLMnqVW67EfCEQm3MiKgDwPb/pXXC6N+po+bV7+i4s9D
KmWhQBP8EFhpFbV2vMuO4//QWzxFZ3HFFKcgIkAM0PeJtJJrREpG4O7V/nPOiMgdOgoz+35DM3Ep
8Yfef/wiM63wuXMS02Oh23C1RU2H252hmdZ8JmutifbeEfWOdZF1SWIBrNzjPEqkDBPrvIdSzIcq
OVmtzrdkfxll8GxBg5pEjIzsjEPWW7YXcGwaFQKHX+wOMaz8lTufy8SzvgDotLirGAT+JZM+CiRy
ySuBMt1vZ0r62vKlMRNq7HT69HHlpa7YMchMrFHCrCIyvaC4gIbarJXLTOrBofOdr1JxLR547b27
IO5spP248CAKC7PpJ8NUW2FFOSORzQ3azEmsy0GfLkRroXNapL8ZVNBIroM3CxpOzxiXPdCSdwgt
tl9nRSGm9GjRo17TAu4FOuyNLS8u0NGvdKEl7vfLlCvu08h79f6QldzzxRFrkumC8C7EAVl52eET
TUx/UxS/rxe2d2wUjYTtQj72ri/bzsDJg07WIRG1wEz3rltidKJNMHj8/RLeWODx0beUz0+5uarm
aEVAPYYfktLgVy++70ogN2FSP88OD6kDpAFp1piRRExJXufw7RwQyGHpmrEFohAWz3EoEpG2sZ3z
tyIIvKhjW9F0H4isLilF+hOzPK1J16f3e2iF9O3qrQLvpfIVLDXp54cwGtfdXxqlkqpRDUZRazSV
jSoLyAIA2hiKqX8UVmgK2pHaFh7eHPdI+XaJ/5Rj/Cx69hMyrZmhl4qJqvRzqwCAIy/aF/w3NPwq
BbgCoLT9Jy25YJ/n9WaZmopLX4UhKkM4ywSr4P+nk/DJq/1ecAETWGgwkiyqCa9o1DgTe3iyyqCW
55f6FWSJpUB2XD5j3HhvGtcjI8/ZPgUIg+DE14KMvJdvcs+nxw+riGpgfB+sA02ltWCB1MJuI3PL
livuhNR5Nq+ezsopRWkpYp0nopRaOSIeOvrK1/Mne4Oc/TB8Yp3LeX73+RUtf5gY6ZW6q9XDq3Qi
g6PI/wqBCLqU+eepUFxsY8hlAgc0JX1Sr3Q7IAb9zNKllfKE+/m3J+3rMQ9Nk/SZXa2W46FSXGIj
Omynw25dbBq8f/xgqq3eCs0NL9M/eVDX7CF1QiYYKVIHDuqIfal4iXobUbn+wF4uC/ezFkAUoHdO
pUzQCi8J59LMMgrnjtqVm+uyIVPJUKdC/g8iYhixjPhfrX7s1wTVY2U3nzTHqhGVH+9HiIDi/zIo
NWGfkpuCeYkjX97AloPHQ4rbAdK4IFE2gxQviGXkGS3S2NqdUos+ONJ/KwgU1iY/lfmXrmjZxX+V
ZW9OV6cYXBDxaHq7ASUcI43YcPodJwBqGOIPX4JD3RC299s+KB2HkTBv7MWlEMX+RMtSMgNC1nGc
VzzyDZ6CZdvea8CiS5+WDGJVOjqJp8XjsT9gjgzmFENF6hHiGqUzTuWfbZM4347o8R6/sfdw77pF
jq+WfGpFExBN7PlfpwxtwwOPx7zvMqIlP8Faph6K6xAa/SC6xi5ChuuuCH1vcbNjs8gZIzEepDrs
tBjLBw2Hg932fXufu9pwCZg1FHncbGvn5ZsKYyk6LXd93ZJIAijYP93vpjF2eIWhkoqctLofaPII
F2nC3qGbF4w/gTFp21H8iPmnLWFd4lI23ZAVEb3Gekxy4hHvU45FsbOiUHknOovr3TaYFsdTEScQ
s9y2CoU6+zpsTcChe3RgObr2tbMQN+nVVkJSvFvr/5jSt3NtySADXkBq8m02mytxBBA1+i5Gp/5k
3dNH3heQk0U2KmZdQGbfIbT8rvL/Sk7nIACwW+2N/sYd/f7Uhqa/SpoLzYkxZYuDUO9svS7jjYaS
16uYO49QeEq8JefZNZh+447LBEQmvtFOXXTv6crTU1bqwbeBzDeaTmlOXBcJPb2YVWgjOECGrIiX
j9dsoNMjd3lUdy+D8k+DR9c2axCoYWRtCtI0kT6FiAfoF2uwrfYIg43Nx9eQNTRyv2sQYpNlr5qO
Pssi8agFAodvBCNQgNpFfwv25c0bnwX3MwGtMHYRv0VIGFnFQ9svw3+/s0gjzakMw0S6cSojH40f
jdrPwVW0IeuM2QuWCISD9aeIphsG09y9Dk59bkSH5Jf1XSi16bB6VejTtvOJtNS4+wngkx0DznRH
IMyuiQyvWHPMEyR5hcFvKuTSkyvvUkm5ySerhCGNNLL8hzSg/q9wxalaMGNGmiOE+a56vkHa4szm
SMQX9lw+RMSXFwqZcYKaO1kJqC5xxDrRJVzUc/+IuT1+O74jwjVEavvyN+ZLGEcT8WgKeSEtP1Ss
NakhtVFb30/07ICXHfc3eH5oWkJw9i868BruK6Ds2jgf76LVmkFqNkfRvPu32EqoIN95+lt930K/
RNP8g4UdF/J8jZSj7Iuzue2t6+B2U0EeKbTctuzSRbInbz1lPoIgvnku7OHWud9kjSIh2bFA3D/4
A8WHTLxRAhMuERyY19GbTWClhhwOJOzQPdT5a9NW7cIFfAPCkqA9BZNej3SaWJYVzTLtRRKW/ln0
npe5G0eDJifAJb0/Q5uST2MDnmVlhC+RuEwv1VR51SZDATstk/PYjbjT3VC2cxSWA+om6nW1BZuq
3v7xFDvV4d6syqydMmCVI6vz3I9LBWsEodowdv5WsSvWobzrhlnqzgu9HDWasUFearzpTtot1T8/
59cdzEpd8FZQLdYP/4n2uqM/BRA26fXkAmyUB+G67GmuIiDgN3tvuAs/C+K2oUwr8DFWuWpk70TV
ytMk4ahlQNymWuiF+0dKlA5rk3Qk34CJz2b8mYEixbisT5gCrCrvBn55YzbY1GhFe8OlEwrvhMs6
9OY9S9QZ+5BqZiJftZmHQ7SMNpNJRLPOqqGD1SeP5Txq1A1SD0zH72c3oqTcuiShm/UdAaftCh7Y
euBmSsFxvfvkHLhk0tuXbXq7M7Q9W5/74jNeG/yWxxSXA0pFr4RmPxQUKuBhnHKwEs2uEYTpHyrw
pqxnX08rSGNrh9rE4Mb3yTQlNiW7H34Kz601c67NSU8907RK/Mk1N9TCHvQB7HsXYcPdHZ4tYJm8
XJEccvaq92gipTyGSn3BFZbJ/zOH/8lEmnczZSqObLUNuedfC76Xx6bZu40nnk7d9h4pJ/gsLAwt
SFVt8SObC9q76lzky8l+Us6k8RTH1PZt2wElWi8zqI9ey2Q+SOLKpgegJFt88aR/gJyB2pxFtMnw
xKANU4YpE9j23jnYc/Rn8JEIBn92HNRSZHw/0EtoiqYBTR80WMLicRdm0aIkroVV6165YASAaJOI
e5dDntdyu9PsNrtLzNhsB3NFJlgX9qowBRX4ptLJ86wU2z9HooOGsx9/DhNhR4XuLfPN0n3wW62W
WPJDeNy0UB2ZNMdp1FdUFShQsDaJd7C9O0MU/+nJGX10BppVoj+GKVzm+lBpwoqMFk4+mdrGZ8ph
v0VKl4iE8TCapdNZZnKmIu7hTMBZSgMmXEiO18F/2RRFSb5cLJZ4KI21/L1+LkkSizPt5EwJ0ez8
DuGIguogDvZLB+tQrC1JMZOilr6GwHQm4S9dBGkgmHsefi0Wrm+qvgqrYfIJviH3st4PBd39BuQh
RA0pd74P8agx5sGfw8VSMgOCAmt72xqynmi7XyHfZx62LUzSJR+PBH2+DoJd41BWVzb3ogytCzpG
oKL9rXYuf97N4KYUxyVNpyvBX8rtnfUvHTySQRFbPbUomR2cCU8ayn4OqlPio0zn/qZjuwRf3+1b
/q4sCFPnU0saaKYW96jBjgmEj6htUaFJPKV+hsMa6QTsWuGXAppPZDFDHbSi3MUb0drMTZaSWIRy
XirFeE11CiJYayvIZybDHK+3Sht2thNwsSgUzJZwzxhTX9z/Zs8pwPrhnG+98NoZt5fZWriUB2vJ
dxviOzD/tP/JUXo6f+hRGEfIUo4pbdzP+KXHU+t2W0XEdOlq9DKx6pIuZWYBQJmCBl4HfrxX8K8s
BsIaCKPeObycFrb1Hvjzz5kXE4bmkW5blSEjYLyGGbnoPQgbz43PhnTnjh86Y5IsiC9tv5KFPTyY
z5RCCmLbhciMGs4F6Cv1KUshRRo19spLE+FHWe5aa3uXev2HTcXvdYQa8d/mx2KiC1Ofp4RUlxwY
7RmKcuWu96YxGEp4hRlfVcwq7Al0u4zBLkqMs25nB6xwQUIRXWrtPlFpYJeVssxdkNFbkaBGa+ng
e8aBmyXrR8D8QmdbkCudUadKmq3gPjY0yGI2I0RC/VCrvekLJN0XoTtOgE0CPxggK4OVM5/SfCby
W0R3hkqtnp10gZFqBp/xh5NidUE4PTYQjuDUgScDmhy2OUbbyW81Cy8WsqeZxLf8IWL0vQ8clRCG
ze+ka2jfBvAjM+eCdnroQ1U3Agc/2hDXeLjiMzrQnl/SHKJSsI7AcmCSYMLmp8jb2di5wJ3sylrf
au7bg0Je0XJbHsUumifrhopVMleyTMi92tuxTB7knXD3eGkHkR3PIMcGybxXQdHW2NVuhG23oF6o
X9cwScFs+Wr9AXnvTtGwH6lLUc8hhy8KeJiEn7jGtb0LcvbPNm9eLKXJHcBy2jSjQYVtU0y5P9B1
CPoXdLv2JevYv3uqMHqdH1wrfBuTVMqBl8wYsafVVsuAeS2g4ikenmACAnoeLUBUV/39UfZO8b+s
YBRgur91GTkdjUML5yLo8CbZZToPZjJ4DyIhckaCTlH11jI+A/99RgyFamdUR9f19hzqGK1H6Hu7
u4HnTTV54L+kfYxM2ynhUDQcQZO8jvkezAoLynCLWAku/rl47YjfG4uU75Yxbpf1EGS+eM23h9/x
6zkf1BQ4if9Ahs4T/Vkr9SvSdb7f7DSJ1DrhV9Rqp2Yn8DYoAsl+9BKA9ahNNKMYUsY3qJg/aIVA
S98Oq2Pp9eh/yAUq8wPOKj6KQ6KoWBrZl0q7ZKx2wmAs8fvZZHyux27bj71QJoLEHm40lrAqjv4y
klZGbrsK7O3GaMumFj0KSo8EDnOGPNdic2ftXBw3H5PrCdixuMWXvp6KNOm/7ysXg97Qdiiy/bji
Z2wDaTfrsiHBqhP3VYR4sIO6vICcwcZiU+AUFkVFbREn+s5d6Lz8KHS32y4gB96lDuBePyYPCQ2k
e/ObMGk2BMUHXNtmUQYdQtaxks9P54Wd7bOISeUxihnfkosTiABb1RSj1tgFajoshkTBjwftRpTt
P1KBs8Fyn96bAxgx41FaQvxoankLevaJ3O0ZgGhd3dj4iAxh1PsD6LaTHxAerFFQGvy4I/Vmd92x
0ACPpNIPrcIhYGu780wVSNho60CxkOj1uTb12U4C1X+fOUkBPiFQ/luGuRucbqxN3rbkRSsdOLp7
9a66JAiZJVwhAE15WLDMZLDNyCWiWz2d5F62Hez3NUuST2MrC1mrnkvM9tiz+I/QVe1dm8GOSCim
/QbLiI2kEsx4rpP299/AAl4qsw42l5sUBpjZTlGupg1jpBcz4OSEHUnIpW1hPKUn2g32GH6cyF3F
MhCJkAz6O8FYOm8tscbcnzg8lvy3x2S6bm/5hGC6q9vL7bu/iBlYa//FCFvzB80yXq6VU1eWp834
cMaYmJHVdZInhrHhlRkF23e80KKI9DKN0caeV+dJ6Zy0IV5Xp46osCYYu3l8OSoW3ahpNr/F7Df6
jcYNXBgxxvZLujgsWoB0lQ9ojseQq+BqSqFUreYWHYJVyZRpyIP0/HhEezXFzMk7mLGci5wgbXph
PtgsX9JlpHetWrR8TwvSco1Dmu6u5L7kQA3UBWFy9YeUglKCmomZOYpAq0lybFbxsdtseMFjq/pw
0HbvAqkmBagvqU/GUr/FeDVflxc8aXcViuQSsdnw2mx9YzKlqxPJA8LWnSSlg4+e557U00bXo6pC
kyZ8SGz1YKDAGyGfcy7WRMr0F6NQG36dZQVixzqJlq7UDbQFUFP6asOeSk6Ip2BmhqLRcEI6e5ks
PCWeMB5i3/aNIeOlODQFJaFPmu3h1fUwxMNC6tdb9ZehHqoBy04pSUWzBNV+oXQbzcAj7iBBny/k
nrad7VseN3e2ExLqEXf9LHaDsPpkHaxKnPzsk/rWKqD1SoGQeyQZihUyQ4NaunAW8Zlm9zLIzJRa
Y39EAzJ/29gKAOPiUsqbRQvdjZrx//+JUjUVpRQi1gv9c2fMrMNCQnptV33PoIpXtSriMfv8p9a2
LIkfeez+x++L/dQeHcMvl1muKNNuh05LYIBU2mbIq7PbvTWgRi4VyHb/1n2AcWUDWwPaI2MX1j8d
Po3x7z7y+vsRP519xqkySMWV/WzXOIhm1VlfFYzrzGIw/QhF+UaKeWqSIrnon5xHf1Ua1Td5kRJz
2xv8a3CMe+z4e6kZ5MP6uUu0ysYU90/MoWYaVEMsmDHS6LgmKmej1NqWerC9dqWlSloSzTe2i4Bz
7BO7YbVNunufVB+vsa03RbSiRum7IUzNKpo37xVFSu1RZmsR7eSh9vycPAK3huA2IPMLuHUZaTep
udkmxfWJFGHDoCIiZIfzSo8higqVSOuBIzbJsMqk/LEd/01GQSQrJI9cxT4kvHbHce7yTzawNNfb
+1HV+QLamez1sQTjcdY+Huotrf4jakx4VkXugpG8DkxOphiN573QAUv/30fmNaxKCk2rOakuyjsk
HpMsVrOKdkGC3AhmQljegm+ru3PvkaedEG3WsmnjuglevWAWs9tsVAXH94UPLF8CQaI1mbcCDy1q
kOHY8MVhcyHzH7flAuT71KNPIQn9pjEWExsjKthSFrpG0SHGPOwsuyEeRCHvEy/aSUcS8P3h34K2
1OOHF+VQqE9gCmyPNslEkwfvfzZUjnWAvd7HBc5yfWNcktX9265RyKv3Suyp4elPcOZ7UuLrbjXM
67xvmt9rSfDA5yqTCkA4vdJQ/WmalFsfFrHa0d1Rck4EDY83nsBAeWtpPi/1mictvtUN/5Dgfj9M
7gyRBP034aXxh3EU2BjTP89yKDrD7w9NvImfJV06mdinkGmkXjY131YsqqkMWepH9hHsX2zmGfAQ
nKOdCsnOCpiU9yEphRNK2scRZScGQFVdplsFYg1k7nUYHH7lR76nV8ZKygxXAv7abaAJqdLvfz6X
7422s0bDKdivSB+0qyZztUe/dRW722SVMIkdUWWjEPcvbU46Oytn4msJHGFgWuYaBR9GL3i2Z3vv
hLS1mOldOm2vKTo83IEzk4gnmz8vlOCUvsk5ULDNiMIoKU4mXQ4G2McHsXB1DIk0t/KmZz2ApHcL
vmP/x8lDhGDV5hrjrpEKowGvYlCRGeQZwckDlByTdlrA48wAEiyiwA3qvA0LBqqKc+GP6j5jLFa1
B9hPBeSe1FamH51qPywbjS3QI/jpywae4RMxMFoeKmPdhxdxp33hwhCZ7LrKmJkcpQReMTCe4PW6
QzGhmwe+EncfnXKMO7kQOJjQtOR+E41Nr2qKQ0QMDcRIp11U7PXw9iV91RR0D5b013eQyUDgG9bG
V/UGFMjtDDLrAI5E0y2R806WJaBSMLb2Iqcs+CI+ItxUeyhYx0iTFNVendwOpbi1fN1oxEegNIrW
DgxrItoC/Ehh+69/4PsPw4bjpRDGzN/x8RqCWYyFxiknQJoaxn7m4rIqaYi+R3nqqdcsBR7SQttA
FPf8UCJhCMONgj0xRGK3k7dHw8FkXOJ43foue79ArEwrXYnrs044i3i2rLaVI+RErb9lr5+UY+zy
4jbd4kA2zo1fJNwI6NvsIPwSxQGvH8Jg1hrUIfWUU7JNlVFIK+FcAgpKlWSagb+dRkW+wq7x0PZ/
pXpYS3ru3wROpHcr3B/j8lJQKMhlYuOqklLHWxaPa3sJCAAFBgBMc6GltKhJYoHR6xBCmb8GkTnF
sxZrQEyjCqXOEn29eNuC4jiN8g6CaRd3JqQKqIwiJZCZ8U2FfRZ/+auzbrLDvlEPC6ITUsLXJfMV
LQ8ctdJvWb9b3lf4rzO6mQXKgzJuJ8Zkw3lmSX8YNlf1hUwMmMHnBgyUDvXU/j4qJhp6MaEpVljw
tQMO8FBmik2RmwaivydSKZ7xy3Lge060gQKRa6dGRtd69q+p92pScebKXV25Gn6K9mqW6BLdnlvS
8Lxnu7XvXJbJWErJUCBFZPWj41iEOL8bd6gjDvljoPd2jx9NE2TkVSupzFjBz54rMjhM5nco2MsN
z2lM/n3dB4EmasOm4ZpoziqwGc7sZ1orc7SAbogoeTICUVg4LfuzlkFFoDyBq6xi83CIw5XuFZWL
p5PX+HkB6KTqn/R06cxBb93ecaT9MoKfNG1n30MTYbf8RKFHmKUgahgUmmigFzpLkpJVBbfR84CV
JssyyI8ETHKhHD1myzR58k33ssyWYvPqCdYKr+Cy2a6FBv+X6cPdxMGqgqMalC1sXk5s4t8drwfN
FDuD8UW3lFfXAyKTUpKzozIO9jpjmmXItPhZMOs+ZBxMmBr7/GQUwPBKA+AljlWPCcG0mjdweFcd
fQ4oaz1r8nFpn2pPUWrYEdLHAlacUefctpUSpq8mkIzki9MfUxOtRlGOGZ16YHVSZtyY0h7Uzjut
tHHXAUgkZfJeAJt65P1b4Av9k8MtnlGtoLoLJSSpHvOzJa79q5Q953X6IRrVOWZQvBwADrY5THo7
BiKItaSCVkNYrn4oVbT6uM6oXTTbcJVrh4IwWxOAAj2zQdmEyBNdwbTCDLMFVrKNPx+GqxQcEf6Y
XZbfqAanL0DmrtGGDAK4jz/aBEev/nUgyCCJO4hbMpFdE19GBG4PzR5e71MwSa4iDCxSQopE/uBy
sslXus8h21E5YC7jkyQzGPcIThamuYVnDE7mVVsYtXtj4zlcavnUouMfSEofp8tMEeaySmXpwrvm
92J4BLysT/nza3MyRjqz70Hb9iacGQOTQtbEjxuuNe8VhG+O8WNSEQ9Wk30KKcBitU/S7LW1exlX
fTFzFSi+kKMxC8gMlK8Cd18z3n5APZPiyaEgN89zsNBy88F23fenqDhEqw4W5lv5EMrLWvddrkIX
zFml2CBPeOJXTs+lIyTTpAax9EBlSh6T11BPEW01roCiDLNWTBonTjXtwSZdoTR8gcqS3p7/vhCW
3tf8AkihukFdMZKPzUy4BUyiJWBjKtVSogv+7pTQaVL6PQGMU445ks3urM5a6tKfTq+rsvNRPu0I
nd/vKlOa9TiH1omOdpApalSi/og+mwGqqIMENgbYk5uUXMCeHAopHicf4jZYVhzWQ3i/DD7f2HH3
RIu0z3nFqii+2NoG+JrktNe75lh2W0AmB+zcW6Jnm9VU7UVUJIC/WKjkpEyGy8dQbV1ZCR6it2OV
7/WOQP7D+5lsAAF0usAPfgHdTPHdGMnnbv+1QWpoV5q8yGzoi1zCUbuVE/CFz0UAQiprTzrlOxmF
MmM//IUU8X5BgKgaHEkD47V5B7q8eQrzM62GK7vjykXD2bL6SV2Q30qckUJtM04D4m5LvaH5cI5r
Uk49bviTMDNNIZIgrGdysmHCgFTizJ5mdXsG9bwxq1kxqhFhqE9Ch9+wmh4RS9R09K7e3CsaUF7+
2PIdGLq5qR6/0+MpOZYa4kjBBxKS8WyLGiohdQUoUW4VI/MFNVUbdfwqcc/zrMjWIRGDYH97EOlf
C1mezMelBEBx/r0KvbJtmLJ6H+m7YpDFdjsivdPEZuk/duKMnkswHF4NBWn4XR8V5z+mJQZTX4dS
wlAtbRYr58IJ1UyEzjiEuTXswDl4c13X8KKzhc/hdrvYO/4aSheKFTGrbwkvWrRcRXv+5MvK2LmH
wSbBfdQ1943Xar9fctnBBAL73jRh7nowzNRJaKPW2ZT4BsBJSgf43Bf20mpUXaV4VeNuHnSgzPwS
ti2xoTvExGoejLIbIPRHHa8sLpuelBOs0i3LvRSjK7C2RWzZX6RLtKJ4+EMv+rNtrxt10VNIxVvW
z8uYxBb1oFVN5umceeim8AfOc6/NZBAYT5LyiSdSGNR6+h5e4jCTazd96Km1w9696lbm9GW/Rzq1
kkxTvH3X75Y1JvnVXsYWjC0CSLiIBJaEZaS67a65U6AOZsAbivHVfjaUsz6kdST9HslpyNLKei2T
X46AqN0MbdsBly++jLjwbNbHBDA6tAaVCCXyJ0dz7e0AWRhPXGLrRkgkMorqqxA3iYNDJXxV6CCO
Xnpz1C3dSR/XyAPYegUdEth0Azmz6ACcnRT1pIhUS4I1RSAjFaozZuSxgEwMx571zQKCncl0fzI8
xUfUMT1VO5UZe0rKylM3Ur7cH3ryqWD8dPLbnxHS3R2anhnVXJ1U0Gdpyv9Rxf89KQoKv65pwO9Y
JRbztPgfflrpWnPTRUBXmWUL9L7yCOsb8Zufo/KF4iPcX2JqL1aafrmkR40G6F2kOtVWVFEPxXeR
/HMxaTbelKKCtjfih8c10yTR7pp7T+8vvdjjkdcB9+5SGDua76q9EF/dU0MoivqvleAIyhDgyEGF
BEb0AyqxTZIeTBqoMkaxnRVjtrbSQlVXtKItLK/HlfObEjiNaWjKpia5WgiC6nFQB3adoxfEl10h
E2LHA+Orgu+kUxLG0+FdX/LlRSJqejt7xzv1EAR+U/D28Jcz3l6MOStosrK6g8RNAsZq6fO1PwTK
nvIHrynZnhxsbYELqlm8TU4ztjiO+7hoKiCIKPFKmtVjggmRxl1MYKZQo4kc6zuOjCnBELhOLYBQ
IS1FEwBP77xcF9qwbbjbZLryrtZEUHbfyjwirUyikzMi9CFzYyATUWDKK7s+2myC/cXLyQtx532S
JN0b3pp3U+MszUk8/5+MBxYus0anO1qIZYNWa2aGyXcDNLXFA4I2gFkMr/fJF8/QhRF1VYmDlnZo
HIgi0SCQFd4mUUvfVffvRW+eYdSHaJKrbzzIABuZlWPB5651txugl7cBFu8DIAXwlvIMDn5Joh3q
eONqmV6ZyLGxkzcCK8lpk5fVcqdZlBP81GlBR57m7FJgnR3KG1GQr5faj015ajb8B6TPvrnr4GGy
bVsFryK3HQMYsOss3RvLXZuaRmZlzwY87DVTkRG7CsLWWzeDurQEr1HsADozBPYorclfSQv9lx+a
iawUHn8G2KIh1eTzijw0K6EIuBaCnvx+t+LHWdAbGSgat82MMBwbuNcNhGyFwP5GNoEASSfAQl+9
7axMCasnn/BFm1IPIWc5AI+ilXzEMb4+ktZ/b9AmMSFMmoDTuYLCQC+EoBLDjbtGAG+KFS36XDZo
J70fOi6+mZeNtFlz1DJJjVO00Ca+n9y73QpMllJP+F1z3JmCbjj7d1eHr7ekuDKd8HFcXkyaC9UL
C5sau8MZW2CgmEhibrGETk1S5GS0fk4R+qqYh8qKL2DmbPW3ehcXb9elV3h6Q/ZgPuv3OY+RoB9n
LfUqAU0wkaJQoXg4g81gqJk4lIGlUMd2LJPcuDH9KjbF1MAjKZdxDK/NxVwbH5fjXMzuvkQPUy9w
z/YNHCTaBrxm83QB4wgSayETC5oV/DbacRh3sCfQP5CTK4yOxW4gUN65Sd/YSr8+RD8LVjoC4hqy
gb/+De0seyzQuptkbDpTRqYLBMZJAYVg068/lUblQfiRjOtsQA4ZXKXfjGkryndB5ekaIve291JE
8j5n7nvzI9PFkZ1eKO7FoeANzN7VyIHjbOoiWbcofYXqMHGV3Gx9my81NtuuxSRBuOEaPaC9vQqu
932qh8UL0vej/ohbx6ojsek3LkQz+ikpR8zwmGWw2boC9eREqBO35ndSFejugjYvApjzWwo2Y8Yc
iyuMXDwL15GxNMNQIwZCijZXP7hyN2wzo1OHauxH0zYK/Nmc3ehuiQM6O/QHjLii5m31/rrybXa9
dP/FOZfoAm9I4WgjfbL7X4oPw54cbwvD4JIhiDE/mNwog9zNz3FXL7rlsT2E2FQHXB8ml7GvxK0c
M4nStlJqV2+4EA3y09HHVy4cXzN+Jhy9UHb5VMbEMhvAaMhs00euuCNYoTOK+25P3v16fmVwgvCT
9GtEtIaDPlHfE3p7Xg8e76+5p6AuIWF8mov8eeojB8zPcN4Af7JhvTQ6MUUMv8nMCL7VmXrwgI3h
f6wr6Av9uH7EAlhFNSdDPM8CEr3VmoPE+ofQtAS9Txfy2GZW3ixc+EPvL6QNcoo2FoKgfMg4dG4u
J5nWJMM7CSFEQozKCCpcmXG7/n611w0BRJC/71cQevTXegJJ6SoqUbrhQunyWKUsZKOQvYURfHee
Rp0fVxR6hkVUmtpG6P41QsUEVPyvAsJM2b5wrG+lfKE5wdUi9uc/8VcqVLrmzreUHmOafqPXH15F
/h3QJ9ikyi4g2/+Xq2/XKEK9ZS4MpsjNyVEJYZMdbHz02MUgondy9SKKT9U8DsjnwWhEBP9VtoHm
GoQafHMlZryrzek51nJ55iah4OI2AvmCKqNF/8DT1LddQxmfV1m3EU8LRbBg/wYHt9bUnP629/mh
9c5nVrOQ01LDq6qbD4Z0+IyrMWTyyo6IKldrWODQX21wtI3XUJSd5uHwky0IGrX3rzQfi+2ma1bJ
6x+eOUOu9ld226ZH7kF0NmGpbLgUXRu0T4xgER6aBpqCRAVKFqchgQ6sjsaLOUSbhDekZy9WsXRB
vrwEQl1plhcHQ/s5XTAdSHzALPP1jWg58JKvzUu2SeCLk+pRfPIukSDCesymJh49qVEzFZVYrEZ6
R9PwuDCM6P9T1ur9enLyAgrMqzj3RAxyGPeRuUPKCDoDB7EL8PQZx3CFomg191nk/H1m8iBPwTmb
abNVA5bZKaFigosuXp7LBPIF9f2oLmsqbTSpVlmyzJiguhTZFhbuJ6TJi0rr/AjMgw8/OzWw8hzS
tYZMt0fJKrqlYGLkRwdIoBtrV4fTe09zqHBJStwzeSJJmCtxDjhFjbQdb5hoad4LHrahukhrPLEj
yD8+q64iwR5l0YNMefluirKEKZW3X5ge4Rs2i0d0mIZZcfN5ii/OKqiuQwwv4jNiZwv8OUrcad7L
bkoC05Bc+3Iz73o1PhKQ2TabB6aq5QPyvKoa7WhqiL/KlFO0RUoNWozElShoFmUb01b6fY/GqZrb
cP+wERRvIu55Ce6Iq0+wIu2VZ5Lu2QcIqU7wYlEpF9IcdyC4ZJT1C7soY9TtWR79PLLRYw70onLx
5nxpAck6aNOSXcbRm0y2HoShPIBAzGxymCkd9zSflguw4MQJhPnqXnjz4W5ngmsrelp/L4GutCxS
BGFW8A9A6VrOfayjp5ZEZuGnI5BJTi302m6VNdNOJHZre/9BUbyutw8RzYZOvG0kRb3yD1NTuTnG
RhUUG6XJmgsnvsc9N4xnWNe+iPQ5z8p/wVCYyMByjfCRaicTukR24M8Jk8+MdowikHFZl+SBhUJv
/n9+TvzCKOHw3DLSAOT9D2+TTfzRr0xOzV0ScmF20TqSzkotzgbLcrdwp0Io6zovNAXrL+kDSDSR
W0uiwOuGNnBw33a2L0RLO67+L5m8mcm6vY50ZD0CuZVfo1iqVEg4fcXNFKE7AxI3lyATHxmQgEUG
uYA9UtZZX2NkhcSKy8AOi4DOUXFjkj7+I2S+qRnDpYf/kET2D4tK35ObVrfrZj+4up3dvwChEHUq
Gd1xcHQtrt6C8kw+0tKvCmfMcBS6PmXgx0lvnz67wgu8LUSr46p9BSVqmqx3tdNYVtdwxbVMZ7rG
JlLc605KgxTh8Yh/TgNlLsC36RR9Px5WVFpUmlDCS831ppNYiAFrsPbta3MCUysW20r1WCYiEL8k
27yNwA09WYZPaPMgwGxwiD8riKPwTI/bf+1ChDcQoEbDpHOS/ayR/kPyDVCgiwmzR53cfFHiVx6H
ZC0VX0x29KtlCJQ+dSH/lIhS960YTsnIpieCPexOwRyBZxTTMYC91oGb/1nfOvrQEH2rv23e5GjK
nEg4YUQuYFoPuuoWaI5+4DAvHoe/NtF66dafGXjvLDNdkXvqbwhGlIT88+M0EbhKXEC1ppOKPwWh
FI3f3+1MHC+noi0F32bDVweYJRvcN5tp24oXJteWodtY/cdbK1Xi/f262+YCGT7ifnlMCOpesxKu
LjTPayiwvJTx7gHMa6JLyleeo/go3/Vx4v47JRuAMh1fwgY2qTSwZuYX9DhipC63XKDhrVLdiI2I
GgaD4UPPqnhKHeHYEDJ3UqZQSnVBU9kg/RsObJeAzBX2VkD7TuSdVAkuV3gfyhBZGjMFsDKRYi1h
e1xwBLuaNM+cxZlzdpOVN5A9k66j26Mo3sXZi1MMdIzdECv+Md7tKeSsUHaPM7WBjKfhTifGHK6V
int1/CNXAQ8hcYPaxYKxaGXZBKdPbE6L6G+r6mD/FAlODnrFdWZxJkjVPH3gSkBTpaxXDUWbL50n
nKH+OHNELm0eAF4qFO27GvLFY/B7WughS3h+QK4Eql2A6qYES363jpm4ap/TxoGQZytvpOZmERMl
BI1SrsooSIPIEoVp14MuGnoBjsUhxxcgHhHpn8gtEmQKujX7uBEerleFqQ2o/4Z1/CKBxFg/QyqU
Wr3C2dOZZUwmM3Rh1fwSkhis35Qxt8Ru+xkULjTdiBOZHshnawbNgeRaL76ZJMuVhnrM99z9aNBi
zNUUs1O65VeaXkscGeOS/jMxGrYhKwDC/MWnZgI1oJ3z/et8gNBn7VeI+Pna+oi09LKOWoqq3Li0
VXowLwzGZ/DjfXRw61qp8pAs0873GfRshx6hAiltBXKX/yg7DZcJDPU5I/v34L/JaBPiSX0CWmHQ
FjwDNQeGH5d0OGoltTI+qFmxjFNEaZ8mE2pr3nrhQJEC7v7aotIoYC+/M/hDmgoMl2EWfY3Dlp5c
9brYd8I1HppbFA7UC97SwsykCYZlPNrdcbS79w6h091F/vOUs4L18JyE0CV0CJR62gsEJDdBoSfD
O47bnMvMs6YJLKEV/DZqKR/R0LzMQCzxtQvUVe+Y9AdNxxQWritb5UmTJg7+IRiHHzKHSUdoQiSu
YAGQ5NuoRWBoBjzDQVK0x568MwZjjPGzDuLpeCglK/hqKWNRz8Kd5gdlah5VqUqWyt7wViTMAROQ
f70uEZhhCKG/xyFNm1Hkc+hL5SkebQtpgPpHqnwSxZMq6wrvpr+pcnDsFjp4r4AtKM/xRDGuoUXL
WHEN3GYqfb92xwarKT7OUiQO40ugBOvwXWeM0V7tZEZKlG5g8gtsXoRZZFHtvP30HZyvn8VEqWDS
HSJ4aeKuakimdZuc1GzvCOyb1aGD3gl/N3eWNI4APsh2Tnzd9w6N+aCZIeW9v7atOhdueQIAcG4A
2stw2dBUNcDBr7/E4Dh/Q3+6BfojhL608CktkfHZOi2EEv4l7k21OuiawcUVYV9HFxloz7rNd46p
XKk0peEpvoWt7/NTuBgZjhPBIafgl3IaRe4p/S2HjBq2OnQlJqs8XOSsxA6NlNsSkLXqKTOYE3pQ
ysDD2JUwHyvHmBp/2iuKAG5dcFOCFspbdaa/HggLc3QZ3g3rodFOhjNE7wVkVrzU18FtUdH29sfR
gcjQn8iWSRpsnEaeUnYidbbnfAXhyu/tr5QnN4ONbrudsojNthpmIWJ5thZGgejNZLaRJ9b6P9lY
JURIOYJUs/qQIKTM0dWvpYA0kTRAyvD1Llc2eu8q/hUgdFTDAuTcp2tka28Wg5Xm/Ar3ExG8UAeG
bRkRWyHsWHRUUEfvm7wlDC44uj8J3cnwu9Ay7Fzw7E1FExkd7lZ5onyjxbwl/LHxDmb7CR81/7jv
i5bP92ngzBnYJM92uFKfVWymfoutM5ZSPieGhssKZ54K5aFbEEYqVBxjWdDw9MSuXqmU+ehl930G
R/4iGmkNwoFW4KG3AwA0rnD6s4IJ7DB0Ah6asVvVqLV5jJ4MhGISLEdBvfK8ogldS8SDCQ4o0UyW
6JN2hJc/XY4B7gWA6B7yGU0NUZRWEiuXqzpHAPUk6R3AcUPV9/dXtBws29ClTnenCuyFTwZ7EuhK
OWwXiPlmCqkzTehaKrbu4SePC4pmu5rmNbKMYxPX22y/DkaEjg5+3ClyJrHe8rc7U33WUki0CJOl
FxGXuxu1RvpBxWFA9DayK6+QKm+Ofa13AwsRscG1zrkSRahoOTqzNXMealB6P+DKRL9fESK+HHg9
xBFArkelLi2SxXbKuQTJXcZPFhJkMNW96EY5lKU/IzdDmq7uFMyBL08MBW6bzbcqS2K2s4CvXqOa
prgEs1PRNFyzHBFnwO6lT71pGSnyrvUf/u3+VKRGRq6e7SSurRckzbP0W1E0CWwpajJxGAd/cMO6
l/4t4fbBu+NVpfMBSuw46teSowrSRn2jETNIN41RGkMVkUVULsgth0vHWJTB3d/1mFUFvDSLyH5c
MnReOwsMGyIBGLW0T1ztQn5InZzt8W1UIzGbMdBhjveNSF/x0guMXSOqnGFe+x6lKaXnQ3+FhzD8
m+9e3SHEchM9/s0sZ64AtNKXs+ZARPmJzTwuMU1g0w/MibNnsQSmAz7uGQnYjjo90LSHMVKtX+dN
n8eocQ9aOVLLXN29J+LR0edYhn689ebLmNaCjke7jd+kiVtaM85AimHFEshuwZ9Wclhxo+U3Iiet
Cv1iYCZCUzKLzrxonG9WLWxxRHH4yf8zdCEIxMfn3AADIGQC57gxJO0/ER/mP5GEOCrvcy9eTQTa
OMNMjAB7hYFCiLVP60dwIEUUmzNlGDNa325GwZoYTGVhMlGBEIsYAt8CkyRYdZ45ZLnU6Xo2Aigh
XdnP6JHdN/K953fheIbt2t2auahpRw1OpBsrCUnjzi67DRzKego/a+Bytn9Mez9l+i1q9Ejr36Jt
fhWskkWrdztxHakyE3SOLNaq1cv1JFs4ZaP4biNX59kRVDuhR7bVrDJbMabQA9jHXdpGrNAhFZM3
Uc7IBINGFeosPAKP9pEG7+ppdnwiXXXzkrWaSaQhZxycwI3vE4SyaeNc0O09OyHzxtBbr/qvYbUl
iZZmIBk0P1vwN50vLDBQ8hUA2N+mHeJZ7ddze1cXW4+hph+EWTz6q/hE5ZSrmdyTWXudT58Y84dA
nfMtD5EZxEufbMS1qTsAx0TGzccDvv1drSQYwHnL3z36LcGRdexyYG0Bi6Hek5LYya5krGHHlQRN
ce1MW9Nr2Ft6TrnoAjUsO+3Jf3g5CUKYai6y0nQuQaXOCy5wpskfjDq2Q2MCwt22GhIVuZ2HqbiV
b3EHtunxqY2aNQFXmrcwElAkKNXVdmCGJkXMaNp8t98sfnXdxgEKyfT+UWA++IStgGn9YafepNsX
zNv9C42jxbkNIpHfLIIIyJhrDT8rFWVG71Hk1TRadZL7XggIdyklGnv6SqO3IkXopk7uxshUoXhT
cn6zveRrX+8RBSRCQ5NQeEMMmpGKvVNFxqH9FnObhESZTaLCcLfAvklDzzJb87hZh2eeRko2qroh
ECjIZRp/9ZJ59LbftU1f3A+RtefixGGmUBeFdYgysAqB8/dcJH4Tp6WpKxjBCc61aIIIFc0bP8Mn
kud4PExVXw61k0GMPk9MnBNON0t4SbMHfh3JxZbHVGEkDWChv3C7t6tFVPceRhGzrk9ohqoZ/gfj
e+UXLUS6tC2clsMbC76mGiOW+daYzfHFK9OZmxYteCJ11Do7QIcTiCYHQfLke0vZo8fKmMM4Nwho
/04MPQ64rpcqePRZGcpCOnJYOdd51/BOj5BagKK7ob4EvIq60oEyQqRFZ9y5k0WFE9NsEGaK1Xdb
hcxBoi6z45To/p2XiwxXtfSIB1f6JdM+ejDPwISc12gbSnqj/re5xk7oN9xIJSr+itconSWkncBR
ho16wYO/Qcrn0azHfGk8SkBTzTnnrtt/5h9aaWZsaNA8icUHCOiYBM3zuPNLnvMel4//j6o8tBjN
RsUGkt/AmeQeTvmQeGYrGPgAS2kS5DRC61Xt3jwJ7F8QgruLY1yqjHP+05A0dKoM0y7iFJb1fbJV
okIMUbOQpuRZ4b8vYg0VP93bkD6w+jKraFfBA3aB+lmUa4fE2plbYA79zvyNG1urIcv18Yd3M5kO
nRecQ7DUWPS7+DYlkIxIAN+C6NVQOA1J8b2+Rj0BoVcKmCqz0zbjvyRb0W5Hi+7NIHutUr+5k2G6
+x9L7UgPek0+RUOvi2DTJk8uAeTPGv29FHEdo83DOAlIoxwcfy8bLUZb6/70vRIzS2Od3Y+vE9EY
zhq6S5ZfetNMPazXCo4jRd3UpC3LC5sDRFKREbTh8cBeDRjP2H2mM3Kah2MfZgMa1ahooOAy7XZw
ALp4ymOipHce4GMPyzA/G1BDcbczDSuykoEkHyDfeRYKIdJkY9oUmk+pk2PHG1TZsR3lGI4r199l
EkuFZgI7jLRapgwWhOWyDKcMn7Y1mTgx/VlJiP9o1Q09nBn9BgX6YLVUm3YFmhNfKxfzWNyCYPpu
W7m1CZaFv1lIiNLnCHsd75dP6cxrDH3/q5RApJ61s6B116kUF+4marMRT+J6wJqbxKs1jffgFYpx
MGGIe7MrJ188hqxmP3LjqaQIzYPncG+oGC6x4mfEJTQcTWHrammDeJ6UEIWSmNlnOk1LIVwCrmKe
eHQ62XQEywMGWjqbOwYPwcdng6JWSIwDUAYxu4DkYnLDf+YJY8KnYFuOVvltNk2Cwnuh6MdLOEta
67yCZwsveDOkEaPCxhH2lyiyrdAxN5hNanBnltVcWFds1RJt0G0eagHpirXaHwy4xMEF5eIo0RU5
zLumzRcIbHRTW9s6lJjF+AkChsH0nFAniz8+AY27o30qteNBjHL79viEFxSR70ayp8lOxNmG2hIa
2EcxdsPlPhErsDVIBj4YTmsy2g0WG5byhVnxRM37M+xHlx6n9jgTrwZ7A8mXbNEkfJMkdDaR92ca
J7/uYAPwrrEdmyMnv1VNHtWUG7N/HupSiYQDGuKbk89gKhH1K/trSApRXQGuj8EEcOa/B2RzvpIf
uKqbcZNmJK0zd6j8zSh1CjW/fddRRogA4nOgl/lqltVffOiMjHIu77Oqb6pYi3h7QRJdtjNAe/DO
Bru93Yuh5xXnhAm85tCJimKn5ezZPlud6sS92elJ3HzYLyWSQvUPM9ZjRTLFRWblId/0W+cr/K4P
+a+Dnozq/l1WWG9r3J5ZmzsLUH8gWf8D2JIjikNaP3eyioT3ZLRL8NHXa5nnhRXgOxNIIZ8Ib9Bp
J88KzBkla2D6s/kGYY2/s0lbpbGak5rZs8aNpZtxCcJYs0FCKUJp3eulfiuYQ3zT87O5Mgq6C4/7
LoRtJpI75e7YAE+/vpEN3g6zBkYsEGauxgweC8MwEyByv54UPBgmpZtamWGkjVMB0jl3eu36JjNC
33WgwLFayLmM1lxmBaxtbi8pXM+6z46i7fbuUMf+seXoFXlAevSm1+9+5iR/8NFHQ+2XdafanO/Y
dBkLfInhrLdMgu82gDrAF5br++UlN8GMuhAUm2K+QymlHYAGpZPNtFWLSXhQL/9bqe3Zlh4+yeA5
BawVJhl/SGfTLYSdAH75earUyAj6CkWbElvKL2uyScIYsMB1cE6cg7gpk8hzM5a4wAZa5DTQx2wD
U8m3ADCNIdG6t34oTsc3tFBSqcgUyVZA/NjukuyLY4br4h038EmAB36KS2nyA8x2LJY7eI9G3BID
dZXb6Vl4u4l7RAcTL6B6zWs7ATcbrmsygYz3UgHOhmg3cU3ExsMhzki0POogh8rgXdqdTRmyttYU
hPen947bHRrR7yKUOQ3PqZZzWAtiHL4A/jWhS6VO1dspi3VshG/e8xeRH1Gw3verWQI/0Kg9K4ES
hUhquhgZ9/G7P846bFTX413sP5nC5tKJEgiIUUbsiNX/ORynTHJrrMCQtV+8/e5AoavaEs+YOeq1
ve42+EA8TFPuzwu0Hq3dLGPaqkd0k/vk9ljXr46sBkcO9fQJQcNvqu9w3kJMvVh7SHNlz/UZzZt1
SvoOfQ08l44gHPimTlrYBzT6WBGtumdltqeVbQtC/8ZmUZGO/r99uz+g76XP/EGGZeGjIH/taTZH
0PfxGofvj5W5TBqKKknWd57WaweGC6PrUj/9ZZcTvHBpWWBqC4Zj8GpLoojQhrXqFx8S7cCilDSn
8qjxyQHUXxk01RWsYxzaLfTQhEIlgoHSHzOoLJSqfrSI6ec2pv98tIuPYrYsnfVeg5YVgyzcG+6V
GivUJRqopwfUOXTKr0NciHWRJCEArdGLO5YtRUoSu9JEB0a9eK/fRqJk7kS/LJXmb24W60Sn1X3M
ZQ9FHQRqsUHlErIni2V28L+JHuzQTNLmc9mnZkABeAP3Xqz74LgiRGJ/wQD/egkHixWI4r0FXWDt
PihThrUJiLx/aLqf71XCH6LkZqBtrNQC8R+m1uL4vNDF4Y7iEnNA9aYLgJlyRacZukXFoI+imbtZ
ozd/u5kt5rx+GU5yx1piEJQ0V+dj1B85/GDeHGKeSqa8gSAhAGG8fGSaQ4SHzTyd8WF3LPbqAcIf
nqKtJRHGaXm7KB+o01vGFpIfnykoj9apLjeY441uJ2C6h4l+dWdWvZg71dT55R853V15HJZ3xYco
dBAew9Vx7uzyYE+rxc+ewnJ04Pw80ubukTs7fpVwqM5Q6Kgo2ewRoL0akWQJPzqBDswuCt0yvK0p
0HP2SNp0c2rZ9dLk9MtCqPGtlgocnA5U0d90RgYTGEwVfq8lmRQlSg0533QOfpy4lGqB4+ZCo1r8
lJZjqagF+YVfZscUZWacxh5EVJ/qmJ6Ln5PEWRO/C9XFjDzXOvES+F0AdXx7xilcsO4UPLBp2p22
RS5zBVlUku1tMgUWs6k+YS6VD15Uq7Nmkr1rbLTT9s9f+Rt2Ju5GPhIW30yVWKSzHhV7hYWaag36
URuLkEHFKl+sbkpiSSBrhCM1vrNOvPfJfqR0uP5Zj1e4BXE+xQASA6pNamm+bSY2r/gqgxTncMJL
baHGhd+dZioAwcfX94NfTP3rwtn1CDAMBoJpOXmVQelLNxFl5SQnQFGtFbYefV5ZRkF+p7dWD+PA
abo089HHsMMqD8y8ZLup6oauDoQXnKnmKWTdFFZu9xK3+NDQ07lyF2qDiOCpDSyQ2jTdVMpQnno4
gxCXdpn/BrfzcTziiOrPB2kCTTzjJPaGbsGNdD0a2KX5L9+wGMXzu8UQt/+cRKgF/M+WMZtA0uP5
bF/L2kx9QICVYPujgvu2swZQH65bTpWD0D5vu8yvXjY8eugdRBLJbnpZ17Uxh1nQ7JCTv74vm0Mt
5IoDL+4YrfUf/zv5FEVK2dZGreI19Uk1brl2vOb7UJci0ln3nLA/xHotk88rwHnp5YA9672nj1Ii
9FG2rHVBHbn0Rvys2Vt3gPlPkfyvt1jZirNatN14OYXSJg4ATI2tM/EEjSF3RaUdWHOoYy8h4QzK
sEnyoi+TSTOOKq/5SQuTq/aiYdchMc3Kqhu+G9vRMb3qVp67wBqslTaug+pp+8lGSGV25Rku1wmm
bqmcAMa0LqZooBUWLE6va4gE96ZvQpilRuw9/88XH/c1s7/B+L9gd2gGiWIW75adcsh0HFUrK7iB
TUSBsgcgraahxmsJJOXLm5C/BxQ+aObDdWiSVQXtz9sXpykXyKWnAkqJu7eHzyRN+eEmOtgkH1zX
VJ7Hh5TDNlBg1irBmCGlSbmmN4TjQL9Y6rFGNTO4lBQD3gySm02Id+TuhQmYrs893MdRERXf+puV
E/E0Q+TGkxXstayeAg1oTwj7cqUXnrIFylCez29E/Z0Z9I3hNRmAr/ZIR35Vyihj8C3WIa0kNvgs
xu2kiqO1Y3YAtrXlKGVenWQyfszqshMMjNY8XbDVrr+I5/ZvDA3MyAOhLGZQHgmL1lSHceboJJ8c
qFq4J9HcSaBU6Wbjodf6G1Jm6+T+UmR9EZnJixcqtNqpZto/rnTlrw+bExtWus2zqPEpbsOjS4bS
i4oSZPqVqKWzJEXU3PIrwjggfpHY6xqZBjauwX0Rguud2xw/ygLKVZZU3bCx+3dNEWQnqxXGUV7A
XYrrwA6ost6NqG1+eluaWMj89FNgNPoAMhhNiZLBbAitRrRp3pNQiT0C0MQfdQ0OzkYDj3cWLg/l
2mUHSgeW/fPP4FPFirylLeZpMHjWOdF/WYDjdjTUpjOfiRNtsG0oLy5+qerJOwF2ZPHFJzJyl0VZ
9XU+Q24QdlCIS3s3l4ndNcWBwCbrLl8j0VGeRjH782rbqa+rfB72bDQxMWmwaPkaDvN+MgDHNsEg
3A2VKowwJEe7H08aqX2byL7dfCu5rEbMpnDe3cH+t/xBgAk4QKES7WCcPDeDNbMwPn6734uWz4tV
+Mon4lISi8hqJQ4D4JQA67QnXtYBGoLdXy5ooCJ8drYWAv4goBQwWDAombqcwpyl8GJ45F+cXRP0
pwg69O2x/h3OHI+CzLsxQlqmAvdf8GKiaFIIiVBw1DSZTGskxIUXJ9CiAMz3p53Ey+HIVb+aKoX2
ijRWDn5t9aCJkyNj0uvmz2FEuxKpzHz4Z45gsagD4bxpai/1Lks5jpLigWrxjfyYO8JW7sedSvQN
6ehMq04GzNNJDT9g6COMeq90nzWdHJItfR3aVxxfS+MJq3Zou8ACVv3QkGdqD+9C7x3BiSG/LjlT
cVprwPwO+PkSIiEWBTRvLmhWKeTGLu72KKimJAdqIm+ELi/DaS6yJpSqGjW3tVpBy49wJujRw19/
alLnKD1LOFAy4qVC/zp4qEowSo/VTEEewLfB3peorkJ+7ar6z4atSP12+rx37kQ5zPebRiy/Im2b
MZyxVudknJ01dbMlDUFcOHyw33H652tR6an6a1DYU2E8yzdNsoAiQMbIUOVAuy0z9LBrWT/RL1cr
5304yxj0KmcHGehMb28euiUEwUq9sX1UlCALSR+vyf8RtJLogaN1HO8+v1+lPWGFaHMaSY7rEQvi
UvCaqljf1FbC95kKJD4vk41Ok5ZkqL671oV32EhSdWYoz2NdWAMjqE0XQRbdZsyvC/CqH99sh28P
OEEkDO9TApBwD+Krv+6zTIH54LPPLNpRDkZ5HruVonR0l8pC+XwERDQSx5vhB68ykhStY8vTcLbX
7ZoNsF1ndCZbGJzKQMdU0Q/pHpL2iogOPlCnToCSWGiC7CyQPOBNbHmbB210SxqBb4KAf7AWwniT
CyFGdjKcuBorbRxA3ZQMCq5+5Xm97PF1caM23PPyg2OcUMVj5vavNnaCsqtBjOiOQKKBOWyt/+t3
TE3yIfq+UUXol1ajBnIlsJUja6ALNM6sDSHKUqhYtmkvQRm8jm1nz99a2I9f7SgYL93E4mrL3A9w
I1tVPIQ4J4cxtoXQdbu0LPyzOhkPOl3t/QABDmqrYdNxeGy/IOXkhvNRHjTZ6wNCwKmiA5qG75kj
Zz0vi6SoDtM6ShkONmOytXi+jFTilT3ql1kCrXUQ6Am2T+GdEh+lz5RPAYLgnCVZEUII3v76DtvT
sxV0aJegscxFWT/ambH5HYF2crZOMAZhhmdCB4M6+vt/88hua0IKa/I/HeuBD/Kn3SUGM+1pGTDl
DEh2t4ii7z5PCK/coH2/6A/DQIAQxZPKr5n8UW8+jo9WNF11F4kTjXBIzPBlShPox0iMvHDNBzXw
eaJdZUECIgW1Y064f47LVLXsRZIXhLBllNudZOU2fJmXy7hMR1kS+40Pb9Wr1HgiBrWWe6W/yiPW
y0CmdkTOJ9xJMx6oo4nRjYC8gR8/JQ9fwVRKgpEaZ8IAjlKbLDbfYQwfH8lV708J+G3HmCJUgj76
YNJSWogxGeN9Bf9MLBgCMFNMlGM/qF5WJh+/2BkHdk42oJqz5cpSRlxqeolda86LKiZtDhB4ABnd
Sym/QHj9t8mmRGb5f2sJVsFl73xb6kAWIErNZhHv7VuU1pTL43U4zSqbxw/R67sJQhHDp3Ukwf+Z
GuGT8LhbDcqaXrGLMNQu09Vn76uoL3ekz5/TebnrMnflNttjbcbuQc+0dwaSLLpU9GWKLJIeQmjE
k9BTVDVCCytCBLb2aWmlQ4Ypu51uDnaZvTkpad09TxVxP3XReym3N+RCKHCbXBD9eb8vS9zDVG1+
i56Xfxchf2l0pmHcSA4Dx/YZPhBF/SEeCATkP798BGhVgiie5YyODlkyTyIqkozDGkDFSaAdzVod
SO77pKfdhGALxiCt3B9OUDSLFjvEQ3LKkFNKAxJt3D6wJtNnvB1bdSBNZrWZIVkvdJCFjYVwltgc
UZEW+mKa0/YcPZYBf8niPvNbLMwHnWI0kX7TeMzl0Vbu4kwigbsNN2JTaU3o1vSP9qEHAp/LdV6a
fjf3nwnSE21c+FumAHGLGB6q/UGjyJTfHPpcv2SWCN83eYHROwirwtsCsf9O2N7r9IVjuwy4kL7R
GLjH5V8sqCJpHAohQI7E4vrhZsG17bygAaSmPINMZ27QHHdnt/7EV681obag84qGJAjkOBtX1LB2
kymfmUk/fxUj6xUN5OJgUmMMghnfeoX8gekz8pK2aXwWVu9reskI1moDjuHY8GIVQ92Tx9+1579t
CWHDspY7Cd7ajsua+BlyelDDv1taZ1SLvS/9NroWgKnb3R8SM4b425pm00SO5POnaLxzqsB4tupv
iWZSQUOxwGLmrLlKng8O3VaybRcNnBBuBeX3iFn9HyzdYi8tg8DkF5Pdzic0hwFSXFmKY1pdwu7r
CedqzgXGwvEmiWQ1cdV4CuUPoPQoTzoLzhjUyqVrB/CrNNuSXbn+ojX1HiYBbma8iLGDEpu8KErT
Ldmv5dSm4p3VaRG4bKVveuP2KohryYKN8+heQ22F+reyB4EV/HQAZaK32EjDauuhtBOphcOlmL00
hGcDKPh5LY/yiqSEEdcc4FuGCqR8pIvHvwYXltsUZVrkPjB+GtHoADnafdIW/v5kSQHWBojbJATm
pMi/K4G4BSEW5CrXgGnTHVtBxkWDBy8ZNwX2iScMy+cZKieXrdnEdOKb2JTYsU8FlhJrsIiQW2mc
XTy1pqy0CWJl9L0Vp+YjTV6/fDf5meVkjvQehjArcAFpJcdrEiKB/By49VYYeo0xo7G61swd85Mv
27RUFtSPfYOUlhd6Z31xPK8ZbGQYavgPC+MQh2+uquDa6ldj3aQoirZ+Nnr8NXjvA4jVa6vB44VS
yWiJ6XdIRps+IRuP1Wkj290wmB6kUqp7Aic2DrsQvWKZMkjEU3PFzS5O7ulemRjtPTeJg++IeXNp
LYxgc7VI++Nfbp8kgWwBcs7wzKXy6v58XtqdLikBQdhkPh+97p/YBu8FWW9ncyq3B2KFZ84MN47T
oRkxnl8MX9t8JOrdJS9WdRL1bKlizGX1/QeGO5K2D4sMBALd5k9AOZwtR4PCtGHU5P1kcKb9lglV
Fmlg5MAteuaU9myEebUEoME+4AUUnXNBMwTsQyr7aJb+JcKJ8JjJqNcv2lYU6zN97JxMF8t4oYwJ
lHs4MqndEW28WFRT4yc/hiQbWKkf/awsgdCtx+aZJCsJ2q/Dvl42ceIaF4tyPlvsIfR4ELxn7SdI
dtgj8v+QQOw3On6xXn1iBiRuv0GLqJdB5QUaHDMUJi/R2ewe5XF887ENlJKuAqyWPmuwGlxz1EJe
9jgMIeofokM+xQAR+5nlSPbKHW6HN6nSbOVivl435/qtglt57f1wu3JqgfwSHiHDH+XitisafuJY
oedZpU+0yC+f3qZsxDgSY2B1n8uscejjGrL4HYeF77MmGQ8vcHukgnKR1T4WnElVIBhWDYG2tvCU
DOTnzM4vcTNiNtljQamWQgjrBS96mB0rhh9YIPQ9tel7qpbQHplQMZa6sZ91yrBUmkpDwg0PrrQ/
hZdBqDuNnZnUOfZAlvsXVVaWxmjWxaTOd+ehykpHE1/ML0pEUHZua4WagALopyZYEUOEm+w8aic4
SuLgcUIwRELqiHjp4wwkgjXKTdOiNX35N3VyKyqhXsEZLt68KjSb6xlxfE8BMkKS7axFU6Qr/S1P
/uVRpog+inTys2VD/M3Y/omH3FWK/cRv1EqEuL6wbLhlLLVZQvd+Cs0OJa7n/zDXiX/H5i/6wbSG
1Hb9FgTNfh5ZXk4Gp17g74VB8utZfx+mM/6zBmOImztOkqZmhd5F/FtW2NXM1AL59sS2YkjH0ZC4
U1Pdj3OlSMgOq+spBzUufZ6VkX5203Su/AGc3Na9rs+cRWJWEW19vJyfm2DZ2IBIxr/RnYX1X/WI
KksN6+Ze+8ylx90dRVB+Tci5u7vXvOyrUYHPcZ6tAehml74S6pG5U5xF79izSiBK9QZPk5uga3Nd
GpZi0830FoDnrHabhRallumYyBFGLZiETC2LcTR/Qp49IjIGdMBeL0iZW6jA1vIdmM/tXRra6Ey4
3ZV/hh9i+Pmgjm5FSYP4TB2hR9hhcfXSHLsYwIacUUDPkBvTO/iL2aXApzRMLMCPC62JF9umo1/j
kMIJpD2VV+aljAjQ2QeZwqxF2vOrI+xplOIMP0X4i6hVwJlMq6GE7hH6oXTjd+RTwCsoR/OQami8
qaXFhUKNjGNMJHfFdkzciB9sj+I0snxRq0krIkIVyn5Jl4DjTHz6xGnJ09b/Zo6qIfeQ8zv3Cq+Z
ncpb2uVFJJoKB40q8fipZJGY3Mq/DX/HtlJyNCiIjm3C5shqaIAUFwQmodzdlQRs8jGQmIkmcHPV
thiGKaG3vYdXI0qgCkTB8vGbUogUkAqz3f/iczuL20l51+EAIGDxYvC0INyBNxiglbP/vBkNUUuy
UYgvPqOM/4V4GLH+IeF5+WIzsBW6xC2FcxcgeoSClJrgbgnVFCsBkF2eYR+UekUv3uj5simY7KJ0
9dwMOv3pRHBFXtbY47D1UmGqvix21GBDH9fzhvTjVPLcdfoKL9iwCHlshTXgy/lpdin6SNFKLerJ
JfTA+7YdZnwhMIH22Pn5ki7ZxyKayuJhP/lxVxK8whleKwGNvANv9+R65E45/kQEytPqMZvgQkZE
SuIGPKPuThPX8vARjdLhd5UtDszyyTtqGnmVNM3aoVtuLD8G7F9wgO4b9WKYn6k27eMUH7WNH1ar
FxE5nGS5rD9jgvSIIuGfRgf6wp9aAItnqXbMAjxs9hdcLdbrL3sZsji4+G7YRqjd5wazh1ql+Ju8
TibtvEXfQe2t8JKSIA/qps7t0lDQST2KJdOY9hyklpT7Gm1ci0AsipMVcFKwiNE+bWico9jfuE7G
Eji8zib9lqf3dbBcQwzDEmuwPXM4TdpUHGjoQWj1ugy8mMERt3dE447AjQhHN8CDLM5rWk8BxWsh
wV1DxPlqYgyitu95mXENgs4kJzl5K2HMqsZfaRMSPRX6MqFf3nIoN/PGNqXKPNeMzg8gZ/eOmJb1
BaIPNJX7jzsyzuTLZK04WanbqVjU5ndhN5P1TG1hV0sYmDXGQ3HFwcHqVtxhi2YOfKJzTtw2SzSK
eQdF75takINUUz9xTPxORcwy7yJySVr8idZ84ZtTyseYie7g9LfHbGnvttUGoeIhFqR8du2wT8bE
5vUTpvmDiY1s483DOsEwzBD/MDMoNy0sxuhAKcCA4NDwAsWXJTfTbyOimitibDNVS9owE6N0cvxf
RFChvnLxDzkyuQ6sRxoiE22PDc9kTIYp4TxlGu+jdtBjlMab/IxHY/xXvyTEmfc6UqiZnZP66/Qh
pMCC1hRoY+qCUig30deujBpqtHbm2GsS2ijqycR9Ik6UO8jkdtLttCQAP80Ottz4nC1mXLhTMKV7
+5LzqvqPdbrJbKMhRG6VmqNMcyvs8QyGUlsxm8FvJNJCAo1AC0tOgh6JFY2D+Zrmw6thA0J9J8Ob
H1ZfALmI4kEd2CdNLar93tciagmeag03FmaQ1i0iI9aBjdiZ1hrg0PvyEQZpYdBaYlwDXVLPNHxg
Xlq3xLNIm8SqlkFU4DtzTBePzfvAs6aoRjV22AhBIP4mpeavp4aJ35W8oWpo9/9UxcwqrrvAt5JM
l6JJrGuDJORKcmKG+TaUQs866Tg2veKZPKEndm866QAZgR17P3cbZtdtpNjMwsUP0NF16wyRxw8u
kuVAOM/yCnI3kJVTcs8WTGrv5CpJT+RE/2yVzGEHBV1C2GoQUyT/edYW//KZR9ynnnoGeoyVNp18
/lBGiLuadzXFRE2pC6BTWCv46Wxdv6ty9wXTWAD+QW72Ug3/+bNTV/bS1ElZJFJlLaF6jOyp2DR5
jWIxQ1DBpxtslKfvIyPmas7Wi1wWX4fnCBrGsTtxwnunu18ZhnjQEdV/6E+3iWB7ClUE3iRW5esI
zV6bKP0d1sFUBT9Y/tTVbfokvZWsx/1vKOKPP3+tNGaD6z6aon9Xon/RFeJ5Vx1rEXMUcq6FId6m
vPEpq2MTtrsvSQvXgQfNrR/4x3jak7JhnMjjg7hFIQM2uOSIqz4hj5EwCbgGrDifq6O2aAL3dRfx
BJL8d9beC1LnK+7S7ax4DhoN3BlZaJw9RogcfHyEyRY7hT3c12PMsM8kHVMVGYRaGsSZItUDKRNr
jj9dncxuW+9LBawyrolfX8Zvf3xGFvnkmilFsSF5peRudB619gY/oRpQxxaeTnI3juVBf+Erdf88
O1Bm5ev/P23uZ3n8xLDAAHVT8QKcZ7XM+WzPkD2mXeIPAbqxSD5BjgYFQYyS4HY+yBi4TEpBDknt
Dqh1bDd5T/qlDT92XfnA6W9QPZOqK3wFtJrCoRgCM+r/Tbm8GJklmZqDyyO2rJ3V4UHTxHWWYI0f
Nmvwc6I79JUnV57MI7c9u2YIDMlh5GFw2nVbVLmRQ3bjlP+Z7QWF9Sc6jWR3koUUvSsFI7Ny71zo
GNOpE61ZWIJWZyPxpJIrNgctLO9r82fhFTp6yymTy3LBgFOyLuNxeblCZpfGpBsfG17/R6SCQgzc
TdjwrrQm/4xI9tp+luQmjnsKJPENh0ZipLX48Rq7qoksHI5Ex2qvzWUpyB0zURz6ySbWJNvJCy9E
1YIwv+CIpjNzmIUu9ZGIanz7/hsXc1nDpW1061z8MKWE2ORtXpcukfBHocCpTNwdX71zJyclk9Xz
5EaYk12BdfDdhaIvbnTr621OB5ACdweUQoA/HTu4a0io+qtk37VQkHaEbBRFAf1OSsidNd+TfXAB
G5gTS92zTwn7X+/dalyCvxFx/NGmfR/0Smyc1tB5jMWcjz4nhhB+3zOFoLbFI5i0k1xyVtVywxCu
nwaBzjxka1ZgU9T7xRzj2V5JQqAFm3DGEWHGFWzlbd3Q2b0FhfueniryGxwzPHFZS6gKIaG2w5G8
utgG1C0aKbfMvQa4HTfktteruhvlkYiFdpx/pCEjV0Cp81ua2VWZ0XP7Kq7N7HBY9qP7tlo1jjCL
9QQM3cqVHwt18FyIqzGKiHtUBTjedrb2pgUnLaq3fT9OK4zB0/QaVZNj1156XMfLNDLIvSqaLsY+
8c1Jiq6Lpa9fPEQKaFZLb1pYv6t4O2gpSGmGoZsDMaNoWRMyIwfxxbKGAl4gTx6BQr1gpb/w8AWN
qpJtBirHbRtg7M6O0XtvLzANWKVeUCAkYsEcbw3TGdzepqhH2Ao4VVWzsMl3haehJMhebCaqqTHH
kj/szx0VykdTu9DzW8rL9s4LOkAAlOgj2IGlDzRJgRsUvvfJKGlrKyHfLCTFc/DFD5WuiFvFJnSa
EiHWBcKUvelcvh0HKO7xR9LmImp2inTEBTPhKtuX+rMdx3A7u9nijWdHLRpHc54mSB76ani+12Ha
k6Gto/6xUbxpAlHf/6OPg5Skq4kH1eveYaRW5ql/cg2zet2X8Vtx3Sd06m6JETZG1tj7sXWQVTbr
TsWkgWZ17CDtYriewxG6x92MzxgQv6hU/H9fE447oDh8m6B/ztIDOskIwRtLw/1x0V4kcQoePuKO
eZz59jjXiJX3jUFVmiLVEa9peVH+ZbOGTlcFR/vkmkhGlRk/X963+aKo7TMS+HVOQ46ICnXKVbmF
J/arGiRSxtO8H+1WNCbk2gTQQh6rYFjSG+/en7kPkJoRybE6G1kk4gOkBX5qw9C/lLvbEeijBapB
R1HlAWOC7/m1m0gmjDIT5sTSN6XiPdwDrzS1PcLPoGqpIJt7WnIGyL2t0bi+vvqqkJOj/kFmWDo0
PswTnEsKOp3uy4odG72aUsLlTgsaBSvcW+kcx2kZUEoCjrLOOp3Th5wHwz6X36NXZVtAg9gKK6hi
t6tzy7fu5uIIpiMyCx1Jx8gYkMAEacWsptTu09fPgleQmesszuBa0s/VUwUKMTdbDivafXPqxhB0
lONxxo9g9qGWP9pqwtVJItETBcXBMkd6SOFqX6LQIB0lakU1MwA0zs7sxZYYYOjEtLMYF+Q5wLXd
9PyOn9ekDwDhQpX8cCAaV6X0CpAzp/IZH5F2tUt96U/VGb26Ta+k4fMmqHS4lFTHMrx20m6B1X0n
Lz4jWqnmjEkvNoNLbLh5eYnXyKS04QaiyghTVkeTiEb8aZ4uhAP1JtvFhZ9oinS2VKYxNaQqIivu
p62/BZuSr9eaELId39Fpfd0w2HCZq6JdkgHN2RwFRdjf+WV8OfHgRsTHedrcQ+d2v4sYzAyVTxEj
D0q3ehckTfcnxawPn16QajRXuHut2ueHjFzzpo5ZIJM/jkzrvt54xmQoknFiSr/t85w6S7WnM1mG
m54pxPWZKMJtb4fiIW5v9TX9/SttwGxuvVbeKhOVE1TwYgiVXt+Qjg+qijbaSagZuz1AZ97DD7mL
m0H9myIV0wpDxII4TpJEVxd9SyHbNlFbbmLhyDSnq/n44Tgu+u+6n5HU83j2Wg1LV39eU0jMbujc
GpxS4zPEydGu/TljMG6Hud6pO8hc+eOncHjtLugxiDWksv5Qu9jvIAPlrIwQO2k3ESBXwlnJG192
dTGviggR85jJlhpzyFtGVtWoYCqL9Nfp9s8nYjsjUpRKvjHKn8rQSuYyvYMss4o0rXX6ZMXUQK9d
GQqDMx4glwmvEFsment5B/QVqD+qC1LtQWOnwnuP/OmIlpFsNp4kVkKoWqLorQdZsFAVV/lw2GgJ
4YpByZ9fJPMbXBeTuCZounLuEmhrIUVfLyYsAodQ0lYTuieeGrsl1khy1pKhXHq9uiXJQQA06/4R
mkKv/whuY4PzT6VKdNNFh6QOsWmZzBZDLv2Yn5v9coismtRiU/6kYQ9BoruWUXwvmPnGg8oUPf+i
VfRdyxhxwd+uqLuq94vbTD5UU1D+9JR396zWs5C33jwCHK8rm0OivDanl+O5s0EgInBL3Whh2Z6Z
EEnQLN4qXWfDONtmzjks6Ecf9+IU/XUjmzD1i9fMyPGPncUYi+Ov0obP6Icax7RJa2/YfKOwF9cf
7gyBh96viYeanbDLLQNxGMM3aowuaQ7X2iejJZUTO+hHeQPm/8dBfwImWjCFhX/QG5neO0rdDH+q
yLmy4Ot2D0fp2zpU6SvpzoOUje3HAK8FQ4+J0zMHG0uLqSs7EAYWlR8k5OYl1sVyV+a6l2Bw5+XI
FgWQpwrINXqjxyXoIsfqY+ExHAhc63rfCTPpF808cjaxH/HzkYlzbeDqPpUYuT4WuiZ90TZE39bS
FdnYAGW6fYZ40wH8B2HSgNwVuYAo++G7zaD8DxWdXQHOPoVSXp2f0iZYe1cXScwuYrF0Ec+WG2+g
FiQk5sUnBxEqOPEf/XFgedpma92Kjh9PGk0xBVUzUlX0czkyC1HeNrZJKEAWeQD68aFwPukQDo5q
2YE8BlQ6UikGhR7nTxCojWUlTzd+YuVy8WCdRAugKcPT3H9cGVk7nB33j4mhOGAA2UZzSdiiK/yq
GBEk8shFEDbUxMJ4F5hs3O+Gsoosw7S6yS9HmCqNiOrWI5K507uFQqkD/ZEdbK+mszqoPjERrMXS
klCwpXjaK10dDx/EQXcvaUkmUIX8KBCsXmH/P4LPas4hh7P7sNdPGPhtnbcDcVfIwgLcH84LpyDO
meB+xyjYURtt0wKJ4JQsT8U1O0JKJOlWkEQm1EG2NHZGbsjBZ+fgwmG79rQfDxCHFgwCW+NcL1Zo
JA4ubfC8RGsOUgiZxqCUAIc/Mg06Calm0zpquVFi0x/pjdVUOmIxnXJfweBn2RQcZDWjqydYkMUX
St9BVL9QIaaHZF+tGBZBFqc+V0ODlJ6bn7D2Qj5Rriz4a0k7l/rB18/BkXJ3mDHZ6rFitK7gS6Cf
L9RwkiJbpneb+cjsyILKFJjBgu3bn0DbhtPhpgpi7lVNXFb844NUy3h7FNM8GeHmRdQKa7OvzrfA
tRfxUVmMAwzuBoMn9pJ/4uiNU+kR1rcsyQUgnslbB+g1WU9Tgqwhz5POuqVWzH4JRwYxDk6Bpbg5
noM7CkDpvoPV4V+/13fcBmUeE7wERtvGa+NikW1dOlV8bxau8AW5sNajvg4RUhFh3lmhhMAsYxpx
gZ/094zzQTmxKSOwxBoTdUEGEJ2zgtBztX3Qp8Yzi458Pasc1w7y0/vfOI1HZ4IQniI2FLSq+S5L
EoXnL+qADeJWzcXa9cYnOJZw62N7w0YpB/VeWp/PUMTF7lkTCl+99SVD2UDfkr5dWULCTmdoh5OB
A8b1NAdH27lZ1TxSctPJWGWMvUB0rPc7gIJZ+ogsHuALaBbeBbHcnThuQHE9MCjFaYDXsx3KwZfR
QjEy2F+czpq13UPtG0fWnfDx/H6nlpU39q/8JT7e17gX4U2++487VS7Rb3DM5rDBZYf6d5LRykGf
bYEImtFMpDm9+g8D5kBguHLw2xofWwso5yianT0rbWF1M6cVeXHYEPJkdFi31SUsgcjTYrRzguvC
1+DgxV1JHUYkz7p1ugCvGNJOTUCyG/CbL5JYugVsu2y8jZA6BcjOrLkIOYvFEbQs4Uv6dv8EjUi9
aQ6eLu99ipFOz9WXyw20QehyKBV3z+aCqwkzRCvHr+9b8m3pJJOvbsRtJ37kSecEeBI1U3QwTy6o
5OYX7VGoUAg8+tq/APfsRo0N8qzL+nJdOAV7CcREo3Z+KhxAULVIS7qAeCP5USjLKJ4OXdrvHAha
hoVPh8RRespcDL/creVP6TcIlExhgaGx6cKaWEaOB8aH2TIM7zG3+wLHnMdPYmDUWsJVWlzN9zSU
6M2hDuD1Ngq8tk87IV8xmD40stmJvpnH/PtrD9JqxH3Zp2csGRHqtAIRFCCU02voKG1iVKRNWQ1G
rMDaYdHpvfXRY9xeqigdKAygx/fiJolO9Wa1ha189qbZu3N/YhQm7NFI/Ge7uywBTgEHHrV0RCqJ
wznTNFnfXdxAMKoEX6Rq0Sh4u9W3RB/FwHsclsJI3T1my8PMA5KGjfyfpXG5NJjM75Usc5JLM4MH
69b8x4CP8kl96o24B8EaxfGldsQLbsHMklImqYUFR96JUZC12PXo+shL6gcqZg0ubEuGR9lC48r6
xHRCZnx3UwH/Meg0Ly3A6Em+F6kJcFodtRXCLxlxDpGyMBr+c1gxEU7gfEgzBx15IR/hPGKBZiOH
nhnxPM9qxyybnH+6Xa3dML6xTubAn3u9xX8M/Oal0G5Xyowv06NuuNAhszVsi3SF8uyS17BulR83
9ZgJrG00B3M1usmZTMSEEx0xO80qOCiTNEdR9iGgZW2b9ez620Nds4/Fzqhna9kZKWBFxDHcwSj3
7byBlCEKVL1tYaaQ83A+0qFH0PBFhqr5dhMhJGaZmtS+Kz+NY97jnsJPO4E6I8RRZ9Vax/mqWs6Y
xfDylYGCvMQ18e5rY74ddjJAjb20hFlMxJpojDwA10MkXbvr6EpcukSws/UWcf/BDoo8zqd3/qDK
BDlhEMx5bx6f9u0UWDir0fCE/HxZNZAsVb4V1u5bpeTIXNgC9WjV3Omo2pyIiwAoEJ8Y17rO9pm8
drckV2vbw6xeA4vLtEGqvCDeWl82E4+Bj1S90FoFMXaF1ijb6corddoaQ93IbS2JGbf4euMSTF/x
2sfPoGuTzhrmME0SeCbFCkMChATQp0i9XThuFWneeh2BziMWedW9VVLWJuC6q4DhbtLOi718k0Xt
dwrvkXktf2Zufg+k5eHrsrtaQ+k7ksZG4nTxg5bOi/cqyo4CdaXUgLK+UoBb7CSm9jZRrHgxgqps
/5Zy36OIiaTro+3lV7A0q1X/vd5OvHdJHAEpGToG4zshQgXDVgtSfpBMJgZvFQ2zNvBsM1XpO2qC
Q9BpuXh5PCu+oql+cQdwS2a8yATZY6bAiteRhu3Kn196kylBYTSYZMah4YSe9Hc4SWWOkto+AjNN
dzxEz6YrY+sLK+2UqOOC7ONG9pKKle5uyyeej/6O9jRhnI1wBP0bkBBdefuRwEE5NQjHhulvwFhR
q4EJ1+P4BzaY1wgdtGv8W/4dxCip/bdY0gFUKxLnvDGLjui0TgdAKu88nQ8JfLWWE2MjAWeqG1iY
/fzBro+vdUJsLJegwjgcu+YC+mX8G8H3kDQtXbtghKw+MBwqA62ClexF+j9dK7ATpvHb8dW5RWUM
/9PHC5yuoi/xow9/SckiLkhi6x3uyTLQThTQveq9DiDy3sZWq0DXni7fp1l6ZODcSPV3D6uHXLie
K8FbycdqnQCuzKHpWAta2sr5ciyv2ucmpe0myJxbwpiGe79vlG8JuMqtM3tbh7ihtjyiUw78+slq
eCwCoAw9JENrnsTsiWc3miXvnp3YR1AKr2QgrW+iwF0TipFtHDeeb18zTIwcdxcjW4kAwBuprdd3
RIpvJ/axT2psMJ9ULRpYA7U9fivvRc6cbS0fK9EJRBXgMRHFK1bhm0M9ojt/DIxEYrdL6jrgRZYQ
5ClgPb4PH3O8NSAaw1teCPntXWPDxWPs/c8XuMwvjVglsjWk8BgT5Von9tcyIFGJ7B7GvDWlOuzO
HkzQB3GRSFQMPd8phfggMNVecIeoS7vMSOf2t/u0cfL7SoPiMi7AAc/mDAm8Hh5uDzdAZEVblWNB
Q0dGLUCZxeBx+VEXEkPrycmfA/NRgto50P4nPvBwytTvSx+Hh4vSxEDGAbl491n8JQY9OUW5RC/z
VJ+XluzLnaLevP31rw4Q6qenzTN5KPRRKrwYGoTykaDpLP1loWP1v0JReQvDb82ia4aSuUZtP8p6
nsX7ih7vieizeGbOvg+dUMvtkDcxbUCFQ4o7ZGayc6x0j0edxBvzG8u9R0B0MmHtLhDvC4St2g/b
HEfiVIxudE/aYPRdjqOHA+1AlfUwnzDICwME1EySLk8a0l+4m58xYRQZInN8B0nOLpht83UEFPr8
iwRWDIkKpN72LAs5HW9fIYN5ivN9oCf2Au1rbanDxMrRPrLzyDZ8OJjArEche/VoZIkNMkL9mP80
aqdlQSftddyPUUn58qHUtKo7dubcvamA5/97kWjFaUl5O5tLl17yFQgdHvapo0f1RaOf+z3AJn5e
PyYtlqGrW4TA24ulfyRpei7edvALXtCOiWvFl6TVztLZfaOVdwlmSr9Y42J127m3bAQpj69Jous8
iFClwvKuYuX4xwhdkF64q209dfHTcyXkFiryuvzyV2W38AA23ww5mBvI7IpqQ5xXJIkP45KoQ95G
fHK3S7a6ZazCpvoPsrxeGHYtiIrdgf9Zo7se1IdD1KZcbHa/YPRvqbpJLf29Z5C451WraKvOwXeB
XHuuYunKufQMXVmM8fkuQEU111ZyEN+ld0nHFMnofEJIw915LMDC25bbny5Qp2no9jSbttxZC4Yj
wDeuy02SItTr5zBAjE8o4/FaC6w6BuWpZolczDHqqagmv01hvFktKBqR9QaQxWtFvrCZmmXx8rLN
g1dPGXPnnlhSA7W1XWlJCThPT4+wGjHg19XbIoRKV/PlfdxNDH/WEhCHJnx9iIyb1UvRIwwR2HOi
Fp/H41aFQpe+IAvDTK4o7SUp3a9jr9NeEpa3CoZMl3dYpJ1nQe5SO9BwTiuVFbf/opuO2biF5uld
Sv+0C/TxdsmAedX5IsYaM6gL8R9Vpfh3aSTOtzVHCjOzYFOf7/aL7Eb/ZFMixwlO05a+kMruq6CT
+d/pd2JEdtwzJgj5bN45nxRE3CaghQMAf+gqP3rcxcgUdtqca5sCqrpZJsiTRhUXu2pgPalyoMTn
tpNW9AUBx9sp/ekoi2QT5SGztwJ1VEHOv9fO//rYnN+pgdhwSuCLerqfcJ6JyH+oeg5ovOwYgX21
ZElKkBtpctWrToToRtXd8iNPAvZ+Eh8xz5Oi9/kxD2I0CGHLVqi5OYrVbt8DTNVOcVKltC+sI3DD
hCy9BG6cBFAQaMmrbxTHd3IBO7983UhsDWQ1IDb1ioHS3VrRq2JNOqtj8Hemcpn+I5ehrF2uCDI+
qSQnfmcxXMVRZ+kNxtvEmdweA0o+NJM1at2il+FLbszhguzymWA+t7nqj6bAVmQbnZ2Hwyyc/bPN
8bxF+FdcQiPwQtwQpqpyJKCUhP2CV0pA1Jb9bKOW2V1amAwjmZs0ovpb/SjQLv1UxlvB71Sd7yc2
vb8iqIbZXdHv+RTeoOvTldKhqRJJxEoZoZWbHjPPQQAKh9KxhMwg4vJ3bqwb6xrI7wwnQ6uDN2tI
yykz0Kf+QMShJogdTZApOUgILYi3M0RqCdKvO+92XHAp7gXXVYjnO0gVImVqCWZlWzUVBhN1Wmvz
ZyYpLA2C+MXgoVDA6x8PzJ7MRQeAHG69nbcbSGRmdmwl7jctp6NsDFnZzMMZa7lbVMPDTyYpMafh
cs3mewDa6gEKqi7IKuGjV/bvBzum/HxJlizeprfrgB4hLPmLPmueTOe+4tcxqoPPoxSXAVBRio0U
JXnXd6+d2MqUBY3OPrBe+VnhZGHm8U9gX1BVKAr/cjjTVTbC8ARGcPo5VaOg3B5TduA2J81qLBU7
YVZ/WNS6DA0F1LdbUPnpcHArVgRL5YVn2IH+of8fEREotw+jcdT634FnI+bBOfXkNdg12X1vM9cg
CMBs+HPF5Yen+sTCIW/2jDrU627ZQgOi7aaY2wBX36B/qpSX/KtdwZrEwwaPG4SGDY0ol0lYSHoy
XTzBzWLEYltpPKwCwcBYmHu+Mv/SdHcYk20+KxxIIPjkNCaaXO9N8G3g6aHQl3Us8MWwKj2NTd27
jm2yvwPmHY/jZq5NHSd5dzvZ8mjWPwE1t9SeYsDitvpOQLQVWlqI+AKC8zbt5MvrAA3FmlDSx8o2
kQYZ3kot4s0pzoHqMMCpsxPhqzeSXJp1pvcC+lm1oIxXz/nfFHMwoE+UgsLMkLXP/bh0iaGt8lKz
rlMHNXG60agKyxGbUAs4C0LbWFVLLAdoSRdCrMIbTe6NbkBNZf63W1X3uNnaWWrwD+nko44ZXW/Y
jeazS9W4mbvlFB7WeqsDXsBtlnDV9VnLQ5XY1JrB40huBIMlDCISzF6IvVByjqOVy6roujk1tNHb
tgLN8EchT9w6rmVlfx+MP7w2ABOgntIwoIzEu2qcXSaJ2PIV6EZw/tsOH5hdm3qxIphJyS5OmxIA
eMyGskgZUGhu1w2oEydLa6T2bEzLnfohW3NEOH1dhayEjjYo5rOVoXH6CqGJRAK5Gx7gR/OA6Iy+
fp/vwUeqkowUJjL2e2a5RJHKzGy4z9kg37CzlSyk66+H+GJEnskkcoywSwVaaH9Yrj8qjCOGYzvL
a+9eFLgURkh0D0s95mj9ULKqIb5+U2dR5LCgzX085dk08Xpp+YpwEtB+2uxkz6V8QD+mxmPG3c1U
Bdjnf2vhEZRGch393B6sK51KKfnMkftJqPUJUYT58TPkyUEUAOqq+45Lrh1qrymDATMTeZLw54Ng
bTPefeFjHUxoe8yuNhVu1THLxaoHVYro83K15VNt7IYvlofDLQHSpqWBq6D1TzvW+roi/Kq0tMXC
rjWWmvu05ClF/nxn3fKFDeC1fB+9Pyj1PWB8x4LFo8mFvwbFCCp/cq2dQj5TJ4oSWxazKdmQfeag
am3QEUG7lOVILmZiUKvz32b1vYyIDr2n4IfAzI6L0O3n6XkPeJFifBb/7K+rCyM+68NrsFmGdRkS
nO1sxNSpUWFVbfLS1XbbiDSFAbvV/KdrSylbgb0WKl82igZoPd0bdOxG7t93axPfCXho2UXmHOWF
tk6onTE9Y+y4RtjegWFgJuSJ+CdWCM7D1LZLw5j4NV4uRnIrggXenMc7aocq7HXA+7QYZIH5XZKf
pe5jiZJnX2gu4NcOVBfOXjp5H/q1f3X2VYpuGA1LZHbs3CPgTPvAYpNIM5D+FTIcyMd4j+/I6VW1
aQAHzRBT+lYCzh/HXAmrSKfFoBstARgMNxC1HzDMLY3jRt7p464J9ojJ+Uqfs+N0iTjCrb3EGmMn
Dtd9YkDQ3OqLm1KKCqIsZV33mITXqK4RGJyeezIwQWzWSvUGoTtp/EMEKwBCrKPzS6I1h22w9TKb
iwCMG59jvizVXxkbhV9byGLHHlMZfhPG7O1jXonh1sRVr354cmhE0KCu0UASkxiIZpgZtrybSrAK
1gX5V26CHMzxKNdiCoVCkl769SZbe/UdeqMhyFJKU355F/8t/70UYXGqtYSx+oQmAOEQBfwj5tlv
zRVKMDS9hdjc2yOVMNasjGuFr7XrF4it5dv1I5MPD91f3x5LmeAvjiDbLu4UY1AhCRqFHMX2tuu2
BlDCZEOrNmbxHyc1sGEDoEcn5I1UAbVRAGMnfTkRnoxAtcm23yf+iipYHMlbMumjlq4ANsZCxwmG
n4jhdpAPZNV2hzjg/R1ReIgGbWInDoFdcB3aVCTuhwfxH2rmvbeaHLMdgUIxbnyIW5u8U4wP+NLF
hRQztPCKaBSA1KNRzAPzHbWVvwjZKsXcVa56QQcxTTLNuV1fRXKn+1p6JwCThyr1MGyZkU8xltYv
rAWna4YxviLOyNaIqicuV+WfCjlAl2LhPUmHJj6xzm0reJqPi7XYgQkP/G+VCfPWlY3QhFiTixZH
KUZkUU2PkoeXG+vVnpdjt9EMs7SA/RNxKeK4ny27XEF1qmPvopgz4D1aorJ3B/sXHUwhGoOfHbZO
6Z5MOF4DFXE0tIM35QRX0d1DTrJg6MtD1S4h96YPobaH/63WhegH+2n/tnTy8U6k2YjYeApnLvLr
bLeZOSVi5jlgkyp6el+O5U0SEzzyaSZdwXuxoDfuJzs90DDEoNUbwfrsuTWnkLI609vPDQyP17Gp
hXa5FA5oxg17jBpyx99NOPfdaRhqFHNf3JTVZilRcXpMY7uq28JDwgGA+35WMFHZlIeGe5/wkszy
lez5SZNsWhO8aDOr5u0Ub7KWNOQ/dynKrlw1vi1GRbzUAskWcyNz8yLyMVBLsY3WXVkXz0BTkVQF
AdJTIkE6kAJEWjHKFcTch9Gp4BzDZITHq2AiDwoGN/85TTYoFijtMsINz+njUN0eGvwnm5kAMEPe
HnHQ4QR9lRaCkMYfRg0d2CE2guIkIhNRuNk2X1d/ddaKRKUUj4AV52c+aRVVwgGUoJqSsxOg4Kda
mA8mzo6CngJfnbnqiLBQCNQDTEE3cKBryKtmvPkodhIZfAjc7eUk6/OjDkXIW3KmRL8aCZYRVWG1
HLJRVhqgZMks6Dyng/loPhrYX4vl6GMViDY/LJRQSxv2SQ1uOkLZ8H5wT7MwsjPlXowAue1Wrl8q
seOWFcOSj+erXsCLk9gSakyo/BiOCiFPVN11i16FtBwqPS8FsXaAKt7j/rag+a3PvdQCmbAmAWd9
ncHLe7/m7gmooZ+FUFlKeUif5SystCojaKJHq3Ka3LZoH890ikRS+Sm59XgWJNn+TtKKCU+NoixO
htsqeVwHEqyL98vhsyAeTx1cpNSFgp06Sz/u7M+OaTTsC/tSJvlyQ1Ho6va7kdRqthiqKrr2BM4s
ILvjIngHCXTCUwZhUuzCFpz87OVKcxySoQAduYVVVaC3rvef18zzcNs0BeBC4BZaIWm2XkRgJeJt
wN3ItwxGJaU9lsc1uCLNko7R2rFIGnNpwsMz3+SDAyjyHocRjUpCGO+9qfrLM07rKS/sn5ALa9GY
VdEMVjDAYU6vPhkh5TQR0oOb4VXGxagFzcTfhJ1trh7hQJhP4zIwIHV1j7ko7VJSd13T9//Itmm0
FKqBtTa2J/caOkKQiHpotTH7DioG272KBQS1jp21uRFwd45VwK3KV7xiEcyjR88CGAtXlQGnIkXx
mqbX8igM6CCsPxrvX//NTSTxbPq+uimLbh7N/HwzxSn69wY7Ls+INKuEU81nGU06vgiAg7dDeiyW
rTjDF1DteinEB4Nu74AqlJqKL07Bs1AKXg3rB7mT7cV04aS8AnCcW3AslEXMM6AIb6HTQXUQe76h
O2o5gZARYZno97z+vt3VEbX2WLxla2gfql+5DJwybrkLOeW8kM90+kFowv+bTaql75lkkAKMXSaM
WSJ/CaFTDXSQ4Dd9z4XJ6pBKVMIBE3CWa9aSgh44Fei4xoFi3hvvqdFoObHBpbn14dCE9Zpgbzni
HZBr4ODhF1N9DE2YyOHCKXmTSPELze+0Lf1h8I5MD4GdEJMIyeRWMQ8KY/0CR+/77ualcbdeh9GG
oKeTGFoT8nXfLm+uorNClRzICY1CVuy0VRjlf42Hsx1FX0qvd8iiauL7Yy+nJLeO8LJj/jQ6dMDz
OEKZ93mf9YaCN6OLLWIqtZbGiEdhGJs39qcjLTkQJjDJY71rVAFG+Yh0UA5UTu02RV+fRNZwZg+X
vTi25oFZsqTHOGcLcc2Awj/hRnBD7VB92Q68zTb+0LIPJLUVfsc/F7EWuW0S7OmZNHMhLaCqs/Kd
OAad5rCsgO4IJLyl0Fua7nHCZaJ4lJNEAP0VfQP2mJQL3V6/1Tk5Z0ggChdZUvj4EJ7gdkxYxcw9
OdCGTyHaGusFhYT1lUkUCxIjSuXxkm49alQN7dAaHZL8SHc736x/uvHhrrKUP6bihEOB9PA0JIZH
zQvyj3DEQAuf/6E5Axa4fCETrm+LbFO2oy+1Q8GmvMFNNhn9I/oT3aLrswl8ay8KC0G0W5FprugC
rSaIORal43FRJRaiN2Xeve46DGS4TH2dUHM1ak7Goer7EVjVchVtjU+8lIHvCVVmFXgH/MqAz+rB
7dgIjbMWQIg9dCkS3fu28m16FzVDdyhx0GY+kNynyolhu9GVt6u36VeIGyimnhe/uXZB0TslIPKr
8hE25lvmeK5JPRp/qi2UXNep8GExNiVC2+1koQ+NCoUjN2oFCDafZX5+LjUUmrm79//jcjn3MEVp
zQB0XxjXULtxRggw33CqIcI+E3YGvmh70zpAQbjrTx32zJMf7h43HPxVOEjGFQnSVQaPOpBxm78g
yXTyzTanXgrmjsbn5/iHCZUQogPQroNaivHvFqWcm9SZhap8ObPyU2alTByXgL0X+yaL3UqbmAuM
HI+f+bOrI8zRmlt9rdzgNOvGRWGqWRzdNBU5uPHpqw91dQ00sG606+RErku95lxpmdIn0eYy37An
oiAdGzXSba5xyiWLX0rk37B8Uq2t/CEevINY5H3kIFTy7sMlzx3yoaFHDbXe+nXiwKXvDvuY2Ol5
DhuAaoHm51F7JM4sK1QBYKJNdZpSD2YET0DjsGwO9ntiuuxFsbBYsqoPYI5YHdV2SHaHN5s7tm0E
SRjQsdI1u4PAirOfMXg70Q4OOi5QJEDYgxXOY8MAjm8/r/tEjPfrZ0/TSiUuk5dVgJ3NW2K7XAte
roZHIZ9JfG7Y3Qc0BAtf5MotIwtcLMtFm4mWjREjjT9pzPXm3OyNj+n221yqYPhDXZg5QXlr28QD
eS4Jk0VVKIXQYMPXw/1I4U9MEJLII7DN3TwdiRgtg8B59XSedWAu73Wi84ImEWt2o2bKsu7p1LUs
wJFaiw9XlffVBImRQDwBBwIGD8FzJJqIZm8ay9sAjWwbUW/LDUFnWdzFDujtZ5mY1suhekCT58d4
p1eWoLTT6uvJ1x51ovy3bFkyQGrVwB3GkhU3tsrrQP9+tB+VZo080hFBPOGp0/q9BrBEzPtcXavj
c69l9jIaphCBO1tRY2+Z9jIFFwQ0cJHJBeF4g+UXc51blNsd9wHXVEDhohHOY9LT5cXlXvHvdMxe
wRJMX05iB1OlQcLlgOXuVrn7KbkdBGqy5NIBXrEscSRY9vjtOxCqO/mU118RjqTvdnQRtdqAd+Lq
V/3EYucslCP+OIHuXnfS48E38dtNI8S6j1R2H5SmsxLyQkp+Nn8pfb22v/meqEpUihMh+eNGauij
psmB01YijlvGTx2/WFQzg1LFgKyOHZOUIqvliGVqsV4cJqTRF1ECL3nIFlwF2HIoQJh8NLnj4H1A
RyBkOTEFQQ8rPnDZ88BmbVayZmHTfEOM6SkulHZIhMiuY4B86y4xFJ14p0gB8+aJXNk+IHMcau/X
qfptF8ytxwybV9HE9P3IwtWIMdXsk9iAUTIM/K1uXBYqzuIzy/I527qTLxP53XdLjGaXpFF3f0S+
Xg/kMKcm9HSX/jQZEqHyIN6yKJMIfOAj4XKRmgBD1KTEy/jRL+OigtSKnKeXwQyPtl9W9ci/uioX
9phIUoyH+cGO5Qg+FHkuZzjpL/mS9y5NzU2kDpQ/Mn5ptG4faAbLjT160qhIbtfP5AtdDjIYaIfp
zjZTZt9YXH3FBDP2x1oAwjw+pbLpc1Isdc1y0f6lDWWw9dX+dywltxi+HBRBQIv5Mdm0s4Va953k
Sfd4lQgYDWpqwzBD0o5FJsZxVTnpbiN+XUD5ZZaMsrdi6Lsvl6P1cw9/yrypZOJLaFxL69Vl26Bf
E+TfgPqMazr4kVG9PIyB84dgVAFP9oivkx0DuwBx1927IcbekoyksKNA7Yk6w+J8tCDWl+D9crMk
uycpTi4c15ktV9/G/9+X/U5yKN8FJuXXf13LAjcJiyj9JTa0VtG+F/5NdpLAYyOJC/5/NgMNOCI2
GAKLwlXcrmk5Hdr7rODAiqLSyYpOsZQ4Ip/TDf8G7Pyv9P/ckA+MDU+rh4Y2WS1Of+/hCRyqLniT
J5DwCNSPaLzb48IJcuOuLwB13tDO6nBabgSbxVCubMOh1CBpfkixTuhwgCPIzp7WGG0EFmgcUa/r
Terl835e0UjauCbTc0RfcJy93dWvPdz2HcJrFddtQxB90nGpMmVff4NY/k+qybdIVzBvhIo4Ofpw
wkoI+5FG23Itb/OLblid3uFhX8rAq1vhjVerABwMPdt0ATqUyRMeqU8SQZttRQy0Xd86lfJVbOVH
KT5EdD4+8SRonaNJPBMndvMYo/pF1oXirxnjc/X8KNGkL7lzrLaa4dTzGsGuzjBia0QHJ1i3gR5O
x8gWzxXGj/jbdK03+dQfNwg3Qedd2jfoclaJLcKVKAPHlNtYM/l9Zk996ptghSLtfgjt6LGLce6r
Mjabv1ln/RMsR/26mY3B8ebirb4qMeUYR3woDhBhXWZv27mYQvjNo/mDTq4CNzwsT5aD4ZjaXwKp
shURccKTdIT1rFjUAou1Mo7SaY/MbTgP1+J83Y+IX/+5FPSpnBs0WeSuDNrxT7Hd8ajD6n8WUv3u
ogaSa+0Jv7Q6/ajiqI0TIU/JlVIWX3deHTdtbeEhKssH9fHnZ5HL5i7Li84et2KkyaaXj+ZkF43N
5RR4cuLyprbRMKk7OvZOVrhqYSoBSqcQ13gGbOYx+y02aL/IbGE9qy1iAoVFllhYawUAtVORZNQJ
v2lLyq7vHq+yzd1jak7X47V0vQ9SChCOXPgYAcFK7yZ2pEzX+rOZc2WDSiSs0ZGeFgDAfZ3LHjIz
iwQaxsF/5nRLzpD5bNUmGm6UM8d/Sf71UTom0s7OtIpQ7KgApv+5mhsoaVrEnZBj3u1nZYDr/RvH
e3aCBbp/4YJwbuBSZg5fRAtH/we0oo8zAdb4FvtrCCd3mAj4L9qxuc7cyqqOiXV4T6dkhv+AWDSn
oqh54m4TuhUpYatIZsndNaoQ9tM/kpmC6H9V/m0EEtQRj0s8CwEvZpKYfazEWE2+xOG5b/4EkJvd
a5nUSYTCRhowvM93iq/bhWmNxJlOMAAXxBRlasqszwcZwRoaPE9nxn/Igbqm2bEle4c3ff6J4s/y
XxUIdE5grWFSJodMhH+t42PafaQ4GuAe9fuWZMErRe2a8zS7RiJt6UpZwuW8dQ8GhwA/BlLf+Ph0
tNy2Kyc/6S25ZMCEgaPAqrwzx5vVNyNTTxLpUV6QJqvTsCkMd5xg+jbwSj8DZCaspvuRnvJwNHen
tSw8WPt+3MGgO3sf0aDyEX/EiAK9aVHYmYBYyiBbc5Rdbmdjzjpv5AfEr1iYK+WnfS+XX1uvDYrS
CXYIxEnieX6QmwNmpOO5ExJXGFurfniBQl+yyyNtiqd+uks2Hkhwbw5NZDWwIlMdqMZEI/W9JpMZ
zn6c7sXgXKLHz48qLuK0SiDvfuRmOHWBNPOyyiAJY8ELJ50mGeq6tlpqDjSvmiHF4GKVUDF+R9b0
qWANIQdMixtF5WkOiJmu4erl+fWPrwsvungG7m29e+jIfT26itdGe2b82RysrRJQFtql9DDyYEqD
P3gC9abwrTLsbY/hidVJtoIhtbLqzz/WUv2YSfZ/FHJGhmfHv0OkDFoxSvllf5LD4WXrE8sOCDFU
YjWKnfP2hGaE0I7m5B/vyl76oZDdIe/dpsE+PauVDEBYd49rTpDwhJRNC5BR5w/Y6fNNXjBqfCiw
vW2GvrFPv5CcqhTv89Rk9ps+x69zQ/Ps+tXHUzaVsEhHch0xhSZZJPDa4f3UoGt908RLbmDxxQJi
8Sy3uQ315BA/UiflVWi0HUWeAWwJoLhfwbhTtJQtKm5RSpAdUk4aXBP1uZcCxVff0nCdA+tHkSie
C+0m8qpfPJLVijzVYqRLcYQweczvzzyLt2c35g+UvgAfQzxUnHu9M4xndrgFhXurKafh3Ja5fdJf
gRjVhuXwSWEMbgcJZd5Q0z0C3n0O3VY7yjkdmL9KrOO78A/vPAM/VEd61ZAehBGwK/a/iTOInOrW
Hnyn9nGTGqI01ovw12mkrokL7q03MLqWIehD0jLGI9eQ0tLeAOZn2iM28ihLski5bssVxcc7BkNO
L+0Ip8jrE/tn9rvExFKictCNLLOHVWXtSiPDpH74jsRNeqYVLMmptge1VhqJXHFOfj9LZJiLolHJ
8unwUmYbGu2vt21JpwkOTvDfOblArXIY4oJMYwp/YuNzp8b+ote/RR2JrpL6MDf9yJDqV9OvPmn/
PKl0MoebSoz2IFSd0yhSAysgdiE1WpQ8o21DI3f83VDDQR3/rm5JL4+83v1a63hH8vhmzUD/Lb5n
JwQedkIBfzzmlOpm78/ttwbNZoLrGYRq4LB6YUdyPkcklKENqMA7wncRoZtDlwBE22qTqaRtfix0
Z5OQ0qUr875FtPnJuXjA2sBEDZvtp0WuMwYFrCgIfEMV06s5jWAai21QwVCCSczMByRHHDkYCt4j
E2dqRbttVTf6vAEcYr/WLHKw2AsYrgSGN4Av1JUGkfvaX7XqXlpnd5sQEngir60lf0b/WcZmP6wu
gbj00DJQn/DUIWMmzh+IKTW2oIGADIq2bnY9AhbPgqODrCQEUMIQKJO/CR0tjbgibQuc8deTS4SR
rrpfi6VlfMUUYQv8/nlhz5uRuoxMH4aGfau8EruKBkCZgMDKZze5OmppWJAKvLHPgu4xnU/Ts35i
LZ6+XTo/CGNKpSqV+b9raX6o+d3P1oaC4wcGssUFpqgypGQVr4alBYCIIZ+bYOjjMNlckT7H3I/F
FDnt1d+CEURTlcEByeN8hxmZ8BZyr3J5S3GdoJSF1+0Ec5nHIBBh+ilnPyuv3taSwRPDKQ/2J/94
bAgm1uqHOSWD0389hyEF+e/gUXgSg1Hy5VJQ44W+DtN1aNsU82hBFbTYPbDvMfG8Ti2oABd0IhNR
69Xo6GFJYJEA/RExrlQjKCLBlxo8/0P+Ftfj5Igwec13AM2dcUHYqv4jNOgSJViEB75EbyQ3h2ON
Jscg3QwMmKfQ+5reF0PwmxOHYK2nvaPXshG9goXkDyZbZkGNActkqOriSKovZ7ztzOFaanVayV30
Rgjsar7Lfba1i4ILCj5P2qXDqoku0JuP48JKUvq1g0z9/gkpZUclmvA85LGxsmhn8OKISEh5EXrm
CsuWKjFfes3xC0HWtT1o7V+aEjjbW3Y447gAslJFm0bc0kjL1h2e8KwXIFZ6hn5AYHcV7QV5Dlnr
ZOindiVbmBAXi4OncZR9JecOcdgeZsLrB9QNtbFYKXwfVy6dZmi2S3g8fHoXQ+jDZTSkdQtyHau7
KnThABm12XEJSKXBp4oxf5JZ7WzNyMt3uNl+Rdg3/7VV/NarMUsmlTIfShHJdTuH/e0PwWu6V5la
XCKgEQ+oSwiGhNxf7F+EB3Nb9ZjyXYrLo6zLbhmrw79gXzyqytTvjHiEzQHA1/dGRPmJ3RHqmx0N
vuIwYmZ0gVmUGHro6KomOLTuTmF1UVK6Ja/TLPS8IhyGyeW5tR7rTH5l8VrIKHAiLHwiYdk3+hbX
JkBdlPxra15ap3jcZ7WopA5IhAb4fk+WtQD2NxzJam2x+eYJDbN0MHGR0MKbX6WgH+VHr+Rz+F74
rtjxl62K3bUg/Xpu7RpTiz81vp2PVIeh4uiMYqkxXH6aeo6s0Ok67DU0GVF+yJgP6UYOdP2bAUZw
gTioZHilOuNBPp7+Eiim8PaURuWMUAMa5ffTdMxnqi4rXno3kDjgPCcX37J/IeeZE1DrBeNosiw8
d0pvrntKcCZr01g/DfPnv1tjOBLys/LWZgCplyv5anYJ0FdAouVeeFyzNxotGdFTrYetz5JjEHYl
7DA1ehvkJ2wUgU+baM4Tm08gbSTWl8QnJi0KrJNIUhBwFmK6FWANw/iKYx46ZKCa2s+k7VRsmsoR
AjW2tOP8Oidd53kTrywUwc4SUOkveG3Ncuph4b6eprB4TFgEsgCU4QfcJ2Art7p/Vd3TbLYVHo4t
p+xrG2LYRcOMQFlzJbASReubFOODmFYB8fvWW00ofu2ufflxA9feYRGnZYwPUmPuQZBD71tM+dyB
hz2IBRQGQ1Vzy7pEgwEk9RoKUO5WjUL+4E9zUm5U+iUVOZaRaRChBUVZeHBIXmKnhQQPSxi5OC1O
tNtwNuhaxnvSAbgWKb56/GguzodvfDjoJ8jovAHdHUb9tgXn2LVcj/sbS0iC3k9im31ipGxqdFRz
V7s1KYkITyDIX9nNmWJU4Oe0O+bV0D5d+lGek0H5K8na0zdjSGzzCl2waZPAM6/JrKYW3AxEvFwk
My7YOol1T0cyemBujVcrSo2Jhat47B0HC9orEBG6SdXQP4HkjuLOWmL8/RZx2sbOH2kOYSu/tGzE
Cgzlmq6fpKo5hm2Ekm/butvWv4Wfd/eZUxVHAEHGsQIWN+t7bvm57GEIvb70fyrhX5UhAC3nM++K
B3/HyqkVluJo2VQnYl+RAOHXsyPVJq264rOZSmRnE8bBUSonq+eQ2T7EVL3EyBQ/ORBwl/FscA0O
DWAmXypER4iedHoezu05WeZ4dv53NXFt1xtssV0iJxft2dDVvV4Z81NNb93+iTAIaBIiGuApy/DF
MVz7dTS4fWUAq/LBgbaw14j+LZKhwMaQSekRMPVa5KTBshE5g5eBaip7QQUzg2TFTt42l8S7mf4U
HCCntDXQef/wHcwY+Cl57mq7VZHqYoaqlh/SI+ZGuhsJnbATAHKIsH40y5Jj23ZUL+jR73xS4aO3
nRa/kPh/Ix8JjbaPLzEpOCWMJ0QpS6xudaeIn4CluG+NNui0QQuEYuGI7ThdmvnKC9HapHlUKnbJ
SFcdbWHLJMbNwrUlfjhambx6a26YZzBBT1sakGnPRFldYx/CQ0J7yUuJ1eft87DwdpyIU8p0bbM+
4+5ACJfe1R4iddmgj3x52SxtkddepFetA4u3Ey7nnKYkzKeLHikW0WWWShmjIH/Gh+m4+WqvUM2e
pT2m8sCxKiZDUUXUU0SqT8DC62eo0dzCGH/mOMbYq5VJeYe7c68oaBsFIj3OiYecKZ/Uh1aeVSnj
vl4Yu2ZOUuODqowtALs9dse9ytL8C/P41lf9c8K2vbOiURQIDfSVWZHJTV6UvLdRrjk1L3olKsR/
jqgFIFNLVOW0za87sXuzqLxzktaQZfKbXiAokLjpGzTydp+8DvGulDFMmYRj7vPmr842od1+rOmm
hGSUl0VHNSN8HpsAunkQ7zVuKJuaE0qR1/JyQgxPb+EIFJfj1WddHU2HbQv5/d9WBesBZjVsL6at
d6zvKeP9LLyJzWpLbjvvctqQ3AbSv1zWJNi1D2Egb0Mzyy/6Mf773K9rpw5A7yTQJLF/QW2NPQPO
IKWxnhA3cX7d0HawuWG0UcVXLzghlxnLxxiTQBRiFuj7XfQv7SLTuR2z+QPBHLeU0DalFZePMsvJ
ECa4TrvO8pJtV4LFLc4dz9uVPImS7iGswrJbKjO+OtgPnHd1C5DRJS+T8VAZDNlH5ZBG7NJwcedz
t3L6Azf21mHA/d1JAvf7UQLYu86JqzDEY7IC4CMUohn2lG3nYBKow6/XR1XwszJsMuTi8nTE+Cly
ZBRmscH0oXtoS7hJdhU0nzrwoLc3bBl389teAn5jI+tsQ29PakdTMJejSmBfZFcqrcpA49Tng58n
P24qNc5qCQ+v4zv4GQmzQp48CFr2BvP9ZATiNIM4lBwFRh9sejGqAha6e5TvwOshPbt2zho8FLhm
U2vLMkefQGR5uyuEK5R/s/S4JLVDNoa4UK54KiAerYEA4PGE7XMXDgXF+eKcmssiYQi6uF506Gip
/Yn/Hmq5BOncwPqOk0npTSxRtG//txjiGDyegOavpKRxQf1wWaRE5E+Pn18AvTd2rn+1rX2oa7ky
jOYqhccStiA79AZt+2lrRgoqNe1rpiK7wBWfD4p8ij+JhApOgUJu7SPjLehwe+j2FuvtKXT36MW0
r5RzTLQ0IszrsYF2ZeARXf6xbQQh6o4rTLEuFcabaBVH+zMIrupu76di7IpGbOvBApypLDdPQlyJ
7i3JI4wCjq/S88YAE6hYYt36LBAQnxOEJ58eSqauaI8OCwOehN3rCsXXhn5nnz+wKLXfgO6tOS2a
MHtGWZR83HDezwyAHEJRz8K2Aav/X6bnPIBYxYkvcdcc+F0iHjj07RpG5MEsR5+1GpaQihQZBmMg
YHOVW8JOy3oKE9jNs2pxom6ZX1EJ0KJKJXU3hNjIiw0civBNFWwDWgpQPf3vpcdJsI+u2HXoL9Tn
rAVeDoRHxEIVrkznS01+zBn0Lyr75ohg0bxkHJ7pophqCj5feRlCey1j4qxgMVTqXAyZQe0Igk2R
Ns5VjkK82wfywTKsbADPefx/qszq6CMpfM6EFA8IfBVIlv70DviwEh8N1Aoe34DkxfUGMshiWfNC
56moTnFw36a21omsZu8GBTCk/vMHm3M2uVHQjzEJnVSrzFLRRwFvzLRxLTNhH+sTCwF08cMCUDXu
JWDWgA71qXSJfvnIjYPpCGuiUVSBEf/zPpQAzd8CRFNuRc5H9XAbSdiHZu77VYtjszuX9NqDsboV
rXozmJLmmS703xjgj7YNRKyKgNAXBMLjq3YZFYiYK0g0Cc9pS9slUTSpSxKakstI1chzjQJQPr7v
8mWsfBWtWyNciRSZx6f+g1qLqxIT1jpv9k8vXgfn/zAbuMbXslypJpnUIJY3CClOlPtHNkE2vPod
bmiZoiaIV1X+bwPvdUz5rvLv8fb6xLcodIE4zHxoPq/FxI4Np4PyVvqgq6yBIcPy/3qkYCd5bGkV
vUnpUpX/geQu5EDa6t5GB0LJIlGvr0Wz/6VZT7Q20fW0rHjNPryoxMejSGQArrHnB+vdAu8umYHc
sdFMZhLFo2wv06BHXP4tuyVNSA0bvZYeH/YuDqQF+OwJDJc7unyO7fjMD9/wcRfqGLJE3V52j810
ghvUW9oX3QGkLRnTARFKbd7f/wU1zySk5+1DWfdSyWVcIvwanOzedfKTcDNR5UoH4mQsy7rxUMzD
cCacOaDz9ZKAzHDJw/5D98KnBbtzjcVJzTE3m8h6n/Tk6HPkUlxGUMOEK1NFsGJPoz8cq0E1TGGm
L/GIh+Cb8ME06OsqzbJ9xQYZSkvbgMNHodmHaoK6Jwef8VzqD6C6UsVy/sZ23AIp9qNOsGBtCGgs
KQSZx+QxhKgXI8T21mmV0n0A5H3ZHLFMwL3XV407ymI/4YIYujoUjDGoVRsfiVi59qTfZPD9Am+H
1toZix4TLrsvP18vUqJBpVFVzSWjp++Gi35cmB4Uo4gzGieuxQhymcUwzeBM+zX3136i7YvrtEut
uu44MTfMrQFdGeCMGhLd9OMRjBflUtbxrW6AiO2w9NkbuJaNQoh+aBIzaKqiS/sYo8AlrYc5gt84
ZyELc3RlQr4S6pJ2hvJd3qjn3YN83fy5OaBAm3FmjRGq0B1+f4JlDzuBRdaoyvAQ3A2bY2rLJPZM
JO52mLXTjvtgDzMM1AaSdby/KN5rn+s2OIJArU1dCv7cAUPs7gmZ/nOZjxBWX6G8pNSHnIJVWRFN
KMABf3lGQPezv2FViz4UqSfiHPhVRkro4j264dCY/h0fGQy2wctkrAxVU9z7d3f1ay6DULrTjWbO
d9bsTeLUSKeUEEYqHNXr1Kn+48jBW2V9lz+HLPDKfWuXMzGLQpP5hm8orD12PZkLlfhD/OihKAuq
jkCa5UOYqKOqLXxLvS0mNgGzi3+TthhP7st8eta6vmlA/ECiMlO4p+49/ksjmF9cQfJXsMzxyhzg
lQgwC8ayP8u5/3KsGXspKyc2BnisnQP7ugyV/q/+/OaW4DqTwJLZNxj+Ple33iyBrIelLn6epMJY
i/dbflR2brLxPEU67YNB2YzQfiMNiXxE8vv/kclVVL2B1K1OoWcaTVZ/7WT1eWfxy64UW8Cepzie
gR2rItoHLJLXQNR5CKZiO4Ur5eurfy6Q2eCo99UG7xHEud30xU9vi4vEwMU6Aake9//wEFF9AYb2
kaWlk8Snqt+6vSNR3JXQBxY5Vh/0S9eMdFduJ94X3oRfgwbj6MprKvNOUXldSzGExng8OZIIT9rx
9JEPCw+gWd8C3tGf8FaCQZJjA2TR+frlg3D8fZesh3fb1z2tKoJW/LmbGdDgRcFOKtGsgeXhJpGd
H/OcEtcqt3ebIDcD318OnmemMG8vVU8i0wWsNl6Far7llneFQEARCfyVy5Gb+G5sZ5Upp+DR+mO2
+THYSP/6Tc5ayERaBp/PCCSaxgNch1R5yaXYpgfuFlLOkD5TOdDDK1xufbQxteO07RyxZhT4EOUF
QeL9V5iEYbKmXFJumGFhnnPVyQp8v6eoPdGFKGBLFWiozvmL7nkbUVF0ZbozQhDl/TdIXNvdHarz
R1ktQzXaiSwYn/+/7dTG4WRgppTBE1QjMY9vyl7a3GRpgHF71lfKFs8RX4NySCyCGThYdlTwf0+m
mndFCzNwEebyQp+tydhEtwFp7hYbx2mP8gQH9ULESGBnZb/vCCVShZ6trliFp5aZjL9vgz0ypqxo
vYibEmlBSuvtV8UWHD2QkQV7YHYBNj1esMrD9/HCCb5Ruhe+jHh5YD6nob9V+HOO/8ih+Cgjqeq7
++zZ7GMRkd1G+0hMHYNPurcjEprGM8bVhbYQug3sfMPs4Ei40SsGxy0f4GQ4tzEh+ew6Ra6zWkIp
5y6LwqCEtkR4ohNB0ZEC+aNal/e9AenyJyJgbnEDAU6cMnFBA/JD7n20J7BrYn+VmL1XQCOUk45l
AMb3iouO1vetbop5yPr/yXi0/vWa6flyxmB6bLV3vppAEv8ZqzGw4LXIREQMTWlz/O4FPG4bIWJK
Z+A9SxIpXWJoib/OEcL+1QsoVjUYOKxtCaPz4iHzb9Hu8V4Gsi+6g0PL9/0Mwg6JI+jA2ibcJ6Ay
Q13aiRqrZeEIanXPLaZ7gquBQqRzTxZrdpIfX+ob5Cikqayegb82fh+oQmSyLdJLON45+zDz7BFj
g0qLeYT5ao407yZEfyfoISyNuWC3n/zR0Mwmcm1XFzeWgpWKRJ0EtP3W3U/UjCLdoBcE7KkXEXQC
8SCWJdkn1mgg+mTYuxaQSaXk7sjOZG5Kc1W5qxI7UzDSifzHmWMw0NGpNYn4m+q5pBdOATABiOiB
Q+1OQZ/x3gXHN/jPF2BYt/4se4QJsroGSB2e3xvAOHTLKQJVNMRxXr4zWhhRq3LGSRUAXhpc1SU2
HU0+ft1W0qg0KkWL4BaVj/+JQ1Tg3HFUTZX0ZRh28qk9xHFsgHhV6ljFKVkE/KR2+I9H05KA+0hH
a36f5MoA0hA7l3mFvIUa8mPa64rCcvsGwNbehQr4VloMfS+BckEsY5u5M81pGVU90YI5oZTy0ufF
PFJWuc0/+rhWH73GBgqVFmVBtXzVGyzDpTFfFjAwiq0gQ2za117M9iYJzYJyz995VyVyHc6fxJnl
oPTjjHoYdG2nYZYktV/lHZUHi7m9wITrsQUOQS+/pZMaSjc+tuJr6CuLDFBvckZqKHd/Wu37+xKB
79YcaAhCqqqNoF1O1+nMmkuSz/5lmFdqR9BIHedFd1r9EHTGxFhBolo75DckFhsdmTUpHl8KJzZ0
yfvtGDsupokM6e0tHARsaX5cALkpEu6yPZ5te0y/0NQD/o74lIBma++nWQHVXBb6JHyd/pvc90dV
FL0C3Z8l9mYHUe6ZfTP2RcsYIaOYQIi73BXiWNlBSza1CHX7s8PE5s+BqmJFAMRiQH6FMax0f1pp
1z3U9TskxEEny1zaIxH8oedSPpa4XpC3EHCRFVnICDj2kjlv8m8TKe6LirbMQjnqoBCLfL2k39kO
SjMzch3d7LJABZPMsr8cpGNCuMYfNGTnrdTraCmHYBBZ59V9f0F2kivZFQfUEF44LeNzjNFk8D4+
TQ2Z2wnTkMrP2rhzQodkqhh2rQLnLJFHU/1DC0UNlu2MjKfuiiwwBRtiRJ/bfmUZduJWap1F8rhd
837veHPISFpLOTeJ0GIj8wFYuUHHR9D/lXrgZRqpKfVxKTnJ3CRlGWWU2JTDGxSKec7bYq4Pam2o
QTsKr6OzrjSOyx3NeJcIxZ0T4rRh5G5YDKpCVTXkwgyIAm9YTM2GQGvhlcxYBIzzgGTDXK7P7smK
nifuGge7eDPFfIye8X3p/vrZkEi6HEc/Gkc8DkZ8TV8FaIalnnxWCBR+ry5wp7JblvyBnc8MXdey
55pGP9ExrvA2d3ywd8SLmPUUhRW/4hymhkjADVV9B59j/9R/+ZRndDy0Td7FsRHw3yAmIUnlYnJq
BKOYx0bvDSuFRGAApOrho/CYExqlmvpqgkq3n0Iti4+qzBVY70FeiZhwlBegopZOMC/utVXLQ0nO
crp1BCe+vDFMhr9UCox4Nze6MfBXu/bTa78W6lBjjKxW78r9rD/kC1YFTuIsqgtu7Reesw/7xpHL
2oHfmmr9TSNlZOoX+9A5MfppDGRXMaelCKzPRNp1g9njlMpweAnLe2LOPInOpNv1L3dr/qHWvRjE
y02m6NW409jrHsFMEAqsC4C8EpXF1Iy7aEWIARkRZKWxxSmrGQyW2lTb9eEh6anYp+Uyq91eW+W9
6jgxEjpktv9jQiIA0nE5aGY1R+7ndvpR0g24I5TteEC8G6XSnhRGzch1yljdRpdy+cwnqHSjQ8iU
F4tC5SyFNUTP5+jWdZvRjQanZYuq3GIIRjNel97VwV1ZNjnBYniefmzsKpu5uHR0IkCxXDegJzwj
39Eb9iUnh2HYZJnUxSxK2m0GqOFZT4u2XZWm4zdV3Q2RJqYZ0CHYgHK+9Ap0/73+VVEUCempitkO
EqoUc6TxeQpWVfDF/jfQY5+me4GM32msiNZi+71GbFNOiwqWKRDwku8o84NIDil3TSMZZP7KJgb4
Pgj5ymU8cgO6zA3T8uDvEoBz3oaV5pJuOgSP1AKeGUEl+djdnrGJ1Zw3sXp8frWCO0a0sm7ahSc5
tmKPaajaqJ06RaFIiH8zFE8NrgHoxqsVBpOVTUaJFeMSBqpJmOM+mYa26nGoBzuSXdbJWxYLztp0
jc0QDAon+XCwAdZKjcfHC/icxsiQbiSPWcsbL5eA8cUaRivxtWSFRjJ4lObJs9oWCFqWBFm8Yl/2
E3SfgwX7dpT5mGkVdqCE6dq5RkcOMIHiNc+Ua2KHBRAEx22nnF9AqPKJ1sTlr0cvWWqPYQH8i9Sn
TF0eIL9igES9LAeElPMit2AV5JwWl5NPj1ToeXnrf/8k+pBp8sdDK/fLcwcBhXxGpOLyfvi/So19
I77YwqGD1GZHY7+hQgcOWTVbNsRIwGdwHBgutRwJA4QxYHI/cKtbt03vNCh9U8IMcH2I9ZFx3zH+
+7Hv5or8YzL7LV4A5JtP/aj1ftAXaAiY1cOHoIpnQUnxLlx/rnOqeBvnDu0kry68sVviJkaBjkcu
y961JQ2qecgcEDOrSeKPnPt2uSf97pTTVomsghq+gIlSDxjCtdeKjZOmV2ni/xopRmEbwMNp73WG
l4VUXwSvMBUMbDg4Tca7nPy8VPD+9nsjYMVn159s0j11PhFYDedgWDv6PaZUzDu8STmeUJ6k2GIA
tbg1PjWLRcUxl5w98pAnTwNN6dTwemZAX7rpnOaCebCsRT/zwaBRgUuGbiy9uj24SgKjNsHLsDlC
FqHO0Mih1mAOCyVCEuZ64dTHClYr/Z3GgDA/MeQGyW9mACWcouW/Y5FAzeVSRP3vECe8l4M4ISxM
nSf9U/e7nMY3CDLqJ8qDFZFzKTebOfZv/X1PabVDQ5a9sEpag8oVUGhjGdRwU+8MHqDIhd00tVtO
yej5hd1jzA0wrSpSlH4LKOsnADkEIX+fmcmftZpGSX+mGdLne7jIv9ELxHR17jAtNo+gVD/r+7jZ
JSCYiyG3vUBqrzHake69BR4r+Wtb1ooYHp+czR1y/KiXU2hQNT7lm16uyeytht7UYXH2GbqfjMPK
7cjUAHBSuGapYdmgKfxBhialVuiUMnUVBoz3Mc2TL0QsjW7GW0QTPJyu8iUcc11TaoTldRBlaAJy
qz8JHsZPL+5ujOTdqTmuNS2g5kWYfE6+cUp5LGgQlktQWWqYbyxDZ41ZX5+2IqdhG4RNFlJjpR+p
ZexH5GZ+Z/xViQk7bA+GgFBQ/WfsDtcyluk7wUihBCjKUyO9QJtfzml+feEJrPQhAhA5BDQUhex9
sH/KucbULSn6jk9dqWMat7+MxgPDStvEwbdotbILw30+A/ersiih79wL4HZ4XgEH9vzEky1yb126
Sgce9Syfn4/CmWNVOYG0F1Ui3Imclbpjw5G5yNjjfeQy5C3jPcjX2Z8YzVt0Pz4liBl6z1ohl6/Z
2d28g34hAX4Xu7o0MTGLv+j2IkrNPV0s83PVA+H6z41gbumHAk9Ykf06woMFQi8MKNCgI+ricxOQ
fDS/lbkW+0lwufAu6KxpR2SiP9FQG/379+fGeFNAx99qJN+Tc2rRPSJaFBnISbkERAs0nmo5z6a5
HrLa87t/H69YXVYadB8tOjR3BK3hiFjFk22ZNb1ZJfgf73iFw1XDax0Vt8vIIB4QVcYHC1uVxPIm
ydOw6cbBCiTXURao28CayWk+mOTJDZxX1PusZ2ywvX/gV4T4mhv6fEyQw5AAu7cA8VxWZ4oW/BLm
95+NuDw7pYSst++hy3Y82WzH9g3OxopV2ojVoTW2zkujv7mz3J3RFD4CmxbJo63rkq2xM1A/lgLP
nhACjMpLjq5I/6zPOYAa12vt+td2D4hJDI9mMvHslNzsu7HRBXcwQ7AhnMYxpIpPkSmkta1QYNz8
rf1LsJc8tnxe00MqF93Olpeop9v8Pf/n/RTQn1+dzQNCikqtyHuhLgnoghu0Q4LjlZfkN/pd/zN9
jhWj9rD4Z8jNTyct88DzISUcA+Ww1ZDV/ErVzin6xwkG+iCACe3ze0fGldpVf+YLPbbRW/xgMhl5
8ayouMNk+0X+UYw/SK0R3KU/mgJBEqH1ESXH7U0eH3Io55svrrUtDv9eofeeSAQzraEWtVXo/WmO
TtefGzi6Z6CCg98+YaWnRYuKromR2ujjq9yGCULvApERE2daTdgK/9pva/bGhhFXMR5r7Wqemdmk
NO3UI7akV2KHgxrtDsGbnYHFKa7rHiGn15uPuC2w9c9T2SYB0acCPt4y2vuMox+EWJbI8bS7zue3
fNYZsp82T65Wh/FeD4/qELhtlaiEx1HRtmtnlv5svvuJ3LbQUJd8o8Ao+kSbGr6bI60eJmLpU74u
5kgn5mkqsQa6bFO8HZNdM7OcjJPJ6ssfTRo6dhsg3nsGyMOPI7ziiG4pytM7RAAswDLfIDV37Sew
9qx6S9sY15fDkQxsLTOoT0Q0NzI8JkG3C4GRUQo3uGD134KL+8VBmMRP4doz7wFhAfPiDwX9fK1/
y49kReVzHjmRBR1kQBg8of8Qr8xm/IzLfJSEB3CM8cGAQoivNSuLoJw9OpKHn+7x1mF4mhq9Ieja
03B+6xX3tD1mXBaN24w/FXQYg8NozpZL/uVbqixoUfLcwYzX6ohI3zC1dq5OEAJNs8UatZ98Kza8
//yToqH5aRE9lNG3c0UtEs1YVcnpq8F0H76QdPC1JyTMq9LXky4/54ekgyRX7ueVTvaY2jX1lKtf
D9aIWoHZ7aKTSRZE14ZGjUqcQvQHEw3b7SIoFz8MA4qVcpLuWDauUbc6GaoOG2wEDS2wqztelKcS
jneehXZKEQSvFyD16CwlJytZNJXnB1q1wUiFOtbwa0EGtlRX/1Tr462//w0SjNwhh7oWkHXRTQxu
ILtQES68doJ10fGnLZllI+LmBIBPGubLnCCWMZXaCAOL2bIX64jFYWFEu/p2VkFObXxMMnvvNceW
jI9hN67/cqMZ6zAHjBThHxumn0TEYBZtlm+y3w5EVN0rA+xKSx412D7vk79IQVjnRvnEgu90HS4F
KtmyssOOSPFPG4Xi4rNBlECfqFDEqfVdlltIk3eZPMD0V6XzkObDyr7PclwOlx7dVXpSYj9dET+6
kyb63ohb394GiTWkWRJP2PlFfIMIRYWxFDJ6AeRsqkJYt1LDYdJqDKC6nj+96pSO6I1gihXUzXTJ
/9kfOpkR/+0rQRT6tf4IguCYXH38wq/bRmmOa3d/lkz7gFBKTNFwh4+Y4aDQAFzjvwC4PkrI53tZ
jp6Qo2g/xYPTDkyz0bR7J2fQThTbI0HvUs1bYr0FuWn09aNlVqICjr+LGrE/ClXJvfLtgxrk8k7C
Ny8WzPyvHO6wv7Ma1cAljwFqw1WDsnQY1Z82xAG5n3kvXARjF4kjZSxU4zabW4l9I176ZpHnpRPK
UYgAF6PQoexgtfkX3VJnuG0Qei0s7+kUeiZ+e/pufkOothBg6q23rbn6EHeu+L0L9VrVnXqk0dZW
DO6V7GmzmzNrjuQ9TPyzOwy8WmohwK0DCnKoSPYmG8yaG4KMAINGZPwVcC9ApLReYTcalXjJr2z5
tWDxQiKBHehNMTwr3GlUcXfI44OhTmYazYS01jAUSPXwPsDDTfRirfG1FcIww0GX8Ld2UXhBmEhI
cZO3hfWJhOHaGtWWavfuH6iH2Ma8dYA9F7eiq8ThzSLyuM9ZhwjpMrLCUYaLOHdIUsA19OIEJ6kC
Kb0+6eym6QVw2uDoTiNcJyu8YpDzZ2C74/n2+Df5OKOqbT2Xy+tMZ2F5P/M06sA3+8T0mqnqpUHm
or5tg3xSQECyB/ytcEZUOez+cPqjWpqn3FImsyCFA2j1233g3wXHrdV40MphC5JDsUYCY/PVEbVK
4OAu/yVdv4lbtU3xuvyC/dxmvHrwvnXi23iu7sDXQ0QJmsvhz54YR3dlGa+IOZwf2nehfyu1cUvw
Ou2Ff+XBgdmgmFnDKzOX4oxJrk3HUeFQI0KHULryZs8UC0E/xgKZVOQXfPZuxob9KBetDtW7PLnA
P2usYve9I7QIGiYUK20soueM9tUgVe7AubFe719BlYtYQXijCp9AxvW3thGcuWqXSnvKyvjOIwzG
WG7eTbseTl/RmfobS+LNymu98+BTrYUsInxgoW+9nbw5f4uj4YRs/o6sr+7z6g77sNxN+kRG8YV6
xGHqeQd02yV2oKVrBSAAkLryCJ8yUYN7CRCOxFpXOu5fuO3lpyMwBVyM/BdPMcP51pxWMdRHn9MD
2fq8seei9JwWWdoAXdc2o8JWC4ccgzB6CoY9Fqd/qF6ec43gStX7MrVq97Datm8i5tb2LwV2TkvJ
uFRc79kKW+8ftJlYI7rjxTVysU6ZIMSqJeznXpD8bGHNzf1gb09m2tKgTIklG9GxBDXZITZ/71if
wNqqZVBz0fqgCgtM+kNaFZ3l2tTUAK4G63DDd9DwlPL9ipI322mMFw6v+JDE5sJcNUY0iazNcN1y
jvJSbBLy2geVJn8j6Woup+OSBTjesbVhTZlsovO6eDmf6QnXmxonfq30RmTH+ie2X/ouAp3u4P3j
TQKfYSjKKR+rAer0ScyRNbIorOi01DE1ZITCo3ijiC7FswGNGyGaCtC9Y+TMq+X3XWtMVfH1SRUU
n8Xd5YDEpxx8OQ2OdvBb4eQWbnAFIwGJanKUd1e52ZuVYVGT5MbQKoMCYgbV9cT613BgY5gwV7S0
RExITEq5NqZYVzT//HzqnRWRfjmF3gItnATzdcrxOs8j6XFaZd9Y0WqMHl01bzOoLX8B12bmPYMV
zJDt+vLsuJJLnJDYY+5YRt5mu5EcT4gqQlJgAnL0u/SOb/U29Eefrf++1ExjUoWRq4BHnEA+PmzI
D3QPdXci7O6O9Ckg1I0shV1AO2ye9+3d1s0cJGKqK+DowWYsBswbfItwo9+jNOW7aRuScMhxuFoU
470xWv62pSOj35vVAo4RQLkq7fTv/8OC9pn8gmAdQL2CqfWeyvkaaqsYfY0EB3mDhNbKUdb0XdZa
1cdvSGnYJNgA6R7k9vxylPEWQHL+OrCwdRZeLD9fVHtuJlFRbctGKQfEeL1mXhy4+o4q95V3/UMk
dS82R3pPcsuoIt0EpvU5llpk24JjXP5vFOX1UrLpnv3UUrhQ5pCixiNyfzLwovMb1dMFYljITnZh
T82WApld/rTrgYNJDxPa7uFcRj98m0Qf+n1FStJ9ZHmAKY9B1WHCZHizG0GEva7LCNoVl+zlwvDI
lozchhrqxb6Y7Vq0ZRfpHV9FNqykrSGIcdkg8CRGWovsvPkFENqeiuc9bFWMY7OP8r8pt3CyIkAC
dLFeHLo/cqIsO3+9gIz6wto2D0lnblz6UCz4KgKbYyBO4n27yoGiXT6eot2XTAlPmiIm1bU21Wic
pW5TOa987w5Ui8wBSg81BMKuFAj93cVQ0iIqaIhmvY8Tfrf8l7pZLjIYo5rKu3zn1ctRloBS0+5Y
nf1iVun7pUtcdyRcnvRTu99KroBeZtw/v0DBbP2DcqLS5jYPKWykR/3rwP7JMW8LdSh2v0nAU0Je
D4p7Y53NIXRG6m3q4TtqdUhw0Hka1oC1JGbFECDc+a46hUs1jlZyk8v0nT1YnLZa0EITH/xawzQI
+sh4bXOWkxvfDe7yfDgIM0aLA19l7RGS6LEoQLsKYcKwHB/SGBko4gkg/4/Xr8T+TFo/ikVEfcUD
4Tyco74nmuMR+ekW44igHHBrjZmFUDqCrCr8VS9ARC+ojMIAz6ISknAGzgUkVno/VO5iaXTRS4dr
vQ1ATV0FEi4zBwuXtGTJDPKNT6frrtBXAvO5M5udGkBICKqBG0qVZgJS0RN4QQyTu+Ni8ynU54kO
j1JBktoE+zdZOTZ+98o+d2DjugkPFqqjHzn8+5n5DYA0qKuQxlcv10+Apg2KuPvpItvhzsyyqLNM
8ocsle7990zfpwQrQtriNvYJRIfYgG9g7FEnpO1dCn96g4e07W34Rzlq2q7iqPk1gE62lcJ7uDjF
kpHuGiofrdSCsbLgC3kjlyPo13bTbZgkteCIMMFFeKmLcQs1YtD6sdZtiSwuqkjxvf2QEQZR/F4e
Sd4EpQ9X4i6t2++Uh6viokrMTFAslPPmxGRwATwUhQR7nUDxmxjlMQIhNqtWe3b3eH5grhsMq7AI
os8AuoSqZk9nE6+zgPcakZllPT6hGHopxgd+hs0c4ZB5SkIDxV6gjFfQQpWQCmuGuzkwa1WcZNTt
colwQJfKxJTKvceXzt13jP7vwd0d/+Jo03SEYf97tf4s0OcvZRz4nQvikiswvxQ8mGz1TJT+wMTo
cjkyi7R3j8vYi/YBQgjUxy4NwDDlJPUOIuPTBV3770Q9a+38NQGtxP0wCbIVkFkz8sgK4TplCjIF
iRSCbFpDf67uYjVJ/h/p3Hm43pprbxyMV0jxh5pAUMovIf6ZUOzTJw+MruOe8N83KFmyTCTkviJc
pRg3mmG8zZqb2GoK3hXWqv4lGpgxXdmenxtOyQdulQMD2k80fthWHVl8VBncU4Jj1z9Ej7Z0Rska
m6FFJmD3SDoifxJ7f/LV+2xOZ4fHZxOLwW3MVBjKWAbWrUykxEcduPGH1Vg+uIOliODGBrEPWVyI
lQ1PTYMDbEv9/B+cm1cgGcOerMa8yMlVYZ5GitqLNeCLPOOGPLOqqT4boHBEB3T6Ps7dh6z5AYCy
JOWA589RclmrA/qyj2pBdP9wPQoGYiOWArAX7sKIdjG6coSMcpK95sqIccBBhv8hduiJJUaBS1Ww
ZbGlMI/izw+/cx68VX9BrgoVoLcrzbsVqmrL/yknT87yv1Vyongkc4Q/UOH6aScWTx2jbsW8Yo67
9ytLg1U83tgs/Ks3FO1unSrl2qY2T+2Ccl7BOptUFxt8q3AVodDbbQJIrdcfcprnOOzvKyZKj9/R
0SqREYPkuuuLY5i6UJfAlqCLy9/BOImjVf7Nm8ClLsrFNL79OMdl1/sJN34oBStKONQdkbo1sdYE
VSHlhCU7sjijcqRYkxRkwvWOWyTCIqO0AR5QhUqwsluUMDtJd6HXYa4Z1PWJpsBoaDxvfnDSDQGf
2fjD4UdDvAV2jpzvnlBtmBxnhpbtle6tzqm5W5DGG9t1+JnbHD2qaiSydGE+1l5lM+tkSlJsRIsw
23NflhksQj2jQfIawxzIT5QEXTK9ihedlTj2t4Zns0/T4PufX02RCv+HqnVn5mO8L3v5HqsFAtaY
ie+eO8zqnYay8SeNwFte/fQxT9PjPJ4hdtWdQLaychftBfhJAZIbuiIIHtY3+47gIRl5I6E2gQmK
EkiBwaxgo9nU50yBpOakylKs9AgPo4w/IPkNvyay4i4/fSF/2jfx3arwUNe14z/zWKJubtKjeHXW
9btOP3yBhEwxeWhUlfOaP+4ZpVLEiTH/lcuI9pYkTH1K6/RLwCpBBHA12ke+gbEDty91hglpK1M3
hmUjM+XK2PURrHcRSetanz0TDJC2CC+D+XsxJtt7y9Od/0HOhLAtlFJf05M/Zjh0XqJxJkkmFN+W
qXWyx7UZZk145y99C0nHKyGvdt3z8wQ0vjbOM01NBK2eg3nJB7kVisfU/DPwdRVOkcjHGlDvOZQu
Oylq2+fLsTFdX20rkWL5jOZE3RBZQrwhHBwfb0qbGtbYKMPkR9Wne5y2E0yQRO2tUgptXL8fQNgw
5HKJhl45P1sUf9Jc4jsOzPFxjKytLhYVmXajWPsZnmmFY0wu9THwjuyc3bAY6u0aBpwaMOSANt2A
5PvKBHOAf18zVOvh1UOa9dW3fcX4gRL0y90JRknOa4n5AOrfEkR3Uh0bHDkyBzbec/Fhxber7NJo
Yrnen2GFd+aWtJKdjeegxINiYK2jJvCed+qHKF2CDz6R+N0EVeo3dsNJRvicYiX0tnF7YM/kZOib
1Bgfv7eC8ScyDIGc6AdywJ1VYBUGZuyiOizjAOwWP2eYcuY170wE7jCheKm/sZyp1cLUeaZOllvU
KJ2inKZbadHLj2aQRbnCaUWEdfHVcqHrQOaHV4ZyDGAtFnSjiiLsf7CDxx1YLjaRIYlqc+4jdxZY
eIaxn/iB/ywnnEEFzfuDrjVUMd+yET997RKGKOvxZ9T2ZyPJhABzDT8csdgsJAnFrTnhDtR8YAN0
yRM9qrEEr9gwJ2sCexsEtTGFRlg9yD0gWLar751QUnsA3JJd1Vj2Im39ZOG51XS9iFm+bVt5grEe
zb/RXsKvP3UiyNsiyBXxG6fPZXhGp5JBqsCRLN+MQCi+V3K9YbCwO0/m7DO0Xy4l4DE45XpaaMRx
20DkOQAg7RxMNe2qRMF7HmgtUxa1IQIK2NPnrJ4zNicwGooCsSPuJCXShtgM/2x/m/7KXVcTQrih
nUpMR6iR1RQLmgWx2SzlQIYkr4z52Hmo/rU7TVXOUimjOoXS/D5JYw2X+NM5BWRDZC01HQYWwDe4
6KKnTxggGN/ZxSNjphGC96dmeid8R7kSYdquFwbtiQcF7Lmgr8NHIscGRVGpBJDloLMHaUykd58L
aNDmfAqk3VVLcaU1R6ojlw4zFyz51t57YhLwOGkjNVS5XO7jknMrYrnoBWSn6eW9lEGTXW0fkHcf
fhHP3jXll6w+WMEWI0MxL4oEICqd9kYYd30quy/60XOG0p7HOyWdaSeEnixsnY79T17tWeYCEE8H
T3MOXP4wJ5YlV/+f9f96rwNJPQTXO3BQV2f1IYxEatsgSYoCf80DdoRF1qZKeYfFX+TBG/KkArjF
wDnFlHUpWHeuen99+ykiQ7L5IkLPg7prBriRXPkKsl6Jv61v/vc652BVxMTA7+VSq6tSTQKseVhs
ZlWxvEf2MeMoepJQKR5iEw9DcaTkRmeWJywA7F47zs3H8V0WKtzly8qFHiZbIChOg2gLm+fiSQ0a
VndPRtDAsPo2l9ELIsDNmgK7pXPvuSM1/qP1krqWu1vcXpZLRtRo3VtbbhOufXUtqZ7NpjNvMJEE
7KP4Cwb18N5Xegj86RlwcjQQlJiVoDU2g5Rle6JVJHJO9KV+WbcJNU5bd1pU4JyVgM58Z7B/CbTI
+nOn12E8M/vlMWp2FpXbjag6oZHn/6s1lxFdAnjhi1zzHcNhC9MiRSUuNHVib3Z9WQdDEjmX4gGv
pLDQWTJOzL2jODli0EEgMo4lSG5JF/2yBcV80Pv3UDRggen6fMlClVG0hGV1oSwrtH4dskaS2gA5
ZOi+UHVlvPZ334mguJiQpVPOjZqWPflMflUjwgKbOsG3+3lvRAEEGtLlOOK52q6vSGRlQuGIKWAU
KZEUR3wQO+trz2G7b73ic9jSraJzxAYFH1NYDFDUFKOrg5e86Ladaxi7A/KGsj2TDwyk9hCB8hFm
LuQY4V9Q1C2MZ6gdGp9Y2GlWud4PV7WVLZfgvNCrzAFIgFAmteGkkHTQ1kIMM3sYqlzknA/nq8Xk
6ROjtvAVbHtuPWP+0UXr+purPBAGKvZyG8mSRSZFoW5JnrMwPbrYlx7VT+06ciQTLx1xJMTPVR3n
0oCOKgk1ryCA/f4raTcjx0Vme0kN9wpZvKUomYa4JmRWnZNbHJG+1rno8lyuLZ6TidaPiOfKarIR
7uab20+nPobNfLooTQ7x6l+2H+uajqvU2EKbV0yi2Pxzz2kx4KWqifYaQb6InZfDforXLhVE9Yq2
TBp26tDHTZt+0aNKfd3ln2Gj0dwdHfGqwTRK/mX4z7owCb2ScWiRHalU+q6bl16vKWEJurZavxb8
DLMK+AWIEOyqKVWXJc1D+FCJJ81LQNsmFbVZhYDkwmr/i+2D83f1F/yOLVBIFojE5dK3jwFfziWt
u8gT2wgxRib+uPv3jIXCEWYqvZwqZbX5rirYJiysaSlhTCSMZ+knQii900MhOEUh+YfHpXfqCkKW
ngyWdnSpKJFdwy+kBEnLT3FnyiXw0cODmgBerCA9TbpEXglcpjNHj7sFGjlOfY3DK3l6kH8eWNOb
ai5VO/jg1ZahIlNVVXquC0mAyLZ8PkFZwPC2lQKFw4nWNoaVUDgOGO9y9fAP8gavpg3qfLajcmGo
rwlKxbqTRbSSAQOC4NG0dcnJs6U+kzca60w9C7MCt6IoEB/ESeskUWuk2/1PAG4gk3PwKz0qCcbh
p7jJN9Y9CVDXb8LQ3uM5+YYnmjRxvF93KyvRBm4mXqD+hkbg961v3IhT/uGJ8ptqRrI8ZkaiEA8d
Zz7VOzcKsQqrwAvES5GUI07RwhhYQT0trMMwG4qQBCD5FYWp5TVIJufxMROBiuoKyv+NqwPvMW3e
PsQk6pmbmM2pd7zI6sT8/FvAlxj/Al5WehFHKFO8SXXhSdt9OH582r89gdudm9cimfKHwuQV8Js1
NpEuwdjV6oRJrqP3ZftNQNdaEJMYm8l9/l0dfOWRhCv19WuoKSxdtRwNS9RUDwl94rLBfuG40qxI
WdNHTQSpGJ238PR81KX7qVrGExV7h2SqRKw1ZCDenpzF/uix3imKuLz69iRqvCn1Mlsk+Kboefty
1NMedeEghQwqoN70p+knSmvQJ0vURVTLOp8nlZYLryscwZy+yfVQJ5iedIP7xDYw3MsBc04cKuwJ
9e/ZgCySYR3uuHCQ9HeWbwOhLC4UN/9t2nMIeXkJeinUkEb705LQDRZ7hMhK0iJdqpIrKXsJUm6N
AZFvbUFThTtnHZ6s3738Tk+qAFObDsyPkEoqT5IA8jHUGngkBFmqLAPbt1ssi91L53fHOLovk7Gu
7EGtTWxHykYbLZrB1uzOPU0xpYZAs0GCm3dZV8KB75ah/2bxALK13SoRNGAlUhe1Ae9J2wXink8x
IGrZ5WAKNIM1RimsoINzAPLDPIodD26Rz5soHLkQqhKy3sWA8t+9w8jQUZIy+B8Zywo1H2ND+E8F
BQuCwWJHZ7jF1XjpUMptaEUh8YbbFTOvO27yo5HSmBp3A0Y3nxavvccyEgy7XGnzkVXQnpGPu5a1
iMUKia2IR8EvHkzEE2CzaRHTHUHPxCuri0tp882oc5sDGOTxuF038wIS2s4lFAn48tBoOd/cu9Z/
VNV7pDSjOU9XR1v7Pn6LnABbgE8PzXAk3yXTjUoAuw4yI65riFIfFDS+eNr9PHztsXY7P2ETQJ9a
CsSIL39yiFLsZvaww3LXGD6jz90QcnVjgoIZRvJdWXo/Ep96ckFRp78a3mUXN1143htZBzr30zkm
vQAPMzIvi1dJs4NjIbHTAy2ac5Z5F111H9lfPWAe00Wocn3EeWK7Mm6+bZEQUi7ankSZtuMu03H6
by9EGO5VoeCuIRu9kaXiOHIuKutaLZyq3OvSq7y7lGxWYxI/5tGjdf/Jz8azKF+XHCZ9zZffiLbN
Ly/U+M0HulJh+MYljiVr8+KqDbxkMaei9mXMTo0n97Fqys+g6KQ5Ui9vNsPybkSbRbheMMaYdOv4
x2ODK9JQG6+6c62dIA2PCmwcrlbw+iBS0Cv1mqn1m1PkbH5Lj5qpfHGajDNIRbDEejLrkKm0zrZS
LzTEGT1UCkXgwkDvdkPgGZkI23j44GmMCGBfjA3NBfsidzFTT5treqoh9avqFWlFpuXr45M40jTC
Bh8+6rl2j9MkA/4SKQnBQAMo4rAHXrE2+1RAoDj3VbBFEJqcX11YjBLu+f4quDg/2DAJAbR08iw+
Cq/1fBfHn7JxRWz8yNkGtFn8AdlRI3bmB1kIBlulkhTsHTKaX66D61hx2w/aC/PY/oy2YMcZ1sae
yp5CHzEWVM7+92qTNevpXrQcHUq8Nuj+AnFyOkx/571ipARLDmsXilUIjy75yLOmzvLb9JOQDtj3
ZwSirW5KevooHPf3uVYkMWbenWV+X9w/PdFWjSz0vzA4BstVriebLG6ZypEq+w5p+UPHIaCvIE2n
JErPU9iDVdm7sItzGm4gHB1xlCPhjudPteCIDkGOvSL5FhlW4apozgopx/rkiuHMSoWb7ngirOlF
ndxv+Bh48NX7d2DAZCYk4SWjM00h4Vz977v/zmwxqbNxGT5esoyfs5jUCF0DUK0G8qnRTH+njIkx
7Bwda+yWDA0yxzZj2swjCvUQ6tysTSLsOdNPA+fGIexjEn67Z+VKUfcKxZg5r3nALAComaCqKVf0
V2JvK1RlMQilmoZuDTEAFJD3WfkFV91cy8CDOg4VqPqo/n45M7N5ZjiFgQgWeXw8iXg/l4hxasoQ
mUnsOZwfJGLPn0Y1yeqHsBTXE2lkVBGxGXHfcyTlL/cd+vbgkw0V5YzFFbj7kGFYdXNIrV2l6hHD
IfrxAiD3lvInV44vK2TmdMYNZCc8zqWCQej2wH7eEFLgfivrzU5CNBbD88otM2S4jz9Y9pDvXo5G
AWEH8BloMnpGZ9L9z/khmGtI0m7vs4REl7N8eZXDFnmpu0BpCxcaUblWKR1D6/vbiLKCX7X1HETv
jYPszy1txniMxOZC9qc1sba3q6OZjjc+089uxtQ+PR7o65jQavmP6RewMuARUXCD8qcfDtcMn0gb
cAtXNr8HGChnoyJEJcyzk2hySkq6DC1hgInvvWUs3eUF93ajZAf56DlrWiBVP4EG65CsyeQcROVc
cP4bDONn4795Ku/I9pokGwbdyczKsawrHKInu96pGLgDcyDgdOIOxf/tIcaFHeuf15jJJYOrLdDQ
xmxB/if95COUNMo3vyAMb3veYi9Awbrvavy7mbIa3ntqnCrh61JYxC5/wcvdIPZgV+WmRhc8r5fp
+QQzwjwZrR6Rwazey++Fn5Va6y2SsiqYuhOZyFKLsjbPEzyxDAtJsOQLNnXhjGwouC6I55O4j7gD
QVVG+JYZ8fQEQWtAkoWNdjt1CbD7jhcM1WmuWXaWuqsZxTOSx9SZW9HP7YjAMtzVZVetabh53zAY
JXiI9yFyKBoxpQIvZG23RnaTt2XanlWJ02sXypzjX9gc3KARTvJ+XTLZ5pHzYD/EvqjZiYKNYd5j
MbMzWfZMDTKs+DMSd7lzg6k3ExHmEQLcDBIw4k1yIXna69vcXhgn8x7ZI3m2Yka31Wsh7eKCYOhW
oGUoTa8UXpJzDdGwidK54KhaKmw2D2teoUHP7+8TqEHZ9fKnHKtLrdY03f/0s1MFvcEyMWPYf8E5
0r4evy8Yf3NyviEGxqm4eHW2imtfv+IPcPtj0PwzvJiuIb+VKzEAorgWlyARmsPGWda4T/A1A1EL
jxEKg0+3WZ33ayezfq/jOQKbMIbudE/1jid0U3JN4uVHwxGqpmktZC7IfEG4wXPpUKSl5AA7bmBl
qj+uXEqJX8IbZhATgTlBbL00I3EZ2iSkm0S5eRvmiNUgz4+F/3bX4ZqH2Tc3oIz/9NJ1/Rqcxmic
ilxE2NuXfV4YYCGV+oE5c8ujJ0NGWRdghIpE2n9/NegvZWb9V2vzpk3zt2GqB5z+3rXhPvCmc0CG
Ebo1/tfgefS1XIPj/bJz5czYH6R55WxcF2uO7lQC/D69no+jOiRhQr1WsrPRopChJSJj1rX87JP2
3uQ3onIfLesQR51ZCCefTrZa6VfaxpPOYoEiMscU73ZtcWILvb0iI2MJANgvHlD5eTYcv/P5igxg
NGcWUdT2puaN01HcWknXwqEdoAcCaT0jpycVL9K9V2VEJ6AnTs8jIvqmIqVEEmwqbCpfNpciTPhp
OHPadhBrxmUf1X5CNSbY5+Ivu9QLKqXE23poNvHJlORVRNU2GIU19X5ZcUXUrLKJxSG0mraVEw2+
x2HH/6VLD7/4y2CijX/D4/ZAz03UWNwtGCKC+Y7j/VpY56Y15NK+So6ZWQ883DGNePieg5/7kMxJ
eyAgClXG+0T49crPSWqEJGKwS+7TyqDETegbQc5iOm2+fbgjQ2NHToE8B+bTAXZIp290uJCP6QN8
r/Y/9uuZ1FxMdkGMg6rgEqoF+JPixgfNEse/4b/ZXbPDztU6z7VyMovTN/IyNaYP8WyQk5G59wac
KbGZYWyP8Rq5QP1T3VIk0bITI9nrVpVFJbG4HqV5pNTV0KFrxQ/l/rMbaTffaJcMPzLUbR9n+yFS
J/Bps5Wy12LW8u3lprg2PXIebBYzjiR2UqrYoIwUe3uE+27jm/wLE+vkeLZ3cHTqWLJUmZX96MXN
V0q8wTRgrarowy7xgD2WYVxvLulQGqFf8845o5QB7RzL346d8o26oTpn9GvrtMFB829dsKLMQYOA
GR5ki+m85HtRrIY/zv7pBTO/+4GcSbOm1KqacYFtKjV9HPByHRnU3U5HkdAbXknch+aME/9JHC+F
NAO0z1L1C8CUWWDsblEPdjWT+vzOggziCK4NZaBd06NtQyu+N7KoCRRmKQ88H4JmGaPhFxLAcZ8E
AG6zJu1HiLKaN/s3z2uStpasyDZg7QamcS08sIxGXqEH898BO75ZShyGw2CY+6Ye2e5x63aR54H0
ewF2QuSczgywa4curWKWCPhQYHJ25rPpbXn8n3dGaOYfvx5fntTVHZP1IDdm6G8KC+JTa/bkX/ys
Y6GcUItS0S77X+TEjIuwkYvy5E3YQeG1lARpKcie/0NzySg4MNHeyLmPemr5WO++wGVvl0QVKZY3
nA5iy1WT03Xj4zZwbb5e+MsRmD+7Q1yBu+ksCUNoIb1LYFAz3EnffNfPqtt7vWO7yg9qr+Z71gum
Po9YeUxFdT4DbEZxXbEcoAcOMVKElnu+our1XZzfNSOL+u0637/EOxbiWIUlpXqXkfNvH9UL30IB
WwuzKOvH7ichpZwzS3bmdr8yf3M9nNDWXgT+ks3k7LHS2ZNUqZflVMEkoAhU6r46j3Dfe8PcUV86
jcmFmXw9xgRG13OO+glztoFITGLydEg0bKXzP6u/qw4NCSQeBI0EDX2mtkwOW7CYiHjeZZ/+AfPT
h0ZckqgijsWjbueBfDk5f2OB1ilGPMeBRKP8bbVtCdNWSwE7J35PhJkUIv6EVADP6WxkZCn15i6h
6Hw8oTfXKt5J+tOGE+Em8ceTspXlGyv7XWARK4GEudf8+gAQDnBgtepmlTxGaSio6lEx1F3FHJqW
i9he5mfzlrl/rcmV+oE2969L5Ga2grgjn82dpk5H7I3zLopoduVfvwYY+PCy2+pnLcV0T/ufB8V2
wqQsRbAlcT1HwvA/9fScinOHiqficgVDuv+UgoMdjwGhuzkTpsI4AmiT6baD242ZuFEJyNto75rn
B1dh3VK5veTmPE4Ua/+YtiyX3hguIqrJmB3zZor87QaQ9VL20lLdBRTedNtn1AXweLmBvyUcccY9
Y7ADobJkfp5awQrshFP9e+D/3TXVdnQI2n0WhrJb4AXxLiDFWSkQR66wJDieFSYMYyfgwgSwJ7hD
aGafnLDZW3CyPG6akjcQtmW066Z1P5jF212pouD+vf3qZRJw3lTSR/EFuqXVwMmS+dkRkzDFAhQb
kZZg2NJo75q2GdmnwwwpK0UxzAbVZ53F86CnOIQjsVyteWX7VQiqQK8BbBoFV9z7R77ouunUKrmm
mVLWUMAGNp1aqBIDzxfIsl6jT438iOxw6TIPfycgI45LaMQed2AOlQ4gE1qLSk44taCabDGuOXDo
Iwi2p8mDE0YGZcdp16Htp6aSqs0VYqt49lWmE3lf/T9QvdlBKv4ogST/h3FaGzlQNwQiycagP9oz
bTL5/tXL5Q2Z5C+qn55ObWRvS7rW1V1JhvWidBCiO4MTSgLDbxssxPRGBYZXl2uXrBM8xNJBMttU
GyCKcBQMIL+ozZZXE3tI+62K1Dd8ysi1FcqvV4XzTbVOhvrj4HBhjNhiTvDYbVeEVKjj6JWBAIsr
BUwYT+oQgq052pwJP6UaT2kh8uGI5w1iZ/yNgSZGahDK13z+lZH8YzbzcFwezxIt4Bcj5fIT23fN
SmydVGMAEHr7SdI0U4KKx13GtUnfXD5RAOpSuW7qbJCELQwNY/asTT9/sSwcJHMHsKpb9npp4Hfg
Oj3LOZAQyvE1wkfQ6eqq18G1jFdSL1RNJsFJAkfCmg3Bvsz+LeqSNy46j88/rvI4XYYG5j4zsEO0
sOvZ3skK3zup0i0RG/rdCVg6yV9EHmjqnZ5FI6CTzrgRt+rUnj/CMVntlZvk/BhDYpnRmiiwkIGc
QIfAA7T71808jlsO26uZ0v2t/slk4WUO2n7SM3A2d1Npf9n2/M/6aDRgDllGdvjwtYIodwEPCevE
YIqXarWTc+gvHp+hxsdezbRzO7xHTixB7dZiYhhqVDtN8z+Sz+VXIrmoKOtWq9TRaElM+fwdFfzo
flzc9uObtk06QJFks3ltZwcugxkqbCDr74ZoqNPT6CshEKDSADutUZKNCoBLmOQCDOCCupOGilFa
7btUWL8CiQrabkHlbF24mi+LS9ooS/RaeVewU6pBVHVCEJeViO86I+sorWV3mQWB4VBlY4Nkcdfc
mxqHhAEnuXtCzif7iLVQsjGuGG9DuIkBeso/huemdXGq+hANXkELAP0lZo4+jQrhu+/Kuf9Pp5lN
Q6A5JaX9cr0J9aDYETQFZ169826gf/dyF/9EMcoJRHBROF6cbGh8DKc/PhJt0o0lQ/pMcJVqZq9f
HlMszzQfI+ibi4MzqHdL/9+4ib4gBqUY86TNAxIlf2MGRbxmfhEUh3MCd/T8fglEJKrEy/pfxMec
qnKDOwGf0FvfVnPqcZf+k96HM891tc6thFYehvqo8aOSGVSde6opqkrgjnJGtaFkPjUXQvnapt/k
r8Ou50RY+a35EXG/Zg971NPAk6+NW4wzbmmUtpnxEuR9NnBaoERd+nG6J8RJhyFQCqouWVUekFEb
7rs7iI1YzXn39za1Bukud90p7j9fNWW2/A2OGIvnIWY4wIRq1c2p1BAjZo4aeP4wM9dLpxAiwGIw
mbdjwOwWz8cB2X01pcvFAtUcImcpextNlYeT7R41ewgxQjZDSdkX6iKvIep47X/IIl0fr25gY1yT
vmzK6l1UcnKP5GVIuceINcSr3Es2+CK6pPUnc/yOOFNXOWhLmvI89NfBrMTk8Cu7YuBU7oLKmn58
Ij9I2ldMTPW+/ijL+Q7EcoMqr0YaLY4JVX3H7Qtoj7sUwHyw9fY9GaCc43PqEXuq8R3CMpEkqEsf
8vS1DPEfPGN8hhwOTQbgQLyQC5zNkgMeEpqP7WfuFfwRB3x9xG7EpGBFI1x9q3WAPAgSA9LryXwk
/1YBPitX+f8kicflGUMOPnLeMVhuA/9o1PllF/1xy3jJ95r9wDyW/qCWihL0auDSauBzuLik2b5l
1Sh4vNKWgpW5Lk0+jlZzNqAKzU/DsZugqPhjXK811ML6e3cYXvy0rn2ug3e/J+Q2FMceY/trl2Lp
YUe2sRS2KzjAukeYTO7ESihujQhpBYhYDfOCv68uXQCpEPLXOYUCXMmUwjDk3rqwpwWLs66NzE6o
WG7qA7CICch+7KpPYwNH0FGeL0Ycm+G2RVoF12oEZ0kDgZqfyyjN8a/jV0PZxHO6hoRGo5G9mqmi
VfV1mATuQlMJIMc86SKkBq4J1kXYfCK5GWoxy5LtxUZojbYGlmKt4K+8EPZZ985awh0aD7HZ0Uj6
AR+hf2pzfLKJVqNphqokUQAUEr65YAz5fA7WR8e3fSC3vZJcwIvTw8TgYtrCTQf2H5xZd3C016RA
rjtB/BQ3/aimINgssJcF4BakVawAQ9BBPru57ftpx9xIvSzVq+Kg/iYRu0ELPBEUq1/CzIeCUFdu
8TjJN1ug3JzcDFT5j9VGTJBGxhts86e05ykgab29QGU9EBHWSA0Q4D8CHuJ9shEM6BmJQOGK93Vv
JbNbjMVUXqEAA2ZXZMwxP+ZKR6/i7m1NMrFtXx2yOYHWMp2YSHTJCbz31dmXdkU8UAvd26P6smQ/
j3alK6DZjGvIR7nD7m3QuDv/IAnE06QLuiCmTvlwltGkTZxO2/tAn53HTA0vBfIE+F0N/1dklh74
hfff1wagdz0QqUfFLpInN8EENSIBJ5FRbZenE8I78kcFla5yHXYC6lVLlQJFJoNx6Yypxcx+E8qB
D6vvDcB/4sb2dF5KHTiUyyQmSZ9jqRy/5CnhhoSxLAhvQErogxD636eVEqZr0hHKwsfJUTiVpWuD
83+nTfnd9NxYuxdBeX+1y1TvEBbxDQ7sjbp2at5crtzKbj3C+ZXDmFyc0zI874assITqieJwFzbJ
JvjIOk36DPTpyYbMcoARdj87qkdX9DGdY3MAXG8GUHRi0+HiwZ/uWpZqspYtS9OZR5H8peMs2Qsa
QJ1EQvQV/KJ9E8GKAF6VOdl04Hq3dHZYo2u73J56T1hJPmKCcBkKXa7clkRqKjxF6vSSmRHwPjfQ
7zZh/VnhwFix8w45wwnM1OSLedzyA/0mK36S+UjMFTH/1QuWeMma9Dumya3CaTN1RpRCUDb1X4LN
GpK4AkonvXlCX1A4+riDmOswfVwiExJndBDZZCkZcLGtW+bOwKB4YH0KR18oChzD8djlsp6XIiXn
d8J6LhZrYucpC1sXcaeR7KDjCgHEFab8a+ICYACA60OPwkBLFGsUZ17kfyTskn8JyFoJZWZRFXTU
NOdi2LVyNNPx+FL0L9Yr0vs7bSUZFHzOiZTl8LpdzlJhz9ea4XCeLzCcltrgh1AOXz0ZmiNbgDja
NFH1S6RiG78VqzkHyF8ElHDFCOhI/zBtjPLOo4sQWSmDLwxiHu7ehhC0VsRqSHnsWddITvMpgdYk
es8zP1V4oqNeozQ/4NyomwbPF85hHNKXs/JItZr6os/wh42G/4NAcTfa0ZtX5zq01BF8BwKa6/KN
WrjFZOjxaX8+w4KzhZcuk+4W19AF0ao+l0K9Ndn3QwF5RGgkKowOXAV24HC0kUEKqelIAABUyGSj
s+PsuCUlzlj3/5Kivnd+WT39zYY6/Yz1QDmUxVSMZ+doeQxt+JNkw7ARKQzAJ/NlSf/gpbJ+guQt
fwnRar3jyWK5EtI4aW6uox81Jo0KGMHw4r0ylBKbn7sIQyvwVVLAYujG44/vpKxav9cV0d2iDf1P
f02+TTAeqeXORrqdF0+VtXtkrah2GnmzGW3A2r/o/8ikiQsQpL6vZqO3Nr6YzAGAympAFB66iLW6
2b+DACFwCM4J9cvcfXgIqJr1JnjliV5rOc911mznsdkJIJk/mF1pcv0JeEm29lZcCmPXIdFRAKEG
3jVvpFmajCg2VNobtm4+WUxGzEmF1nUSdayqRscCMNCQ1qbsINSKfLpGYGEz9SVOGIHJ1Du8XXfm
MWpIcd7oQCtWuW72p+2ZXG/Sf4vi2LKupm+4FBdz6sYbvrM9cuTtamcl+lWklpBajGu7vXQaVi11
0PAM3zxPj7/Z8i2Bubu6bLvy6SWKYI/42iVnNSxqZMne1fIGAay17PNdoMGybMW0G9dxSerArLVT
fn3cmrXG4iGfL4SSehWhDTF2CHSBsHvFIcmIwnUhIaMNA1LQ1WpMIgHPRRNEZkGjDbCgw62vYA20
/m4Q8eFexMY0RRIm2pZ6qzcsH3eAPxOm3i4nG1MeGrFfkJZrfZHvzjk3SqCmqHV3pRYgLTTeWnHG
+nnaDal8nkcsOJ/XcqdNkVTSWt1QgQbJI1KnP9zKWHRkmsAYLkQPjeGqN/mmtP+eBCFuSGl+1fTx
Wy+EHuU8Ch4gkYcLXCDRCdRj9bV2VHgAGPUPRhoEXXGxWpRozI9cLaCrUjnf1k8ok9uTZMaoo5Za
srp4BcutvmWo8MYE/zOuSTpEaaSyLdhi3PcLxiO+CIdxNLUT7egIBXpuMb0YLwebhpdeJzyUUIkM
vuRk5MpASqCx8X80zrYaGXhgPtLRljEF4Kb3Nc2C1xErumJlsOwY0hPl4muHc1ua6hV3N8LkEnoj
YwD5jSlqqfO1pC7vxxMNgtdCzQ5MWSD+IWYKtFtdlggc0gUECnM5k9yFTznJa70FsbhHAi3qSv37
0SGc7POKI6a8y9eopVnQ5V/X8IaDzxPUsVxYE1gJG3+8Orxz45vSntMhbLgfwTuBArJGKtbCJjCG
2ogVXHw6WB+sTIPDfEgVMsE/OkjO5Z8Yv0Kmsjsl1LZmpYB6dry1Zta1Ln0opblOXx46fCEE672U
RTym0mdGhV1u4ElIHNrMRkYUivOPQcOUM4ZX1JB8zsM3Oh5eSiHuzDid6WDIbi9mPcWrnUQuWZ5u
Lt6kn+1jVsd03ru2SD/ZCJ8TTEsIlLhe3BAuef4nAlWVVKvn0eIp4eqH4e6zhd5W4SKq8sG4zIKt
HN0DVOWnv8zpBhWASsXYDkNdLy24hUbxPirgmP4uOkVAnzaBwSxAfTbvLHGnzcKdgp/auSmvrzwi
4FXH6IcHvDukfH8+DE329bV1v6CnE6QaaMQMXeQvIDknUrovAFipGbaXV6NWc1jU6napaqLV5Z40
TRqlIJsP7idNUDEAglRX/0rANKDL3giLaLBbK/Gat1uS6zqTMsjFKShsUlozyMkKf/qsGr18a1ZA
lcAVw/h9WZ8E0Ep76scGAXmvg/5c3LWWxKS3EJUuwIa9XjG6jOKYUIAcpf9++OXVcHDCkxitklZ+
pdhaSR03bxHjA6gF0noGPajlHZX96kFc/1Ak6fgsXeT7WDiIzvgwsODtHIZqRcTjqQehTPgzauoa
Cc7pXn9+Tmz7HoGDuWXaR+h70obSxKg2jQBD10WpBcajteL+3lt81elvNqCk+zo4DCjoFz2Ol6nB
chyMFc19lev185Z2XEXtW/eQYpJLJtzc3LpsmZgczrUJH0enF7bNVawxMSAlP/EtSvkzwEvaj/eA
QRqj69scrG3ej/Vmcr/0KM51HI1Ov91TpIGGiDmz7F+CrIejhwadOBWd4UMdY64FHwSslMZBeAhC
j28P34humR5YZiGb2Oh+OUTUyyOvSnTzpF3oTP/AQ+5SoBlec9T+pYgmOXmQYTy7N7XTrB41sL6+
HKf3TjlQPilrmn9NV8I918rByh5AWySKwPV+hVnDD49ovhRnyK+gAkTF0ldWUFM/Hwto5+lzzIhH
t+ZP5w2Gbd1KTH2DDoVFS+vYkN61DUCq7cdcgq815HFMVo7nwG384LoigonsMxLljjVdT0gOGmhe
pEPQFQBhUK1+0JMHzKEfRgCjCovnPJzS6eas5l18zq3jcgKpheETb2e0xz6IIOIOnVQXytwHOHAQ
j0wwMKfALxL7Oy7V2Xr1j4AOoStFQnw3uTzKSspzuNVZdRYVzI0bzygBrasP84ADOBMMRcz+9neT
SHKraqWm51FYex6s7nA+vwCgEntDCn+tjLy2w0YG+Smtkj86Kg7j2CV+P5XeihMcxZZVmRQi2meZ
vVYo51t5j5QGlSoebpLirXxwJxTYtOtmPaj0ybKoCe2waEiggz1IDdj14+ONJaH6UB7bOkxtzhej
0e8ZDqE5p83JrCNg7YWTTrP0HlnxyWKkiZIKreQMKdu5gJnbdHJRkKNTLAA8UlBXOdGWOyGiNG6Z
qSb/eRfJ3K7VZh2JGaNIKABqE+trrfAhNIPuClb3xlI90IU9nQ711PAtbLPAsSSDYcjnIZPDIc+L
KNfjmPW7sBPpTQarpoDERPJ3QHOFFgtf9zQDpUX4Tj0sF5zmYy8dGZ/sbCKMVtEohXRMJuRhPg0o
SoMqsH0ao7ocM000cmhjvyW3kPDVeHGgJO8EdFAEdkOYQcFTfL31a1k6o9maAUnMjK9q7icdRjXc
bBxdvAmuW619zb9bgdRraOs+0v+9tIkI7X7AXf2DisTGW+waJKGuODmC9mbJkKNA3lpGl42hGYJK
rnke3OTyLAjOxxRcg5avo9d3cmAs08d6G0DzSNkEihPL4VbrRuUMgX6Id10k+QRWuHTZ83U1hAsh
o2aTlmTvvrgrJocyI/fHgAkySnFo6UTY0+qN1YkDtP6X7B/oCwVdHCn70iCzzuRsPeWYy7aNAYXU
9pPlQsf8Z9Jkcya6LWzG8MixkDLbovfPfbHGkk7Z2ovhD2pi93eR+R8dQsQcvwXqiUuJnZxZxQOu
mAFFs2QRDcl0pA7/p8ZMSvr1SDKAmcrDIlNpOKf8mYD21GebkLEFiWlk2QsGdKSDRFSXiGCqWGUm
cUawWAbqWYit0s9a5x1NKI9SoMQwATxU+eNiBI+CqshuQqD8wTqEuZejh+2v3PoMNHZrJP66eB1I
TiOIrccd+F+P57jXa4dFRqgCBULQj6nhkqvLMWPWM/7/7X3Bl+fp/GlR/uVxpmOSAS9LTtZj3Yk8
YuowbNRQUIgV6n1GZ0hBnLbj4Ped9FfTNU0JhpuOpFtaZt0QVSrHuJoIJyy0IKU2u9yS1SFeasgv
4gNpxLHrzSTikImm7Wv+oO083OWPnOotdYPmhGsXw9h6TLUuozg1RJzxxayIVG/+rj53b1YQHRW9
2NqjMfNTp6YDDOOAJScTH4oj7VI2J2NnuHdxgTcnWYmUUSyMvVcSBCf96h+2ek3VvzwYgllSK7d5
PoaciCRLmGhyz8UIhzEyUeF8PSwK8LX4tcc2sgo7Vsmo11PU1C2OZuO9t0g0wja2863ribHNByxc
0EnZ/hNkjnqvvVNtvKvyxsyaDu9wrDm7rXjrTtePpZYEIgsA9njceiEUwyBSMFocpPw5e7Vmfgr6
lk8vsmBXJrzwrx4BcLLm52guLXuXv9EC/vsNFUQI7OShbFGa679brTlluEAyP2mnAUphXuqvOpR0
ZMRGnPFfHrdgRHuVJylJ8EI0bdz2CYnNZqDRquwftkzsygTVUq9gBnk8YrPxA3+uveyhqCBldGjo
m103hAyn9eoEK8+0lWndOL2pSVmo6FEjPvWrl7RgWJhqg70LRie3UwSrIomLJAdjmjmJNvK18Q4o
Lhv+2sSh20rIbEl0xrFHkJmZ7NflFkSf4pDcZWky0VDor+XNJo204LicsJ99tW49+HFCVjSBUaC2
4nX+VBMG3AeXfPbnAE7oPdCuy+3L112FFd6Xu5QbUIe4rv1rFfXagmkyQ6gdYmie2dP+ZSd451dE
vgRazjqqrQl5Wo2SEUmko7rNdr2rWw5smxaB87VQuOvhb0qxzHi7OZhWELVWD+rPiZNc5rJ1Oadn
49cwNS1vKwLMwfOMCaqssEGncSzg0p6n8ewjttILY14fZIfNIZoCfV4jDxUTXmQUs4I2T8Y9DmSp
U4XfG5Y8F7cCz2ZfHk20aWrwzEWNizFLUfgnSYax0AZbZqz7xaj3U9DRGV1BH+rBM4dPjc+nJuVN
T3aPqNZRfr0mSWYFK4YL1+wHr1tfZza/yj2Iz2y54yRTA1z/ZxgSFcyPKVn1U0/7vEOqSroIJdzb
23YydE0mue7vNe27FRnFhyLcR3+SfsgNTwW/o9A+QjvEDQMd7gT2oIDPUR0BxBBVfIOoLG73T7+j
rhr5XEpDuv/vQ0pF7t+2aAT7kk22hZc2BNyO1/ytM9Mj99G+FHO3zVf25hDhTaI2ZOwLgBYJaR35
S1rqRY9+50LiBFcM4uEf7d67Ty6Y3pobcC/AbGspWxG6iM4Ieiow9Zp/UtCbcz+tdB+5sO96fJCn
sdFEL1E0IbASI0QZgHG92lck/nqNM9IQYZDdx5AIXWdqkvI6Rp/0+nuOXPI19FmLJ+WXEJXQ6c++
QfH5zLVpsvx4kY686ryoHeNfO0exxOIpLddgJoWAlWE7DeeZgZOdXC7iHyT934YTDGGLlSmQusod
ahCX2KJLORcjmg66+CH8wgNbl/+CPb5YkWz7RwMnWWDFrUUNnUmwpUQmedDRNFfLWygEImtkH7Ho
R0MBoC8zJ/eDCGQGoPOzlCssD4F8ZmLAly4psteXNHDY5mOCb/P8b7Qd9tyDSr8jnn9NkAa6Udia
gFM0utq46pv8SlkoaBfJJWN7FmbWZVnLrF4HQOB2c7msUnZHEYzbmaqofN28R+C7LiluKhQCIAb6
Z1UwZTVzEsOzHFAAZwfrwiLZvJgC3kv7gCzcSeYDF6SZOoRqE78+QuIqcabs3LB1Q6cZoSC3MeNy
8JZGgMnYDGzfj7GFnnh4G7CL5S/rJ26/7hYFrYryggnmjBvaMSTrkiYCrtgQTW4IhgLw4/xDI1j+
IIAetDP15LE8uBO95eRrO74O2OlvGgIk8PYa2UfK+H2qjW4kh6Ox3orwGzEhkXUc0HiWmTKo5obW
wpgzuxYlfxM3u2ZBoewQ5EBQzxFkahdOBIoXaXbzdspV8wRvZKNkLkLvJPCKgC/LkluGYzYmt0um
fCbNmv3Liip/JKD2GKXW8k/PLVKsor4AuTfVj8t1RhMI75tV15SAXVSzC3ltTiBXnPf6oIzV4ZYj
ddq3K26kwijhe2xGoposb/IMqOEUQIoVN4oOXZZ8mUtlDRInkdfNnuSt8RwgFoH3UssXcyxac6U+
xGDx9mze9RKZn4H1fMFZ1iFcFn0K3qbfmzzbwtlYJf+VKt1UmuRgH1I2W+HuZiEQOlXSCrX0ftHr
6ewjSFcLDNZR5t2CGR2/KxXrr8P+Ehh1us6kro29CserY5g1R7YtK+tYtCOvTjRgZdRkxiTRQhMz
fhv0NJuC00ao+BJQhRRcohn244+ZwuAmTrrLqDKsRPw9D6FvkUCCHIx6apiuYmXDL+SpVzB1GSIZ
PJfCAn387n2a3W40nHYzWPT9GrG0J9W5SbP1i17xTv1D9Q10SdtepUzIsIB9kAaEv+5mtHyTBC36
9BznchooO8Cq5Q0yRk6rUK5ZSrvtwOIx7jCJ6hg3BfMkRvKfrOSpb9vPZck5NhuDD6SgSyGguo1F
wtgm2ZabfIUkhSibf2cL/uMofoqivx6fqUGccIuqAQb7rlEKrSLw9gyOL51E0W9zfw01FJk8jFl5
cmWYD3dB4jB9OO5IdcaK3u3H3M4cjQprS94LRl8Bjx7dQvzS1LTvW4MkEswgogYL5Xy5zujzOAPI
SV0gytVSUkyJ9rVkB8KPXxTS3sV8opuDWjaVMw+tfUIORMTqgjlWeLxLOgFMAKbf3joGWUqnim1q
G7F/cW+xcMC5zSu/1V0PcwcVE7RF6gOTUaCFWV12Nh9K0+NrlO2zQWQ6y0JQdrkdrt3PlvRsRWEc
GmEtEM1iBfihtEWHYYBUzMYe0YbxGdFJuo+8c6FTzE1OFuH4iAp1NONR4MGXRe/6Q1xYo1Ciqbg4
u1WDqr3+kYvCsWXTJeInWJGHWPkDuCIc2MgX7+1hafiQga/lKbNSksetlepAaEx5kX2Vc2q/DM/P
YzsSm9aT9VjtWjz6x4OowliImGtkC7zt0nXC/HhXx8P/MpJFvUpSXjn6TlmaOxUYWxYzJOrarsXC
LEz3WryPAFxs04q2BSsQCgt8AklrY2jzLqNPAfhuLAk3w2Qta56aim6fPNrfwqoIWu9nn590l/PC
5glAKqhp1Lqfk1hcoOv4r7SEDf1Z53thhOb4b6Asgvk2Z4J8RQWuiVup67CHgVSjHIXtzIdeHGxi
/yZ0mCvsK9sqRuGbf4BjoHaE1v++Da+TtgieT4fXwpZPuV+YboIBwQuV0YzFkTN7xTHwettDLMpU
PTIZIzChc8/qsbSN8v59Ymj8ARYjnFuhWRkdR731dhrdv7NI61pV3/vChJESBewAdISXTbM7NQ86
Afjpe/aLjMMlVcEVRhVQ8KffWz9QgBv9Vrfwepm63PZRpx+hPfEAdwgbPX8HVdGD2ykF0pCAatwF
6o1f296vAqkPqktypnJF1rO0a/heYg3AilRqmXmXcPC51o3ZQhVdY9YiNGsZXWFOgmmQZPJVS0CR
UqY3or+rL87kWwCSyptFkNYvs8f4epTnhKDXZz9zlYojKFxkenmgMz2XVs4+oW17Y4TQ4CBuazLE
cGT8RJglkorIxe+faRgg5Jj2KwTKkuvdDz44HN1joDWz8LZrkAhqtp7zH7JEFb8rrYB+0c7Zsv8Z
j651MqbsXPNPomR22w811yN+lY73kNdgF4LD/9SirItFXnCdQZre1EwBa2L1G5UGJoMDeVpdiRt2
uhgIQ82DkTsDA/ZfgdEELemKsQ4HKP1UbnNY2o/MG1viMcsOwMRi+L/ypYUgrTLmHfjJjZRfCaPx
kjkWjz3JXlC4+4yKVyrPelNZufIxz1kU/zDzkOM04Wd+2NzExqf40+OSH/MMgwh6o+KEffcy1BfM
vuqRBNwWr51DkZOfx7jxPyasQQyrIar2vaDMw0W4kJXJG2m7/e4BKR6YI/628Gs00NmFpiNGpGXL
YO+TVQqgzm/NsHyekTW+3nHt85tddPJnFPkgEwv8IRW5wqyR/UAdzEMFThOB648TLWx1ZePMNDR4
wzBZ7Y+qRiVZLBtmDWWqwISg/W3fbMAcPyKEDNxFq2liIC/4emaNv037aKr9VEnFhpRFWwf2nWZZ
FNiALV4xPFfXgoFQvW5T8goqbKykGZE31iUUBWQ+pWH3V6ndyCrDz1lK1DnBAlGq3EP0DkRpOZtS
hbrwPG0b/y4ZG5PPhZnd8T6lUlcMxXhZqBrdGZdSdtIqc+PcKxOEyR3xS/ECl95GSaGP1QQ+RH/O
lKoouOvfB8JhBIJPlg9qECvsB+8ETFlSDLiUKby0e/RfCDznQGxFyI1fo9UzLwYLwRGw2iQesPqb
doDNlg+mzqNMkC7TupXF942R/n6FjDaMn8j5N3CDFdmAXMal7eeJ4dQJQl/kXIWTIZBtjdmuWkoa
YmY4Du/BLFbGJoGhbeVK4j/6+w278M0RwkREQ2IID1IMfWRdNzhzQXN9oI36XVwNvGPngG2KD62+
4qnJwuo061icjLLeDyTHZ2fdrrhR1KwTgzEFY0cQ/mERcStlD/CEFpvGs3aK2nqTR+E+hC8slV8x
Rvnxgf9b9uwwStc4M2GsF3h2V+K/E1pC5Pkgm/NNYNsXtylhMqRgjU2FNOAKgffUGvpELuAQRXva
z/+LzpeEeXwG+fKTDuOJdQXX/h+N4pXf5sCFvRued3P086apWPQZKlLL+yM0XEKJDFpLSf72ZxE0
fiEm1Xy6I9VYIEyUXmL1MZ5ZeuBCg4smpU04Jo3WTpevWhjwDQxj1MLYESbpQ92UeWh623vHURYo
9EvFHWEjH40mhiBMWHv08VE06SRXrGkDHJlIs3UbjEWmRIZUsSy0vei3bdJW/TKlvgW3BSykkhm1
lxv+VICDKZFG4KETpIWeDg0zzF2VVaiF3bdKMBP7ntMz2/N0mLSGgkGNGza5xhTVrTCl9v4Hcq6p
pbuFgy6EhpmHmrR5QSiuDy2N/jX34pB/YDNwGmztUw9871YeZUb0Dc5k0HDrQCKmfnpbdbflLJDu
k7AdB9J3dJwZHiwxId+TEbSBkmj5QZIygjBg+5/LRcBEekFhT0O5XtnbGr+rFN4RHQhVbWPMAFtR
hkDcTBsAFkCdaT0XJDdG5+j89oNLAtTb3rqF6UFpeZDJF7QDwnl9mNkKx6LARQvqvEszqHn4SJ3m
dext34BOB6S3L7myXB+YjszOzHoOzOpnC14fx5nggSvVgDavD+E6Z+DMaIMP5NMJ59GgA0xmUGs3
xAfGgiyhRMWi6csKzbpWi0a4sp4Q7f1IzC4obs0yoq6KdsGQti3Uuoz33s7ERsBgJS7/RPccrqzL
I5XnUMrXt/8LvG6X/bZebVZeGVHs3I9v0BOehMRc4Z+yAG6LwfdoCZb38qeQah1Irzj1/WeiVa4E
rnyfbpLIUuISbiB4CX8JGEy0Kr5OvSJxCOVLEqWKZZB1IXb4iz3V4h3gJqu+I4QCOyaVT3o7RYZI
tS2lKtYQKaiOlSpp3PlPHCFi17w8cKxjnG9uboCcl2VVno7IFN/R5Ms5fI0tKZQcTW5RKJRL6nd1
+7yLT47YgparuDdS0kOmk3CjM0YMgGL/ELHdHVrZuEcDp1JyYHlqfI2u/ANGCseq3pNAG5kVZlNj
fNsR0KQAkBcCA4UxI9jkQYbkVzYwW7zbOD6x+dXbFXWrYxiZnaTDZToZtOfpVK9gzApXM8X5db0c
K0wGmzTriYQ0kuqKeM7DlWuihQ/SkybUkYKYMRd2/BTiUctd48VqNFLyPg9BXFZRZaHkCMKibwOV
xjyo5RH9MWWjy6ZyLE5hE0mhYL4ZTJJLvdIg8ltnyyLNkhhIRKQK36AZ3f5yBUHdelEiAoY5rfvw
XfvOX7FgiPaLR+P11ZOb0ijLC0gqJ7AgTGgJ0Gzarqkf+flakj93qALZ/Ve4MEaVyD/7ggB4Z4D7
QOAHzNcRpWbg43jjJ+C0d3mZo1Gs02hdlBUlplZeh3rgYp1qBWIzpjjdxd5suqS74uHS93DkKtGo
HhSavO6otwyEl9xSKciaZeGfv2pYnSwdzgJ2k7+puoR2waVvQ7e//LYpERUMqLIvApH3dkBiaCdt
VMxIqAp4OEO71y7DjiH8XUKRtrAljUpc2SpKV85s72z9igGLI+lu83ACWeYsmDAS1xy0raBm3gft
WSFJu4CQdqQXP7B2Bkmq7u2nwmeZ2hWmzzh6+dcilPlNgy/M8V6tyV9aGz1BDjsp2tcNZW2P5aRT
xeop7uyRjBTLiyJf7TVmzN8BDeUz+XxB30PuC8xmWRt2Ye2LjkdlJKZ9HLGWkbZ4mX8w64LBSJX4
4FdBdyMAucn0quPj9mfOcrIl8bs98Ey3FXdRYiEk2SusNZBysa186SpNjF54e2lZqdfE51ftWkIC
PJ8hiuNxQh99bqNV7j+qYHOqJEJ8AyfDlISGrUykREsqqFh2OIcml/bey0PReYBMIFPKpFMZPLay
GIqFZYX+jURmStq+il6fr6WThP5yyKLGIK0AAXRrt30dixMStpQX6DDLrRZHYipfa0XIo0BW2h03
TRZK0qVsDQvYIrHZqqPywMeDVPlrpahPTZy39A8YklaTRBW+J8VOmdLjfIIOmBFFZ2n9JsESOf3h
bKVf9xhXjOTigIxEvvCsIaG4Y7U7KgXHquelzSSAM3Jkvl7RZHaveWYd91wKJhwueHoJIlE/LqzT
AS+G0/OFVnhkh3kUHx0wW+HCfwSB7HhFev3yhIhJ8/TYihzPQlwaotcZA67DY+slgnHR6RkRfjy4
KzIErYnL3cPkUIRjPF+DXeRn3eFXtygxFMhGzHzOrINCJQmag9TXAyS+Zbxt+FaWCFPr2kkuCz0f
/FQlf+nTrTNWaQwKU0e6gCP1crg2Cqd2Wf5Siaqi/hFW/tvyw52etErLPTZ5QRfSmi4uV+KeUDI+
crMQstTzCOHKUfnBSMa+OI8SPK1yYyjlobn4ok7k7JG4mPq7YtLQB1RaDTKPeGk+fnU0rRPb4ZLJ
SU0N8i2HEdpaVlXOTmsYbuGeSz5T0nv0wdWe3U2RUeCCeENJNKiShvyzzzXhBMUYQbS6963jJkJO
bICipi1l0MPMt4oJsa0qtMXvYQ2ytlqsuBC6vK0wJIgmw9R71ShTZ2viNdO9qKvln/bMRCb9Sy8D
O76+xDAZ0IZS1AXsAyl7HOVd1tHCXFwTLc39cuvr7cEKR3FBVTqlEDabgLv1AZtlXUnnw4i7QCeT
h1AChtzdC5WvsB7VO6hOiAVkL2yyu1xPs/b3yZeDX+NO7Wf6OUkTfu9AQ17YQexmcbFxFk9eXoti
0llHDIUkn5UASlpdY1R2fGZqA931tmZpeHZa8wthHpIl8LZ9n92F99LWtVaYWhmKYja2qGNaKPpn
OtnhvI4sEQ46yYJdA3hJD0dlOUwMkOYMKNzpd5+ilalUowlwXN9FyNqsbDm5r8KE11CyQKfgU/xf
pInZlzaGybwOfCn31crYTV0MdEkIR+miiw8ciQrGVqGUQHGs2tnhN3CpLgwuGLGFAgAOfb1GGyMJ
n0AcL8kAQ/qERNeu4do28TUqWcAaN1fcFHIqdPuE9u6zgxxnYiUCCVtX6nDbxtq4xJJA7Wf8W9qI
Lp9nlSc1SdaRmdO/YVv7wvWOoCjXKEekAD3r/9k1AOQTy7WRs4wRI60rWoCtatkKgSZ9IddhYIjU
096U/1S0jXLe+VxkYtlakxgSELZI5LWSEHMJNYGI49snGKFRvy4jSiufHEwhQDLoV9B++Qm7L0ob
C4RXyPb7RWjAfkk+MWj5ybjGF4iz48Ihi5ffaAQW8KUioUvQPwzC2Kn7LGXAMN0Fi5VUSqYGHwmk
etpbvkPtgrLPpWP7yh/nV2QzTaI1pXF2N1IgcMawhgdsgXr1mEhu9IViPjT8mz8kYkXQABjz2xtg
5rITXP6VUENfFhjVIxgG7IsUORND0P2X8jrA8joL6Ri8IUBuK4KABVdgzva/pWC0Y6o2mpUnk94n
prsh3DY51q7t4O9x4QBKI/L+pUVpAw1tBSxkJriokJ0T6K4n0oJx9AxK75UB9RCtLWcFarxlSoq+
obBWlmE0pLpBGkorAp28Or1gdHXqQF6AffgFqGpyJoLxwJfPy6QHOzyTRehwOILHlP+G/rRz05iU
S/NwZCsLpES3PcZx0h4FZk0/r61gas7dS7hIY1UQVgX8mGbmcvcGkEaRizIEC/Z3ZctoSiBm5DfB
u7AvGwShSmXz6QGDYXIAsZyAPN9xljboc7KC1lSh9YS8D/R88ILWUp6EwJdrTO4ZP3ZcCtQ6UDn8
3IFWbFI9Ek5GIeVlm/ue0sLKv3aPJOroVFdVGAJr7pcsqGxCy/s0sXwIxBvJhpy+ra5lGf00OtLt
eJ0BRCVn6IriWoBJEHb+83d7LYj1XxgLtZ06JvzVeyGMCGYTg7NMGsqlnN/Wj/tC2MBE8/9G3z3I
StPl1n8QxIjLVAH7a886/fhxrNeRCJFw4Yjf+aSuOm/94j0+lDOlhpEFOuXZSe8ROqM1lg+Z7Og9
FgoMlrmpzKswq0IwSslqI5+yLw/CpFnAH1yrl88nscmruS1JOb/gOoFhPBsIvq37lJRGNDLmhzmz
Ovoqa+hMypQp0XatkMyKdFLuAkROR7vPPvFoOSApRrv49R5Y6BCvRqVovFQRLT1D/ot/dIgeoftR
upTCDaRdtyEmKFdG9IEdHrSYJ9oMRBcvGxeX20+MlX6i7pv761qLmRFyyp10OSl8rdAZZgCEVdMz
2RiK0VAtJCHGDSsGGKME3iLZ/nR0GvQJgTx/qkjyaMkC5gWYyqydN3JtjulUQBtx62RSZ1cf3zim
uTD6OeCFld0jpxkeUqVzygGMCaGDSDP/oST6WkVCQYGQkuitxtXt2eF9aHvbbVDPhuA/yd92eMcX
/LIo2mNlX+EAqSJXxMZqTpbR5QjddCFvGnhEq+1F6wfQHI/EjK4DTh//A0EmN7eiUvYdNd8x5ptu
xRbyMmeQa6ke9qOVxNk6BdY8CMqXnZUbr+Kxr8J9VYHxOSlX/RpZeC9oYIZzVgxUVnSA37aZ29Ez
wb9s7f4CgcKfOx401YUPeIE9Ju6kWNZAKDJnbEDJhreQObiVfwOMalRqHQtcraKW9S8gdLOeNcxa
HuJIrjXDDzJ8iF1LkXK+T8Al8xMqIMPhcnQK//1SCpYi+5TeZPxMkRmcCK0PkHRYsnB3GdB6LswF
iBoNxVmJoCuQD+x+ogbZDc1udUUEhw+VLdM6HXHLTXjBlvRsmqAvG5MHtOAUEB0SmCYUlUFPttCp
ZqPIzvYvQf9VFS35/8dUNHBnUK83VWbxgR7nNkKOHu+/3wz8VMh0BAwmV8N3/YrKy26f9AGU5F+i
l0heIV1/AoFbvUQbKUOZBgnaFOJ6TIEYd3fPuqPc3+1DcQKPiwnYiAK8nkhJaugcd3TYHwX0pM+h
spYZ7HysDjmzi1xH8HPFaiXL86ZyfpgqWqcLXGBPcV3/9Zu8jF23WO8xbsB7cfskfDPcb3wZdjFg
MEF90UHd3vKgIK44WBiOPNBjijbaYe/KZwC++jioWbztZA4QmYKa6uHfyEv40bZ6sdfrD6IsAnY3
xVt6E8cfsDESNIj2sbqtccoEOWBwXDm8GQbC3hdX6IYUDch7Rqku8uGfbKHqY05E9guuCeJKhUuV
HWqOlzW1iuHuhEnYg7XHRdGy5FYqXRBnl+IEoWvY9x5deaTIL07Dh5kBGzDGABbIy39KPnwtSFkh
BiUo1pgp8S5VOcLEczWY4K32neSOxoe9aqp50cd+yRU2UsraYYZrGYfu3ws7g7UK9PXuvne5Avak
+UEDG6Pzi161Jo2Q6dsuBDu4k9OBPmCxBW6kYelh3nkE2m46qfskuKm4a2YiBHI04r7qF7qbn7xn
hGx845dG3mWDF8Af1pwaaNRUwlYXl5qtMQKKKjloBjJ9xmbSUvtLwrgvdi5hGi3XZBGbnE92Kd4q
tLgW80aMZwBHrltu5DXr59k1GnN0DxVhYsdIIAzjAlEs8yw4lMsmVrv28HftymZj7sUrJwr7j+hb
1r+NiaS+ZY3QO5Eb1ILx/d9ayMhogChslRBhEKqeoreBJvq2aRo0nziyNPSZUb7olLaINxNUc8/j
ECibpZGfV18pbeEt9LvHuCLXXIMO6tySGrMD13zeiyhUzWsBTgluI/RDhCCDbnUwXYPQ87mBsVYQ
UfdJrLLrxmJpDIMNsRXWjFid8zSsGk4Z0uDAZqxtQPXsM0Oua5/rbJKr1nAEXbWZgaESJ5Hptd3x
Uvn46lTV3/zvGxNfEUzAkE+2cIodrHw3hgqMBJ0k4I452YI7UR+N8eGgHWqZG+kjzxniWfPqu9hc
IK0CDnb4/qFuri7r7rPo+Dv+MXRpArUfM+B9YfsWKVO48wkebJSPei83xiAx+1xpFjnAslPWPSan
1zckEGIwsBcS3Tcozp25jzCIjmf8hF7zDc9BFfbMo8s9OZBc+OkVxvNngjx+5Rl3jEGnGCR18tY7
rlh8iAPAZP/wh6HNh0dOpv4uSNe91dx24xjoyxvz08gelZa+tyCHgjFrXEx4FBYt4zknproO4Tpl
zkLgC5ZeHMpvVtXg08WwyJJSNOrsHz56b1l4mD+STa5ExdSvvVPX9lTEOG3D4uhmwjAYDFtj8atQ
y+eVG5qORms5vuT/96/2oprohHVJ2xdwlK3vS8R4eoZoMADyH322dhjCAdfIsNZDF+0IhtOJXIQJ
jsGndbri7rSmXqNA9//FSB9OwE+5eLATkuXanWAO0h3lvRfCqlyjcTMUPcgoQDgeo5jRAYURoN2D
G+Jv7aiAZOUjK05k3sT10KpIBeMo74ko4Dp48a9xVD2mWqR//h9JiUhByA8TiY1P5cKhFPwXDqKW
QHQVwyzLF5ZGKt+gKUkTwz9dPYnRDUeLhAKz1Z/iMP1WghyRtPC50oqSY1niEOK4YeoiAc/JLlZ7
+37irHop6BZWWrgUidIKSzodTWqLhQgAKTLJr2fzufefgZGux+EZAcmFaP4+M6DYPF1XfI6oh3Fe
E5ZcCPAPvl9iyLTUxwcMKlAwL9Efa5xobkLaxezf554VPx1RyyLVy/GOQoxG9sc+2IC6tPJ/PVUL
EMqGlONxBMJCCIAtlSgpYwHFo6BXygPb0JFPZb9i+RlafbkguXil1WYkXoTUKFPO8ROg/D343zqY
8KrEqpJ9NWWrNS62VVtoLN+Tm+VMywXo3XdE+k16QQokPKEKbbz66tVAKZUeIBmFCwAtGPiHpgdS
CBWHpHcfoxG4YjuvjxGlqti8jclXx4dFXsROiFnkwG/2gsHy3omsNF3ckUOQk8Mzz7x8dZj0TYAk
Df12ySL5Gb03UWhafLeR4CWzrhubbmd20WKiZGtTv1WMx9KamZ78i6tJS6eMCGiLBBTyIvibbMCS
PgNiUVsAXMagnCMr80KpHX2EQiNbLu3AGyI0pXlmcBhda75Hnl/r+El0jiaIYjeY1MP7pNNN6n7W
VloO7gVwcfDdQj3GVJX1mWBgAssoVAflzeR5Pgfj9r5ap1yZOQOzdFmP2HH7JQqO8TWobj3IKgxV
BzTEzLKUWMXErpSKdS4IaoenDAAFxPZZ3BW3GV1tEPiNlN99LPUK1TKknoQZg8eK/GOsSdX6xEZe
AsMAcgHW/5qLiaHKhC0VRzAxL2UdrpmW5+sEPLuyRn85qhzquhZ0FeHIvYM1E4dcJQi8iaRwUfhq
c3qxka154+0xshAtUoVPxenc8DVj0GenbUe1AZJLp4UUz8BSQegEUQOI0R1LorYaRqTAdS0xuQ8R
HCUBVY7SdqirMqHmovAjQI+K7tjCOn/Nd0xKAzWw7ct7tTpf3tsMKHykXb3LIVI7IXGCsIpZ39PS
iZJNLwYSjGyRCqHFaMWUGHmkpF8ouv1FcqvILD3m46U6KQdlVOYM8AOt3Y1Mjl8WHbEWza58/FXL
4rNqKqeGgBjYRrjuRhzSQO/cMtTXYxNrrR85Z5kVeD2TT7TKvlTIOOlpu7Dut56NUNuBCiHZ/RnU
kcAt1oacPEeFfk/fsTtVqo8YdRS1OTAQGB3wnvYH7Dm0Lnk07kbwM8GIc0hOdjW/1w2tc8+P48l6
tmWDzo3WdsHd2dN43UWvhZKvydy+ZEJeSeKy5+vfJN5fGLUnc1PrpEqcyeXldVOcFk7MbH76FsS9
rSTAN7VwOiIHw8dVQbFSpcb+LoFEGLIZHgQKwjRM7zrUXwLVbk4++HNOgDzopVPYV7gKS0KlI8nm
S2c51ifUqlwD2JM1bVcCFz4FEfMgJrh6NPAdTvPgqQZ8i98A5KhNQ2kDsEJ/dn1d2ln1oZr07Yfh
NlyhYVdIAZitPVbRTlQuzL/0shGwnNyaFBLCe3Qcjo7CCQLpEy/2u+LpQ3Kdos9+S5zhuHfmInst
FRGdSXSThJvy3X2qPZCGlrVq9KWjmQ3ltCKi5gXWzYuS00znsx1xsJjCbjEY7xJtsBknk/CJl5y1
MUirW7srRuOB4EtekQicwWaUUMuHhaDz5p7mV4xoyvC1MLM8F0lhaUIZyrAOUcJ17zsqPhFjzSyc
zaRBKcB8wX5oLicX5S3nm/V47R8blU/b0aA8Gk9GTx28AWraE2h+94JoCn+ko71SW6PNEQL3Uy1p
KI1ylBRTQnzxCGkOlmE8LylN8+BTF8JcCd4WkC/zR1huqil/DMnCblico5J2Lec0FyO3CqiS8kxv
Ecu6pl2X4I4AAjPxX3qw+Y4/+dENVRILVw7XXg19PPq/TVZ7RbiIPli+Tzh3lPA3hGUa77gxz4KI
0B40mJcvxhQTZfz/Qg5hjXHZYItf8/lNQzjK8vZ1CMazt+GxNJFUPr9qenhq95r7Nj8hyLLsIImk
MGv6t38TbwAiu0u2RYfEBN09jpkf69BL4qXmWCfOYZwpTCxLTZPsb4S2/JW3DvROrjwOxLjczU7h
G6qBmFESHgtn1jVUCCzuzDgJ6mp6A6uhdT6nml45u8mSjBU5iuTwScrxFNzFuAP6om5fnoBaZ9P4
2K5NyEJA9XSi+b9vat1f+EPl/GsMSovt6qaJCKrc09U1k4M4CB8JlNcJ+Ain9LMiX4Rk/E6NGQ3X
pasojtuUORCZfSeF21cxiJCGN1bT9OAHAV3wkAaIitOaZpBBBwrB/e9E6j+aHxDeHnlBPM4uqD2T
+wcYjHet7IxgNnbv1vlOWRboEwn8S3btbR7vWvUZ2fO0H+X1IlLpRy1A97iNNKBs7z9RuGKOOWxX
qykWHEWz0hlhjIVxlszZHTqkodJLiLR15WdySaWQjtc7fHT7Wv22tx0l8hOgGxVUxaK4qutdp/Es
yZwF7iy2x3N40nbs6DDMlDdyifrZV8vM/6Ejsmk8Jvnyt8rSkaqnzPOJlBgFW73pzR4vpU1rstfu
HP37gENhgV+VuqSQpzRJDTNrfaV65KnSw8VjAqCXSzeelg32ggUTr5w+7YyWM4kU5nkplGVswDwx
qjpB1Q3sAq5gL4ZRUc0fp3tMRxy7VBsFPmJ1fnUPLF+ASVHXaak7Ub2P2hQ90ieo/WEe8c+pKHA8
dobTPT1aoUKIuyxzsBY1E65lWy52cp9DcE+MYakosPRjKgz1rrqnFu/ScmA46BjwEIlI9QGyhDwd
jQB4QnGMfhWYdfvnhJnqIT7Le899rVZhXEFq5mbPrNMJfLb6Fj30DHVygHXCpYU4vu1vUESSoS71
8cYxVqZ6o9M6HxiuNFPqtql+J3bd9YzjwXTttUlqqEO7YtcCWtbVOSqFcyxyBJ2DTrq7gegdRcue
siQZSipFzdpdPNbJW1BrfYs4JaNiJqWYAotH3MKegF2w4lw+43eMWQgVzd2kMpu21ibPWhG4rCEV
juv9u+VLY9csIZ0+Jr5GWHct3BAu9yvYKL7+9jdFU4wO9bDhIRlcZKBBtpIdFXO5mgapiUVUYf62
rDt7DxkZWU1fGttYbajf/biSBJeRZ34SW7in4+RU8fa2PtVjU6FTUO65pPx3/WJoiQhCjkk51Pib
jnP5TOmbywPx6yWHoSIz7JSiVFws8t94f94x0noh+ulZ669QNP6Xbef5jGY9uD4wGoNo46U0VeV0
YU3OGZHmTJcaa8PL1Y1rLZezgcKBwVlcR0FHNmTiH4GSklQ8nB0Lin8w+s1CLr8YszxcKxCpyk3b
rzRLqEeNXp1SG5SOArF/k7NCt5JiL+PGfzbEjOirsHvAfWDnKOIg5bPnyBTdVyu8MLBuGwy6GG+A
0DGvZN8TGw90cmHjnfWv7f1VpjpCz2duw7I2/RYZ6nr8XOTGKJdJuqRgnwxVBG+aXj2fRp4dAYYZ
tOaUkKM08nF8cD7Ai68zzWE4cxrhsJC6L6FwqOJM+TCMluAk7wgMrmvsM3vJ8hSJnQhC+mYgI8Wm
++K5ZmIU2Akc0VYkdyojJmGlwMfsYLhFdeZIIiHenShjoNyvVu5gNgUp9I0lSeKJz4yx6W8lUngH
1q+LCmA58gbEuN6ZjSSnvX0+bKg1JPavy60ZsfPFWmbdVyQCsYjMkKIeSzJluwt0IRDNUXx5Oiu9
EwS0v8ySMRHpg60kJf+EIbeFy1eIarbfVCaLdU4ym96+40PD4QfyeUofJu0dKJ0e2LKqL63HKP+r
6OaLts1YHUJ3Si7m+H7ssiWUClrDqZo8MH6vHxhBgOLfsUO/ZVtUGnCsCt/rTxjtdqhIZvN07SVz
VCy7j5wuBCHa7oQwSbQnryC/GPNfXHyVFU6EJDmpBD5bd1Tmn4DeneFbHwIU0fKy6EjqP5e7Op4/
A36bVSht2XIu5Z2chZ7oT0IISwUaTiXGJ7FPmDs5i8dzjwabqZ9AegJ1X3ZhSEC5sImQirMnLo0N
xcOT+T4PClevVlE/4kAciW67Le4W3nn9bjxQYQs3+I8B1e+rSa+SmBTOTe2RT04rvDBieBScbVJM
n1Bk+23BNUuEMCzaMC+RhVfwWGkLtFOYyhX8ZYJ2/teRFZ0bz3IPCpj/kgL0S4cRBujMld5sxUCq
iN+dA+FEMHmOgZ8xTWYPzZDgdiFPWifUvmTUUBxYdjsE8QuFJFSoAr629uKA5zqgKQvSMwmvbhDF
/yjW41Bdo5kLwmg12KMUFgzTDkiXj/ObWu1+fvmE2RwI5dj1e3+K+2A51pcfjDx0rC10YZ+BRCcP
0aCyQ8VFwEf1gtyXpYZR8pkukrN7BjpMtvf0VzRk28PtNXn4MzQlJA7CkqAqDSqMiS0bMLfgrqFm
nrg0A5zxR21+0VTfvYz6qLIaGZC6h7sW4oVpWNqhiXQaodXxK2tZsdE65V/NehLZQ+xEW0JFGOge
+DpEnAaAxxsV4qk0Co6SO1SHy3Rhc0HjXMvEITnhz8Iisc/7jJLSnHGBaB7U263BtiUJVv1axeYn
ZPyTBZoMgPaAfN5DIMpOIIWS5JIcirzKFHcORK0xYQ+KdHtBYRYzpvCKRnEbIpu7yUmDib/aLJjM
AWkoRkXwf/OhkTwt365/xHb0WS7RdGB3Nu7RsR5Bdj52t1FyCm9wE25BpRJKg+CnhU55IsxDYfFr
Xuht1Z5VRxLZjmTwwagvI7/aO+cQLCTmqdV8vMs+ef+Wzv4z7YkOkOqwxBJBJKx58jH9rxzO/jOk
C8AoabSKDbHy6E4GR1d0T0H2GzOhdQ+l2ps0t6PCEtA7NDjNWeIDKy9jNQbXv8iQqyXvHOePC36+
LjclUxMsAiEBreCgHGkgMZ7UfPdULfOTpaC1XJztpdhdzxZf8i6x5T4vSIvkK6QLgRnJ4DrOEAuB
gsi9OFieOwZQyt+DQiWqu/SDMa/OUr2M/d3GgI7TYhiaab3fjAkJhsU6gz01DzJkwcrUIvGswJIM
6tpq8lOl5FTjoFOE/OGeylatmftvE3Mwma0N560c5JBqp6k7h9xlOUXrDGcma8AQtq+trIZiiL7X
Fbwq8P8cgbBzgGYeAu/ShoFaPbtxKmRuMfl+o6O6mq3MPD3jCCjMyltDKZPDqr6hzbkrt0PmmVBQ
gxpdK9+UjgU6ujilIeUKVVgVIBNVgNLHvkiwWunt185ZkL6Sl6DrilTQPf0r2cZSZfufsq84TRpw
VO9wCfZi/JQLZz1wLY+luQCaNEwQ3g4gWzE74001qHxMZjKg+fvDzyn5YKyqlVAU351bK+f/bHsD
VFMIounlTxv5kZut7ZCz81h0GrILmUKiQDpo54eC6LHftaKSwL5hOBfMbxs50aNllC6xMtB04YC+
TQ8VlO72O2AGR0Byv8UN4cKEM9j8v96oO8JrbsttwO85HxiKqP0XqyQG18KaX4UdxGtP8C2iP0A+
m1lZxRWHyMN96XTlnxjiC1OoIVSVTqwYlME6MHl6D/0XlHwebFJT08C02BP6XfYowcGLwWsj/1eo
T4iNuYGUdrO7Y39lzkG3hm1ik/c1iF4v1pfb7On2WICn00DQZmBv/+PQCFJcIq/rrpJR3YQw+K7s
kKhePm/5bqSCIUB0RszGhWPgzTtsXCZy5C3bsdQZSlggYDyZcBTM6mX+8ETlrQ5q9dxw1h2Bn1+/
qnDNv80aXdFW+N5Mi/DrotY0sR9HiELE4msfe0uD40U0wLqHi+GZXxUftLlrbmI2/U+m3wAuZ+Og
ra2TwNtCbCvaGheDfGoN12MpRBlpZHionJBkskh2hpzZhEvTqE+TnUvCzUGP2PXLu9vaiuXVsgi9
jrBD/Equ/jT48VLGbEMq7EcH2uVoAQ41WmjHyL8rXkVUXGfM2MGkf8lrMmNz94chEnKVd0Kg2voG
HRLlurj1z83pgR+I22HusdiQedzxXzDd+/0cPGDL9TkO8lyWTejM2Wd5PtGF+N5pcDR25JQdqQIk
wIEI0qVGg7ZpfUTsstqL/oyYn0FRqYnnsG7tP/C9xxvzVkHlu6CrLYwGHXeS2BpM+93QrtjxT01g
+dONR/QPswR1oIon8OCdXXRUHpG6uijjh0hVe+XDRdG/7UsvzhkHuqueYhRGJ/PzFE24vuawAgRk
uHnqrZg4LAWlIE4DE5YoyUXN2sTNrN/89WskKLMKAQKEjy7Tip5tCQF9TZKX3QLlCJcsZN4zc9zH
mvUmczfYYHdDrMPDQltd+YRIBbAodMP2a9tgb1PD5ZkJ9bZ3S/gUpKYW7CVNt3BaDNG3P7agdHCL
hpRwU2TEpFFGF6+N9R903yb9tyWnKX+m0F8VVZm+gKNHmbpgjq4G4vF+doF9hzlhC68kQYiWteFN
F0wPf9vXbiBbfz8FM8pUHrTUapzd1svKwaICtNbVoAC92zKxWjuKPNCJjwnreKszL33Dv3AKtdyZ
pypU7z8WraU5UU0HK7Dhb+RKsMb4blpDGqdGuqPWXz5O1p+2o3ZvYvr3rLuzguUlbOvlFC9re7ok
K5HBLWUPqfAG7Iq/MCsXviJP2VmYnx08yOr6KHb81KxD3V+INq6UquYr3oDELVJpkla4toklJ26O
rnfTd3Pv5vVrJ8hqyHdW098nUycodvEPANzcU8nT+7zYGyKxTTkGa1A1rx2dp0TqwbqQwSfNxNt9
/knR6x5BgOMlsZ1n4hr5x100B3Vy1tt7z2AsHd6PR4iWTC9KvAyo7J5ohftPamNTZfR84uodif5G
vdf15ED3dlKsnBpMoGnUlvKovKlCHDrFvKL7AGjy0yhLzS9sD2ENKXc7n5xVCtFd1zm4gbpVVGaP
tBqWyu3iM5v+4mzEDe7R7+2tZjQ5BMIvP353tdRF2WYQ2nN52v/vok4FJEoOdoCkyg7tXWu6pJVk
Nm8wnDBQEaW98lnuF/+nVanvsjEkyCludVrbXNXP53NBpHO2JvkzTmnLyHjdBxJy3KsC8wcw4hk8
f3rQ5J6CAP2Fvaq5B7dO/faYGZ3r0wDRL3EMyuUlY/k3LDCLptIv2IhGAiAhlih9UyS18iYIaxkb
IKoIskjTmR1A4eZTKpWELhU0ufXk/uXKYlChXwRfMKmLMO7W/k1MQsiHjq+htuNV9n1NJAcCjGC9
wqD/I6en/bnjFVj+tnZuZJS3DgsINgprqSyhUwCfL0btvH2gyd9k6ps4AiznvV6Ac/LPIfn2j0ff
o6m1sdeU5FunnveLNiSPA0WRCb4UbF3vE19qgHO7vZQ6VgWaXcTbZrlfwk4Gp8SUX1a32ftuytgO
pPDeAzn5ABscC+ZbLqiD2g9oARu9WfNb0BqNDs6Ccav8iBaT9d/pR7WzVTatMo4jQ680UW83Ko4U
iiidrob0Ocu6e9PirEGK4jtFdKC8ec+tjeTCLlSfFXOgfByrfIU0kMyCRqXGyDQbkhggp6Xej6IF
9HQI+rKrLwzfLZBlyq7boBIw+OQzplWj6Uju65HV9EkDCi8ICBIF4zENFXN385bHaCEUZw+Nd2uF
7sn0bX6KqqVk2KFVIAn/YXBibMv5xep6/srrilANT6XQ6P25l8/KXbqw28QF8PESzYgGHzYEtOhq
0a9TwOytR/yveSWqmWMj8UnoNthfy8fBgKiufQnR0UZcztEFdPI8vR7kyn8E4SgpPcjD/HQffXLk
hJwZvglxgzsZpp74/Tluee6oanN23ouoZ5gbStxwpYc5Y2EpdNdNqpzy/yy138txZneSywD6W41N
Xi/WgqUoRpHBg4uB4aNNoRDcrpm8MBwM9yrIr7r9tpUYTjOcx1fynvN3+XHYKaAHOusPioYN9/oF
rdNxxgJghgqJtTs6TDuo3nxvZQwb/CWq3XzW1xBgyxvCGDq7tFjfDwpNuWPj73B3Lz1/LF+kJIZg
XCyymO3xoBWAw2Lcqiwbkm8mM8ZISR8R3YhdOBBA4J5kHCS6YQ8CIkaTy6FyZ7xnBQTKynbkgB/J
cqGFev80EcVSkcbMli4QCGQ91KnMzUPTUemBFXrmiqKMc+cZKNs2XjX6Q1oNnvN1FefaAFHoJNja
1okQsmrmpUIyJPr/ULovBkwZn8+y1ClP/YtaORBk0laeBW/+yeuwEtlxln4lpptqTCpt0UBFpiGp
3qzFkiBLbZ6EzpYTK0vpFjl9jbPQ8mbMmKF2ak07qvkAiXxXZBSbcbnckPzYbhXZ0OdoMWguVKR6
N5E9xM1JSvfWFj2LCBvPe4pkH++GPfHo6Kk2Z7it4j+FF3qiKmnHd19vMfQbJya8cubNgKxgixY8
AXx/ATOv8IDLxfvASOKNCySGczjLThEXqDBiYEzc83ssvRc3fqLQuxXq5CGuGo88WcI5YyJ/66dT
baleHbM9ATsNlqS8EzS0p8liVbCJClAPSh0mF8fpXNUQKFmIfmknJ8lSJ38h4nSCj7Vykonxyvna
Yh8YNi6Y4kteAMU3rPbKbJ2g/nQzkJdwZtm0wnzmSG18AVo6sJFch7FD7KE/r4EpfPtMJhIr2hm4
cpzg/IFMkEENon2hEE9wJkR7hGu8WrbSOhXgDX3OejjV//mtvgGolvw8Ul+kMAlHvsKyTc5OOlbQ
jQMWA/g1zvs+1ybUUu0csw9UKimKRJC+D7/mJjeuQLeL/bFjNCgbwmNcqawxL+V5kci5lwxwgB/8
JYrLxX2ANXzUy8KF2dq++fOrjGPLjKOgZiic1bMNPSAlRQmFd/TJeagreWDen4V4pZ17uv121SYC
zSi1asMNk5ojVSP/Jvn08HOpol24jjVRsbowCiXjyNGJ5XJb/x0ah3zfDWllbvjdDl0g1uEb7B8V
VfzS6kaP4bF8HpMVCgdudkEpy1U8EiK14wDVFc0K6gdiQyF/1BO0TUl2phtbOH8yKyvarFehdrNf
Vk26xbaMg63iv/Zc9ZDXgNe5Bmszo0w+P189aOMD7Ddev42OG2egtidr5MVdYXzj/UcMVJUS4YNk
1ZPe9ggfvd15TE+9eCecFDTxi2UYDUOz54exlTR9QdDQIJbO/gp6DbXEhDljZkFrSoycMR0GBVza
usfwacVWxJSHh7HahPxUAxBLSW3hjEx+LOI/hOyGwThQ0WHGaIUK9L5bnxnicJTMlfy0oDFYzqbG
uuvLHGVkXdPqmG32gmh65s7YKwZgaZG5vrNvntwxoeL8Ut5wYGn+lufSEqKlZeSrqpW5iI2zZpjj
ijYYfwKe0Tpyn2xMH6tYrzSNgbyMLL/hBdSmRmiqhB8Mxq4VRkC9kFYjGZCvg6QL41M23T2gkg5m
3eWFJBcL4LNc718p/mwfYnSNBBIMhklGCiVY1rP2Jm+Zln91ZzEoNBGD8SAnxBs1G2UjWBoalpQz
JQLoUmAq4BiQKYj+iybN+SkCESbvnVvjS3BwaQodNcScZTp53yPsCuFRUYZ+3u1Hmp5XNUN/12Lk
Qqe2TX/2dmUDQcQjYOcrqi9u7mLzQesVf1BU/4gFJwzF6xaQfc4cg3R6ClzCSBXozONpu8bbexWe
Ish4Y7hvmcfeELyciZbeQo02uTBK18FWqMW1N6+z4nflbkkfXze5ulMmclwcauY2r0Jxf5sfcTn7
u++IC6VfvWrxVnEqWyS3H6ic9IrRLjGP+Ghw/fr34AfnzPrk3T6tEUbyAwTAFrKC8HKrbUpdDbsi
w1bicTPXYfBbPZOH+GeT0ek4cpNyixiLL2+9lg4TZKp95gI+BJY1j/p57g/3O+lpc7ISHmi5TDjk
pEa6IPOjN5IkFUnLI06codiXWS61nm+enfgzi7GPI595bWCTyxqDxKj/nm+N43jMhorkPGKM00T5
qn8S2JX8yfjEUwqNpWfwN0ic8FEqkoZQ6I6qsE+1ghy2YMaauvBJR0UE8iQTCRSM/T1mEqE5CCbZ
/EEVKljPbnQ2zw3DsL+NsTNtTn0U+4MLX67F4BvU0ySD29DV+xQK23F+cRoscWnxKNn6245SXeuE
o/m2Ti+w2RVW3s/9UosbOyHORc49SXzY6CZbJEjt2Qcw9E2ixQpk1G06hhErxDsoq+2s9puhp4WU
kd34RxkLpxsUH2Gb8o7UjZWBvHSqJ0msa7uNHn8B64RgGOVH4W1N0gwVrj9cABRyZVslsMOE7ZPS
dd9GDad3oPLKWl8l3vWsocc45UNYgijlW1zovJIiLlarL4QTgVO0mtHJO/TsUs6M62SK6e1WOgse
A3IMVyA8G759H/MkySQYkDFIbJ1RsBrjQnDfP4avfaqbfc+elFyVRer1OSu8zBWD3juzG8SGGT4N
S5RpW5fEDJgL+AqLiRgpH/v6TKTIbxVAMzFGR7/dep6tmkuxrwpHGHCI3jY7idoIjLnwq7Atq7/X
5OVSDbzgkR8/agFyMWaSL2LvENC4C9JTdOu5JZcF1QwAhp4Fe+tFDdTMAPhJa3+bV2rQlJfxaOUO
qTUag6VryZcHjzpGTYnD+A88+ZgD5HHFXcFjMopC846+0sDwlPc6GHmGvCIsMKzc14AbQAVv+I5f
+PkYENli8emtiHRJW0agMRnR41B+S9kTXKn3iNqTFdX2+N0hx+tCRkc9yePCiDUMwwyrCzHhT9ma
jcOBgXGaqbr/H7agEj9vczvMQFYfW0gpAOAVlJXMmQSr/pOjGn7PdurFVDWz0OfTmcGaffUNbdsn
7Oxi/VMaDp/v0jYThofODv7HU9q85rcWEGZuuqMgn+xcC5GHPRIHN2ZAKnm4/ZfMg66d8+dO9tFm
fuYT3AdeZ/4hHB+JcfrAixTcd21gCXYOyH8FaNDqt49FBKEzd+zEVAIlp2/qQsUSoM+0PrrmKCMw
Gwv87Ly5laIgx5L16qKIdeWIf5XG5WjEq14t6M/90U8VecVvetvhBVTiNp/rseALhF++Sb70dOsf
Jb2WXr7v+sftdcI2kFO8tSap1+dqy9aDVuhh8DznxzXOqJnxwVJTOWw5ZJjGecg0rbhQu2mRhhDK
C2B0waJjf+E+qh2Ky7Fe3J6P+l4GfyBWuHky9GT4yaIudawyqGU99RDrEhcWvHuRXV0QHbwua9Yw
474rgFcF7bJ/Zeuj3MqKRQfcvLeJtSpVqoLo1jxnGVP7L4KiDPzMh7klnGJzEJGTKLNxh7CngOYR
4HVFcXYX+xhzlzORQo7PUSS0JzAjzmu6HIbT0owqqZSP2LNlZdM0G/C2ey4B1hpgyoBO9n6kP5KW
8CoHjAIaRRjsFJYqWA/shXudnztjdWzGYKm04aRVxcz6zE/3L7O4lD4W4e+rKgeUaTvBpBKcFR9N
OgU3h7sjDd1CRipS3ebFWDu2vBnUfXuXUM9b8Nt4x/Ya56Ac6rTVyG1P98JSZteozR0Jw/c1FVW7
SEO7naxjJLzqWzrI8qmYBb6WYvV3xzm2uO5Cm2Yd59g3u4YRxDZ0/xS47av6RYnjqaaMt6UlfVkw
GJ3lhsOX61PnpAuC+IOK7WBpOckNiK/gCrpP67VDuWt1ZwGR9g8yHA3oF9fzC6gUz6P1ptpR8T9V
DqmWRnx1Qzl+Z38L0hCX6IGrO4j6dwkvG/JXcg1gduBEIDDQLV7sby3Og/DjXSZMtnHCaV4NbYhG
FQ/o/y+Kc/cMEmJtmhNxJFr6WI41P1jy7KJ9w/IxYTHH/eo4gGzU1N8XtztO/PW+rd6CN45zUVxs
sbBA+0t90Plx+VvLgVhFaFtXALGF1uq5fZX39A8NRHnCvQ1sBKHtH9mRwi7SNwULhGPFBfuMCs/f
9jFtedpBfMuGVoWgrNpncCfmvsT3tJarh5HoXA7r4Hh1tkxqdzsWZBwqZ0iHH1OIiaKXUsnjvnpS
4z9qAZSKQaqccHPz2TDO11uVu3tHoHvnqzfcxzEwf1UwlMidA09Qb+u2uFjCN6m+K5Ysvp6y6hbz
E3uVCc6Pm2xZkfI1GHIzNeOaylE3pYl21/txSuNVjuitl0y51mYa7Izs0bDhcwgICjWjMZzf2dVn
cmYSuOvCy8deVjS8naaVBc+F09/eu8k4Zp/rCd/2c2WSWxF45cbkL26Q4BC+b9o0pC3dw4GAbOLy
a4CWV/H/2gwJ25hMsWa2E4CD6JAH9EARZHsDsIdo84ZwIom5qWx0DwHr+2GoOGE1OwIbmDXSDDoV
OHvJyhCHvTlmPtB6UMWYvS8JTF4lZaGOCF1PX+fE/4zEIzsn30GfT5djYtm6p+31Vhl/0gAFWlL/
rcj5YMlF/tqSCu2XVx9Qqn4dwn8u2yNPfS2s//bkHiny7DEQkDhGOdU4jtS4RW5YKsnuUVi4VC4J
mbpHrEcZGN6ZkrlHUI3gkEU2TFLRpxGspcaMTQZ6jWLVG4otJy3WvVCUDb7oo7l1FUZohx4Os4Pz
aw5zSCZl/MAXklZQ2fBu2pxTUBIQg76I4ju7mdig+LcdF4vGIjwAXntugi1AECxi2cpFO9eFMP4s
m9oSURLocLilQB4ksxTNcKCt9i5KaK8KGs1qkAJCoUdKDXKUaAlHnJ+HMzJFOwdVuLxJQQIn9PpX
LwAQTTzsYn+RY+CefUPAlzHx01seZbOZ03OxCezD/x0h5WiHKDpKp+jrjM3y9sf9e6uc1CQFne01
heNRxx+qTTzqH7ZQW9AO6O0HgcQSl8etuA+SUeS6Bjyh/GBoVwpDoG+Fzh75qBTIihmP55PECZQS
9KoPr4cqa/+roVp1IZvxJkQJx6Jb6fuGTYWYopIT/sCb8AhNKa3w2k1iMInwYxHk+CwJst1QIiTs
zsec7cT0YTvaBBPIH6lRYaGTblced6OvUgm/95lDIJrz//WHfnfQrkuoI5YDk2w3bBrlq0l2nF7d
AfPtYjGO5kqmZfKsPIAz10rdzfT2gtgZOjZPq33IA4XbEHkbyoWKn5HQbBf1i07xPcfhIi4iniVf
r/i0nD6MmkdAL805HkdY3Ffq9kYVS8kn47A7Fff42IovHe4KD1z3y/WLYC+RxNt5c68EqsZgOa3M
BsjjPpsr+vrrbh7GhW7/5Bamb51vWbAsBvpaYa84XZ1d6IA0LuFl5XsZOXy6AuPUo+nBxtSO546T
kHygw3Nzn4fS+D6yiIkbxHcKnMnDAqD6CeyPN2OFzgYtum2mkHhIIvKptkdBmAS1+EhHY3qcX4XF
vFAywdnsgmqoUrz/hZ86BcTgmVRfSsGmndoymlmON/zz64PxUWPL5NNmnMdvWTk+5u2sEPKEZbW8
CYFEs5ZVqGFykXlvpsq1FmrSVq8creiZWNHj5mdrGyZwNPD/Y+pUkf5D8Fm5KUZ24hX/kpmnNUSo
GR4b3JHTmApeOSeYZxTIxPGXzI8ELnFFuGnbLSqBm28aMDolD+jZC8KxCMW30SuSJBp0BS1dPGjL
qEvZdFlrSPzF2Q9Lp5PnalRMGiruoPAl7n0cH1bQgrv1tt/JWffZEYXrBiXfDiwjs4yjHoPC1+MY
pcQUPxhuZC+Y1iIwkWIbVHIOu2sSmnPnZdODXDyE9SFGYn4P1I73EXth5ISCYhgfCDEASebCsRhX
RypYJcPmeX9WJja1pIiR/WEqkMnT1PDMW0Gyh5S5Wl41LGgJLg32Kza554pMfzPf2vOK1Btv1scn
CbjUccu8IedPQTtoIplnzSPY2pr7bjw8GKPF3wK6T/RX8EPLflnHDmdYT1MnOUBHwbGmMAD9bPKt
4D+TX8tJuiKPdBKBmqb2nILzrLNRHr4jwETVyREHluBFzLSyEcTsBeRwKT8SFA759enPg27THQue
alC35TnFp0oJgZ5GZvECt042Vn7xObCPvgMfcxY77+UjLLLuWdzb3Slu8cd8NrrGh6kYXr8y9noQ
uqXzf0etVQ1G6sWGdl0K6nI5B6rUhZGTTZc3YWv1gcnPngbEpE1vJj4W6ZozG4ZQr4T+ygBhHeS0
W+ImCYqSYYkdyWNl5r+tn+yMniVAfc6/q+ZgMi+vx2NE3f3mf17uxXSSh1srTvut/njs2DOH1c2U
A5RcroW/82gneN2n3ZX7osw4Qoe86QLkmte9AHbiRzG6ee5VzP04sW0blZa0clOwJHHWR95GpOG7
QzfLmBJbRhIbcpDTM5PRnnAH/BKW4lOLaWU7SOkfSjfq3EDV/c6a5oVPEtZUXVJZhJafMETmZ3G3
UimpIm2dLF0ph4qTrF3j5rQB61B+oio3F83aj75UqpifB33Bl2+IGRemDbpQjz3T6uGe7KqMck/F
DhNbmaSkcmqOiaYRthRKnlhsMJXlYmFAxoasFwx9tYmkBHAlIx5VHzUDjdv3tpHKMaDOyK+49IbA
jt6+uYSSvjMk1ISNe6Y80Q3Uf7LVBspMgvOQcTBSivevt8NodahhUW4d9oTRdV3YrwAbH2CAo28j
G1vkPbE9UM/VdE/NjI53wTzZc9tPhOj8FmfGE9D/hze9OiqOqjC23bkUhDJArUPR3VyYnEWNH8N2
sc2M57+i3/6b1HtowQ7otubjSTj46sG0oY2clXSiW8OzgPk+DjMOpPS5il8plqYap3BcWS/5oswm
7DGSxeHzjqylQtQR2MH8h+UMHjqNgXj7ubUR0fXgkBqNNGfXoPEsMzoUkKS4rYmDL+SvA8SpTSGo
YsY/ys7IQWDkTN3P/XYH8xwWxmupF9GuuC1xl8bNkneqMR/mdC5YRWTggS0NH5m5F8GrzYatyPV0
dlqsP0uCWqdyGNsNPX5oBEa9qI7stYA7YsSNwF8C+VKfRQ1Ijk7RyhUwqDpFY9VJVtQSeu00KREk
FxPAaE4nLIZRmFaormST4FyqxlEgu/jdxS25JrZ/8td1pKNbqKL/oqDXCH50xjWE8o21fV9Nc2uf
XCdmzD//6q0oJdi1q1UIZwXymfRcy2uKbTr4ROZNwDohHHorA2ZJ2qbQUTpjrQ6ubsP4KJSe60cV
KKCsGT9gfOUfSj/+lkDVi5Ou7lkIaR6IQGAsFMG40+1YOFmuDLmji2sWikOWEgUeKYkAumz9I6qG
wTKEVst5pjjj8tHTgNYMIbIRdzZkTXy7X96yOo5qDKiaF0gL7mU/AZPlq93vuWDghu/HQXFJUH/p
EgIIbUaEx+9XCxOsc9bs5+nB/paHK58H5XzgCd8ByiuRayZ166Ad59XgZuIcaU4NRmWgPCpoSR37
zlzlaH0vHeXbngcDoRySKwHwo+U4ApovDqI48pchq1hXcyemkvEAma0Ckdhk9SZx6qhyW06TIlos
r3oo4Wbm3dn2gQLpesEON/0HFJJW7eytDuBLao9F8yqyFGhk00W328dDMXYvG/zaEI/Sl13CwcBB
YVgjEPsnQ9We+3Hz7sZfLcQyI9btZXVidzZ6oLnCtCgyyWjWUj5l2TmN+13/q39GrK14A/+xt2Pb
KiADKJqk8m7CqmK95SeBOWepYKVFZ1s+69mHAaOfuav4RHlJ/HpPTojD7KKxg6Zc5zwXywDfnJd6
V/k89MaHjkaaIMEsDWQx+cy4NTdylBXEdHm8/mJyR3TbBeQKN9GwxtbOFVspBSWs4aA0jWrP+173
+wmoVijMlYwyIHRl92siBikUU0XYcN8lHCb4LrIJO2tYymh0pDdEVEILLCK84TB+E362SGy68z1s
zrrACiZ9841l5p9iMFZidSPxlZuNTlWAoJK/HjoFJGgt2mU8/RVpqDsi9/WwmAJJm9aChsncHOho
OVk2xShS9RIBR+tDt1Xai4kNO3O1TbckgkvoSCYLpFkbv2bF9S9jU4cypS5QL7bdYbd2Pwkt8y9T
dB0bsB+lXyxqpko5q18CwIDdRhZ5IftcGdcdPQO70PSfRogvuLIT1yn7IbmaS0MzziLX3tM9ZsQ3
wcpZiQA/q29sXRdbzqV9G49VyJWMSE4XRR18VW1QIPfmmPPOTaeplkrr97FBtrvSGKefyO4tn+7b
4AKgvSo/iZjwkmtz05RKxH+209Oc9Dv5TDAUJHNdN5K7OUAe7Zy1VPFbNYOQyIozMgUiyTyZLxAb
oQV83P1hx6KMbk0k2GQG6NfGALPL/H2LwbPgZPiThBFHcB6I0SCCJ4dYXj4PUS6eYcvU3/1GKp5L
mzUg7RpH/uq+2zPJl+PtKIXq7VMZpDPWTV/7uFsNJMZ3R1UorDH24C80b7sTlUJPgNyvi59eI1iI
Mq2dN9rYtCGhM6pWdBZGNYE5HYAQSv/YKLvyFklBPDPUotxdDIZc1hbWMOI8JaCOf7hBmt3DB8sJ
thxxsyBS5MQp+w/+xjIE4DyxoSfcGmS04yNe7+mWd5Dh1mP9BRQeKaz1rmdA6G+yXSVYT+MEMPXP
ak+idJw5OrqTrgWBILKxpZsIlWTfKTbtN5b7UBL2LFCZk0aOUQryf6wBHFZA8b/Wcu42lddp1Rel
czA4jiaSxYrD72LcnpJccOewf7WikWctiydP8Nhdo37ANTr0iEcSEq8uR5ChL77YCEjdhdsyyBLX
5RXOtN5sN5cK/fssPtoXPJMZYAOfT3sFtaxa820lAfy9PY221BS1TWtpuNd6qm9ady4LwimMeEYz
0NctXDUPQxwWuj5NcTU8m1XbyT5gpmBgMKOCo/abe2SxQDAF2trJdZ7g7bdRpW4WjExFmkdaGVs6
w1lNxKzEk6oGKEUencWmr0IouYNcxQnOA2NG+p7xuzyYya0XUaa8n9G3j9VyENCdAAyJsx5+SLYu
neThWVtPaLfHbLnSWl3C9dXBMOQgB8Gy3bUtnoaGdGsw/d4OAQXrClX82PfOmDSxM08n3r8HluQ7
V/xzvhLwD9matZxXQSxFlkqd2kvPCgd3dtL1nUM2DO6u1bNdzZ8GZKMJEc0lUDf/1oXuxdb6oGH4
05+AznsFRbgdeZzBS0lwRXioem1u2mNvuR7PS3vQEQ4iHcTf/ZPLGEjpwwngnmAJK5cxLvsmI2nI
VbYhC5zP6JNfAdEfQnpQrZMy7HPdlit8IW+XxTRBJyo70hl7DsmdOE6ATe+dDMNv0qzQngIIPhvt
m2Glpvg0/9edxVq9n2YapTf4OS/5QVg9Hj2aE6NTKi/V5IFibd1OpMYM0d7EzmgmFh3BwmoI9bUS
KGcWADWMrRjOf3n6OMl3gUKwuucCU6RB+HWHphgFomwU6IGcztkZ6gn08JQofzVxtkuqOzJsabiK
F+yebF0AZynTZpwFhPM5gAPAYE55JgFv6/4odAzHQiufSO9bP9MKcxSADaQWDRnDeZWxqt75uX8R
2UHcUbYV41IYPnz1orNVVs/HQNeD+rFvISwmuqAWG8Aidtw0ll1fmC0i5KQZ4v4UIqdrjn+pHKdg
tKEIMnVYbUolLencFegi3Qpa8csWbQEpWBoZHjEShU1rcHuOw8yFbJzoDilLd7DqCRQV0t0cEHSy
rAtQltE5PrcTG2nexaXs5FKlS88U1DAo/+Yuf0wNDGXJfjmMNu545rHGbTEw8KrsFHoHxIvHLy+A
erCE+F3zs3cOR1DO/DRkpXPqelaTE6TokRfUXLUrT0tosYSeqAaS9+DkzFjSl0OmhHuiv+Osy+Ij
SCYfLRFFOW++KXsFG22E5IrvmVAv8d+jojYkHXUke9JuQEzTqliz41rsn9uLoZsbpdpC/TzK2YBN
S8OoT/AGNfBvSeaDTbTw084Kfeg/NMXcvFh5aQkWFThNqpBIxKrxllg3Xizs5+0wGIX1gjLrphOB
ZveSZTrpJGM9j+EsVIrY48j2bJH/jN0GG+5xDT+6Tf/SOcjCDi20NCe0c1zINoWLK+abVJFvJaA9
EITA7SR9Lj7zi916zprnfQuXFKji3dBq4+HW5rG9Dk85vEPsuzNiGXQgdsNLmMRDBjK7bjnfZXgf
WLN5wD4lWDjE5IqZI/oNeIa7Kd1plELg1iLtZcXP4iXPeI9PAl+Jd6UadpF72ijRMSU6QkxTj+2a
2vblVtKJXYjgWZsL3WYTzTRr+9fsYb0HUBE7LHAv0h1+sqxcYy+er2qX5mNAOTKe2hPgtI1MS/0t
LtEhvEQnFnGWwbPHimD7kw+1TWMsjlcWkBfUMpf7NO1p5bOX6CGfP07Smt0NynbMpj74xDBXMnO/
fMO7DoVoAqCoSuPd3aUXsrjedANckneEKPxcoySyXvRMQsKOLHlmzmYzI83iP7GBN5Ygv7ZWBPa1
bbhgOUxT2hgIoBnTNZW/i/aR53HZ05RVm1kGtwD6bTNlpnCZAKEwV9sRvsZXgxW0KIXsftY4E/QO
jLZnVNgOyZLx8Euzgmmcp17m7MmzoROKlQhtmz8jDFHrDXC38Gzk/UNsqQWc1rlL+jD84LwmQ40h
/JHnGtv2XiO0LeDNb/nrhTCq/DsE0ehlcNWKCp74o01T8EZzgwPbSVhDRHz+45FxUnF/Ctbh+obe
mqaNN3Diwi69sAR/CUBUIr3uXy3p4nKkwu9EU7z5Yg2ia7POahqq7bcd/tkXbtVSFxD5IwzgP8r4
kesDtTDgixdBpX+6bfGfXdo3SV9BlEYcAGHWJ4/qhkcU4e7WUUaZxPxNqYA407lZGBVd32lfSu6Q
QTLMlLGDOiBOHGkrMUFra3/nYvfW9oIAsFXg5unpvuVhhEuOWq0+JuUc6A4zPYPWTrZTCgaWLYmy
YEF3DRu8OVe2IUxkRqSxBm4zctmmUhXcroQtGsYWpxASRrRIGr15F9Z4U672BYywVFWUWeOupVb+
MMR73svUmQiGqtHxHZU6hpwfmo0jRnCRTOmhw09IImIqFe7CfohbOjN2NTR7l5A4NZeNGU4cZoUX
tuVkMV95ZGzJ0afCRP4p+bsBBhezk1Lhr14+2s8ioe8CdtdP2x+CrOE+wGNb6D4JN7qIxNkNcPkg
GUTICPr+LrEI2nsMXFdfmVc5nqPJVgFN1/+V4QLmz2wgG5DXqtYRJXNXPXROtgG5Jo2Ggf1s70Vu
Toci2n6TWU3UHyWgXl7dShHwlylkzDs5r76BIcUGI0qKOTk/zVDfPCGknuwzSPb4jt0k/Yhzfrp4
tyizKyr4Vh2rZeYkyqOqww1fH9zeSMTkeTISiVrEbu+Qpv2Rd7aBmD+yH8p08/AzosNi1+lQ1+Wt
UyMWXRWvWdVb27IwuXAcxExtj8yRxEVhLlek5bhCP6O74Wqbw2UjvZ/QJHtKyPN6zCtEaDXGLQP9
b1LymAaTW9Db9VFjcMk+sqBO3n/KI1iOmbhDVroEKkK8JFp2eGfqGkAWNYvtEPepbdY8qYMw+Mqx
W4yT5kj1YBkgqTENNIbdJ0MUcPcqtJvkiB2OK3JlQC4sQW20a0+qZrRH/CbvkhnwNcGgNbgREHlv
F/3AWXGXTK1T1qonqpCkuMYcDPTLvWSZAB4z6ESUzkvu4oMzdl/R6at6ZaI9yVVrbJOHZp1GycOW
TIePysoS/vX9/y7Gbwh0qhTE+31/xwxaAi3+fbd8fSG8E3w+bNRAT/9ux29g5u9D3CWDuAaBpg9L
G/W1HQLOOvF8mf7YgFE1jEsg8xQkKWoPF6xuDOeQM7S7Hj4zb2rBzzrzy4tNIv8C7ui/lbsbkiaz
YqdLo2BZc27N6dAnSigTOA1bn44Das2+sGjqnDagEAkIjE0U2McRAJ/fw/ZU+7Vn3DyR49K/B1EH
Sdc2YbDYIpDbHsHrm90CEX8SdeSA8EZ6ZvduA4SFen/opPlegbtb10AbJhhV54cLjhpAB5Bxde72
urXWCWijeggEQIivukswWWZOl5yWgAv0kjYByaw+omVEOso0s1/E6vxbvUsESTmDqaKAG+8sbHl+
DC34CwK7O9pdjuzVFJrRYmK1qv2+oUsvF6WRUdDWiB22V/CwaN0S2mCHe6EcSfKd8ywB4msgum1S
dpkGdeLC4lDFAf/gX+LWvesaJM7FTYzeYjAJUgcmFP0DEW/hVTWhFh3sWwHl0CodO1l81RmTYoDC
vrYWGsO8edh4ooXwpSXP/4qVfIN7Np36uvz7PoBgcqulsHQ6BdeWqky9eI2I4Li/8qkgDi/44kQA
XE924CgxrVqArBEE9Ck2lBpBcimw0NJwil0wwueTswmezEs0O+MwADfTfOysMsKFRjQ87pb0Xtq4
dkouCLwz1+hmL4DmlNwAB84CWX+/tblO6z20mLp9nBSxpT7TOVwJM+dHCEJYkCulWiq9ph6bY1Kt
jJAEHkChhie9TqXWU2uMp7e2657FylHKlML277mydInxHbdGxU9D3IGWcGW9IaJq8L+IMxhITxL8
Co4I1sdiCT66ciMoYCL6dFpjy24Kd2TmoaWDjENTTct5D7tL9Km2jZSEHRTESbIrPiNMovzw8Y46
m1awEY6hIGc+YmsF4WegYm1iLgUpMKmLGRABV/n8QrhyzZX+SHAR+VMGp2zZQB7LqNKg/6/xyBU5
rtwWwAdxX+mfpH5lvl71aal5gNAfkPf2V3qR7XTFhcK6bYWbD9S8X6hptSpPYoqAmCl33Ghas4+v
z2VQvsMLUo0PYJGTwAM03f8Y1HR4rZQwDqCBafqrf8Hr7Ap59GRC91D/qGVrShm7QydS7l4YIds6
Vk7Ad2dLJO4X8AWHlXhL3ffPDvR0n7Ot1ezHNTn2Ue0zBvxF/vXqowqgHD9m24IGmgPRh2byTmOc
O3KyRpR92WXMs/Ds+yCaDLu/P84mESfnIUHt3qKNzX5fmWrukqg3xbit58rhcrbY+yvA2GI7sZZh
kVgYVgAIme9/G5sjfkM+PpbzgzpXfOsiBDgrX7FHq7WGkC/R2BgBybDDqMz90sTK7WOt0YD3ZVpM
ExdXKbPEYBoKUB2LYN0eM+AnDENmu0Lk2MEUs5QldaOj/T52fKn52NWPJGOBybYSES3nqgG+RKks
iR+6qH6Gd2+rf0hPAl2DO3M4kPbtxOLd6I+kVawUrp4szEQfuBcQix9nILOhrhY3aq6FB5iPN6Dk
WtZhmhuvDqDD/6bBpEO9VnaWybGCbu62hmt8Xdsq/gka9m46XeuhMHyPeqbHo5f7ibpT3PRitO6e
WiodZtEf7oVK7+s1F00MxAaQEEcw/pY2WO/Q95I9mbrpHas1HxaI+1vXqbTdKiX2J9tYL1pbcnzp
ltYxxIEQPzfU3DjXv4VHz/ymMsKXO4BiwmkN4aAvvv5RudtVxRJNAJdYmb4a4gruuVdbV8LLPQNB
YNuCoWxXgGOUM/jnEdGxWERibGEDe+dH6TK4lL6eq/Hz6NI4c1jFAxDGsI2zZtUZNcTc/2iaxyUP
hnxgnKs5OWNZli/DAVARsnIB4n7UvDfOaGZ/fC92zexCfI/ioswYgvc/yS1TiGtBTHSzqc0SlYMX
TwdIlvn1QAaMqsvD05BgnPzHEcmPeFNyzQwpBFHpkxGOlDcv5rnlLIdn9VtrkORjTPZ1fKIysGqH
UQw7JXtnXMbwf3BFyuQ7r02AqznsKZ/qIwGpDQ3YM7LYh2wVtaFPbjm6+Rfs1kx2kAGqYj8TNSLo
mXk78gnOK1zPXll9OZ7BiP+cvSXaUeUyJBL5iFVP9BRpy1jJDYAyn7vot7RsbusZj1P1/6oDcyl8
RBZC0eOI9msCw7xIQgvJ+rdx04WulJdo1KKvqnQcP6D0O/byZmOk/wpV2kkHjtJ4+uWNkJKBcMHs
t8tmQ+LLtZJoH3PvvpuS4yM27DjIBd6qq8csleeyAxKO/ACg3V/yn/WVcp3AIVZIx8qzUtD2E9vJ
0yX2+FZeE8RIGU2Oxb/M+qq6TbUNC2X2K61t4A3LufDDBViMnvu/NJ9nq/xcmwFgIC9sIkYpoQmg
8mRwzdP/yeIcJVudil5nP4ETtRu/pa2MJokLIVBlou3/UdWTF2Ep976hmgPlOMkOUk4fItS37Z3E
jIMuVGCPmetGUlkaDYYNjolp+iEuoA9mDclt8qjuPqOaN5h6yM8W4iJLjxVR9dZaaYSdqRFPODY3
VNjLsk2g/ANWuUhIlGLGiqg+YrvbeYhYJWJ7Q+NWHopTR2pFygk6uwlGFGTYoQt1BhtgzMeRaiPE
0L9g/uf/7ktSPxs7AwkonygtRfRRAA6fb1CKnD8LYtDlfTiRF5GZHB5trXRRT8TuNwkNk2bQBZsa
u2HiYsHUcxeJ4YZlEQMynP710CmHx7rm3QJ/ogmbVPRM5lLLCvxcJA9gvDeLJMHfCh+FH9JWT3IS
RfJkdMDBSX7e7MpLLcyWLH/KpFJ54yYPlHfhROwl2+LC4tAASCsTv7OY5xhweA+sXRf1dW6xzKHv
tEpIQZe/W/2Ogpij+bTUeb03mNNoU+Lv1+XWLepXyuChdNhOwJHmHYWZK5D6QdxanTNwSmtBGrVE
T78v+UtCiGVJUtw9EJJmPCZpEkAulyOUJAAbEBhann7Xn8faxApCFenK382tWYImezvWUp7GPN56
cEaR675DYWVA6yZ5Mev28+340Dm8+GuzWACllZug5bIXVr+flv98Vintswzi7oeRPPhT9nWeHpl1
s8/nZ2Czqm8GZN06TqYgS6A/Aq9X2DlSwK4ce+vKzIuogFG4lBm7IK7fj0MjRTLUi74YR/Mn2ZgV
W3Rs1Kko5txn345BVmBoYaKXZtj2eRGKgxsPfNg5J7z0DBjUTV6gjsG1W6GehQO7F/Xkdi9h3mD5
JNSyPDf3ZxCGphrcuaxWii1zqc7+lk/e84Eh1VGhLVCfwtmqvUgCKI5GV0YcNIBwdmF5uMpSQzaG
qSeI6AOPPLYMTJTAVVOoMpmO3Jc9WEdkkmJk8J7Ps+yzVaW6nnwweq1xsIWoomj+QjkPWpt3RWil
tuZLTuKDrcq38uXUpoo8+NH07OTdwhWo9OKoGpEHTDVcJthXhcjodWXJKkpRmJ95CSkmwgKRzjl0
RMPZE2Ho98MgqK/MHrc9uiFYiAxuZKwlQN2+EEf5nEZwMn9rHLqqxH66cxbXxwLKPaNb6PhqcKX/
ZGjZknkuM50jbZFVJtLAmNg5SZUCk67Y9LpT5SfqYG0+MH7/I/Ub50H3NFaqCkeYmi5D2BsWn7qn
o3ArzAYCdpeblO1uqN2CxGPUuqZ5+pZgWXVxaiI3rmt3XjbZr3lEXNICn7Hl2ee4JTUh8rL4zi61
dOzaW6Rzm2mciXozihN5ZSo80tgjfRmZsvWHrVDG5OzCiuDkNejJ5A7OjE939pG8QOlpKRqHoqya
EvJ91iJiNnjb45Mv7pcvgVfUEtAGLgr82iDmVD9BptPqoZkmW+OVUxmNKxhW8RkB+0RABN/E6EkW
ngmzJdFRon/2DP+a0uR/IpTE+Nn6gwBfeIm+fQBAG1zjJ2KHRri4XWzqeHdHNV/x0Rj7Ekt6gFkH
lY3MyP7n8l6uD/e9A0WzU0v72fwog6vnmk7v+Jn+UaR+CnZO0Sg7FEvKKFsehysXoJHNaqCByiRk
hv8nIjo3VDwv+0f1vLJvwLMxUSOcgvnQvroBIHq+OHU+6vqQjwqYIDH9MR/3PVGFA/3MknC2gxQg
9faenTnnW8CE5O9x3VaxZCqhMMHqxp2XNh04FTyOEzM0EOFavLrf7NLIL73migzB+mvqJMKcOJ+r
udrb/fBUk1fQh0k+QlB62sK6vEB5wY5DFmxWfovPD03yDPUj2/OKUFKBW6M2QY0Iu5blzQMgLa5X
o8DUNuPyiG+yjCtZX8RS8tiWa7FFQRA93NYYMzOYuzj116GZy1OZm3qCJqFjduO+pQEiLAvJ6MiQ
zDprFakRcC1Z9o1Ba6UY1WbIttD0sOJ7Q1qdFoDKylzecFB2w21Fg0Ay9/FCwz3aDx2lG6o4xcLC
ZYg4oWLQ/+0lYJMlxEi9dGLb/BZ3iPVdDL8peaJymbwXB6cSW3egzI3hBrW1GvqFXE6BEtgAJurJ
df0XdhnpjYmvTyVvR3bivWl6bJrwrA88vaeR0xnfQAj8hmLqgBGhv/IfjxM6D0TPKvgzTSst9FOc
c2O5PSCsBDqWlNsYUvR+UqrXStgCGFcomxrTjydjUnYFo3hBT6Zro/kQjaS4vpCJAxo3HhirMG+Y
GQv/vNvZbN0Bt88RyJUOzFJ/Xw8F3CBaTR74MHENECyeIvd7yzTMU4Ruq4xZFHX+qJcCDbrWgkrG
rSqE6GoFmmGjaGDGyhiINefjAOJ9iJdkPbyMSMuwKnLGNv4oNadkoNQ8FdM9eInCNPjPVssYbyhh
L7rGoX2NAvqM8paWfo01IFFmjP9cD5nkFdVxkF/RV+HuEQYOhWpNhJLKk9aGGEJqeBxUq8vyte27
bY24Tw+7LlEbBQN7SkKJw9+U2YS56T4fCvvMakXA/t1vA1xjk8hcCuUXPG1c5OtjosRA6G5ppERL
cZwHjvuAxdvYOd3gJutzuxwCGMfoSVpynVNV7pzOoIyqCmbijOmYtIQ4upfRJ5XfsvUZHGDUlo3u
OIoOYNLmihhE7eREx4GFiU68c/BHj2bNv0wqKbw+BYnhAQyqTt8vjvo/xaQO/yvUIFiIAvJBMYSA
5gtg1z/5W81gFw0jdw7iKSlJ61OgmbGoQ0CQcPT23NOs0Ak6A0qc3suWQI/SV6KwWbRzcCGEsn43
yVZfukVjmLICUzV0Qx3057I3XAcWCxqehSfQQFutVQS20AA6uGoACdhn4UX6twteLcsnLTAg3hfQ
mIvg9qrbgOgUcyE4b8LLFgeoXkOu2cowUpsJxmhtKERUpuRgV5IBbrlus3ZKmREkS4OEPXS2K66H
txpK9vLGvjpUXEpTPpifFEZEVngJvSVnAlfFDf5SKDgks3nbGXumhxs2qL0kUULz6CnLcBOxi1sc
xbdlbsrxuaHsU/lIwnXUV42jL3WqCo0yC3ew3LeYv/wXwTfVWtPqH7sbF4wjpeFJBrE51JGca9cO
rszkaiUAHk8fYcljhbjePHBMfucfZ5G40k6U4pZ3C3jf8lFF3+B9SiNOTL3oNF56GYqiV8HkYtb7
qDCX3x9tyD+39PyQCNg53lqrlOR/DQeunwtkthOfQEXtORnC9G7uxrmGCOYF3LAEsFXjU8Boyp4U
6usHfHI9I07d+YRxh09r3KOx1cBWpS1J5uz9a0beR2Q7aYhAd1wZcWQDeySpzywFUT96L3/hye6g
GXUD14K5DW7a0OchXbPowIPm2AF/Jg+fHAX5bN/tWEb4JAIXHRHoPKHulnZG2/lHtKtU5tjuz9g9
H2PLck2dVRsCBSNwt+kUh2KUvwhli6+W5RjxnPX1RRkBQBoaWAFjAKLyCUj4/IsHodPGQ166y4aP
2+PBNpmYgx5lvolIeR+qJnlScYHsWpYQAD+FOXaCFI10LDJ2hKnrulHqD5By6LftIZElpGCeD8Lh
o7gKMFh48RTNqjChMFma9colTwXawcBpbuaL8ho0ekU6CNRsxey/v8g9ewVEi8kC1AXi4mHV8qO9
VE44vFV4cpNXyIZUPxpA0QSRWCf6ABE1K+e8MxAcqztECVhYAXuxtxxoqiKBUFpBTOEY6FW7/jqp
nO7bwoVzhqem6ls5DFiPBxiOiOjdlSTWe5nQm+qA/SQZlvBaVjHZnvxKzid9ohYn8vZJ7vJNegjy
rLLoCyQd2wiTpud1F+BZDR4fBR5Oe8PaRulMkriTp8KM+iT/FIc2TvoZ1zoJYOsG3xm7jyEIhdQ+
/foL+E+2dMdhnDOptpFJPAcOtf7+FmsxFvZKeEJ5NpWHq+yZCcVXbKfhQBLV9pONu/cWmm3TrbOE
CGQZGDr+TIxfrvdw8PXu3XaMiO3aUMBqDMAsH0nwUA59+aRKS9FLKcl1XcmW+3HF9Z5UXnHrnlWk
IIQxlSX2Evt1xlbJLz30LX7jmkoDdPkZVBHxFZkDe/nk2xJLxq/mMMP1jQ5DZX70N3Zd3fge16b3
83iYSaQw8hZCGot3DH4+eyZZeYoeH1A9bpWh6Ntyu7jQhj+U7n9qIGL78PnmtZbgTrfckv1tWaDP
iVh8sthuapkHcep7MeXxJtKewWQ7B/VMAFWA2YJXfJXN+S+yw7dK2kyofHT+DhrCtesNWrCGgfeb
acAEbIWGMjMFktpntrmKRtWO6AsYHc4eeiLWElW4B566IsdM4Pa+o8Wd3MOe5+AImxJR72vPNDvx
uWLAdpUECO1xquU3KswQ2qZyBxT50PmGMynKsuh3uiowQHEro9nRRKsVCmmy8v/fyO5SXvJfcwf7
rrWyn5c6AlaUrB6C8fVAyph6VDdhskEaBj2KXM7/uG8xdQh6HA1xy6bSmBqxsZ0eYeTzByV7tcYi
/0q+fSqWMZtGL/WbYuGC+6vESveYAbBjSte3SntzILg/KwWigRbBzualCnQrg9fiAoJxzo5vLGny
NtulBwth+SXsm3dUGCkFF3K6oGMtz11Q6d736OW1t4mcJh2CQ2sCAP1QNr5yF3Th9DD9navdRl1K
zx4rEseQLSdrIp8K/AGGz//qIFToIcoai2T8NaX17mrmmPVg0oOyA1JD74O1/iPnldHnPlWZa78N
F8CJGeQfQnnmgORWIpI3r13fHOcemhBFebktQcPOBds5jnrwLEaSUZ7PRx5s0ZNfCMdTt7Z1oJTh
lUabuLGAd50H4cVVxbcbCWt9COXFtaOkgGuT9+8VosULueYe5hjKy6rmoxdigEKIc3B+IC1VI1nN
GV4Jirpp/QpV31bCwv4dwBmbYg5KHFWYLuApJdAa41JS9OEufzvhD4wWu4nhue+WekZ4YZOU+LEE
zO233VSXoReiB642uHq19ufywCsyLajhnRg1MQ+PkXr6X9LOZvy4iisZAADmAmbl9NX6wnXwDS6J
THMl4SwETYYV8LNXkatf2CRTcR4T/mwwt+ITYHRY5kAGzXez4ctpYpAYTOVnUKtGb/K4PsiQ7Is5
eoj9fAs6i8f/jfLxXhCBRAylQvDNhNOIa85oOrmVsL5BhTJWOmGvwRqPYyYOm4nSFjt2YubSVXwC
v0AwodKvPP5gkjyOLYD/OPL/yzar3pBlGCwD2uj217kx8id1QKwbvAxBu35SxyzUX2ckHyCf+Rst
P39doSGUfMV+mm5rV385vu5ZV67uXct3BHELGTTDolGYl1KseW3kgTIGOz/UxnbPcpgelOiWcp9X
cwD2hg6GZcKmB4kdQz3W6fASXhXRHh7tb4uTF7iWm2cYIKva8BUIfgJbfSIOcML2FNKLSsnui9Eb
SKrPNYFItzUMLHtp7WxD3ezBF5bTpTN80YEjXd0p8vXjNiT8WpmkS+ekrW0mvU+CL0g+ug1DCnU7
saILnDylWgpZw/9nmydknEFlHB70DwmeEfI5NHZba7imh6zqFwLWiSuG/3y3z96MsQHi8OZ7DpH7
JF9gFUbciySPb2kQ8fdEEvmPpssuziOMLd/FYkqe9Q7coBHM6QXFlmIexLhkWU3BneRpvxpSmuZF
a2rLDpjTggW3JxxgQQyFxJNCDBxpDgm/IbgK7LCWu5kdWOHwsQL0ay/ZRVuQk5qbrPj7TDitKcN9
ZHmzDhX/MxmnF8doTk+ID40bSmy46ZTyFIxSPX4UbjWbyN1eRhHxWU9g6dlShHcxHg/2rcoFs6y0
mcWL058BY8YY2Vhm0QoRxRB5Hv+bt/6SsBEyv6IxFAn2epO0doEzXYiP2n8dy2V5W8i5ACbN+sJp
nWRAvXIcUiXtdmnr3oIppBHDIxq41GuGMMBlZAKYK/SHOOOrwU4HZHE2Igaj4KoFineDUjwxn9TC
eogCc8B4j3i7LSvl6aBJGmyTnJ+jrygfUOkzbbBFi49FQ6tynAqcLV47GofmXKcQAwLnUJz1GpkV
L+E26SyY45oMBM7IJnxuyNuUYczTV7AnfGPA7/71pDcnnY0kqbzBseECUf/TclBE3uXeEUtDYu8x
aUcR4Riad/muEgWTJKabQVn+1xh+PTOpQt1Jnq3IJiCINUL95oJ7Pq7CUMyCUza7JcwSEFVBKgUl
vtZgdxQfUCFjwvrN4EAqdhhlkVHwG+nX3WBtNGJum1UnKFretDoK1t4NHtNOrZpqMh5KTwvZU2uS
hl1QVhPiSMcwtotAzHJP1bcznu4Pi2qh/G5Q3nI6bOed3Q0nGFQL6pHmxgl3sjBMtXL4zY5Kndwm
x5q6saWR9xBF32TqYFr2jq3DUQO4shXQFmC36Zo4mHHHRcmrkF/A6nng0s6pmAj7hkYUJvK4Mmam
l/xo0t1IFeiED8DUNxAWSHuwOvfNMIsTgrhoRFHsrdd+f7qoZJQT/0lJHW8qE6bNu3d7iX9XA+Rg
hrAnuq92+ay5r05B5CFs25lFp06eihQjzMVv0ntVJh9Dr7bUrQ8OgyIT9M/EldgN3I4OmZIQ2b54
M8UnNCfNMwh3g+/NaNj4wSjBmwOlz9qTYgV2rW7IF0S/QR5O2jD3nr4JzPRsWHUyZirZyn7uLY0F
qYgCIFOgwizn6XQCH6lvJVnelgWxKcd80kvtaanniTfLIn7upGx40VkSgjcHoOeJnKaprJEpsGPa
EWN35sTzkR2eIG370dBonDU5LKeMH/iO2Aq7ZW89z2gRfqzZTpamaFFHLlqZTCjZg3jGmXo1EVNV
zVxMQA90LFpr9K7aeAB/KgLQPR8UzyLHgPNWlb6xp6pUME+karsJ79AIH6CNJYY4nQSXdP5Ehe6J
jtxKhHzmlcobTAenwa6yuYdvowhpsWxmDDrKznXnN6l1OOCJ097GkOrvdAjiK7EHL/CB2m8NArA0
gY+Nbc0qMd8TNbhkgr2r3MG97Odmp1S+O8PG8K4fjZzJ1wbbhAeCZO2rShy64gALHGEdTkb1+q7l
P8rGSys8/+jctf4vbTeAGsvvYWe5DGgZ8jmyHNoFVfRVM0E3XZDCWLRJhOKf7GLojSE25nLs8Pv3
2atlxgtsH8OZpMKXDbFESMf/PwqNTsQtSfjpOp7UwwlTfy+BIWOUwY9dXZlME0RvXVIeiDGQfvgh
peJ5coJpm4BAqrxcyJBaq6YxZ932mHmEtXR4NAhE94qOhLnqTrM8S1Ny3XT4/z4or24eCYdsWv9F
M3DZdbvROE0jKfJQNtLCVD7X2mCiulsYSXXm1w+H9nRmgxS3WQrWR3nOsUiSEYap0KKrPfIwRK9H
hFj/EPkXjMLibj9vrL/VeV1GexLczgiS+MWQEavhTkinKCrUud1qoSIpA+JVd0aeIOb5P5q9BoiY
innOzLLjY0E4T9k/v8pDRNyQGPYCmQHlDzdaUpgBTsjwEEgsaNahRKr+jnx3dPVjx8Gk0ZAAp4ZH
WI4XmypGm6VnrQAAvP9NE6hAk7jbEfA9YFvDiIo8augST92rXzGcAlMqkQIFXUM9a4+uLSjyhLJa
7jSDgyZCkBUOKudSMHsv0wi25awnpOTzhMbZvjQXoX/DIi5LhuaaTiNmbyYVNo0nWuQsMCXCPrS7
ZB3o0nJMMqYLFjT9LCn9ewWAMEC/BYmud6d1r6T5+iW5n9m/MB4z83ip9KltDNAq3fWigP5uh32q
UiALDO/+Nw8SRly7PQdeEsjDYcbdQeXuu85xdb1Ly8gzkyr1jKRkNK/R7Nth22bf0DRUBLIAsI2/
/bfluPyviQ+ZV7QyKGNrCBgepQ9FaXCdodorFBhRIxk1HjlOv3QV9S7g/RkhZIO5FB9ehXWdjf63
4PiJToGUOTlXbdnz9zyNCIZXjqbn8BdKkzQyxwmw6BFq7gTCL5960mMUp0CrhherhZO3D0YPxpoN
PIt/ljWfO8GEInqvWyS5OJR9sOhkTWX/7CSAD7/RZorKYJQXNzgdcGmhkEdjWmsFa8snYtCOcW0q
2F1v92SiprDNcQsFLhm9txW/RJeziEGoPA8Paxxr782NGI7Gipe+IJLpbxgSjWPpc0ncDIYhEXyG
fGuL5VCl4T0x3Z2upFdT8MntONwLTfUNz2DZgSrI4xQo/KllOMPvZZQMtEo4T9h5daZWFyAzMTXh
4yBDyybl4FXFRRRPrYRcET4HXEO0RrnF2RfItK/P+8CX90OQ8RhOkMgQuKzL17jMjZQ76V8soNFu
g1RBAZE9sY9K8ZcEuDlGQ5LJ5whkieN34Jg784YMkpduRWtY7G9gyTGhLFR17ugwXMi0BFNkxmaC
z4al+bQBXChRoe5jZu4OHf319AU2fVuIbq4HWpjlMvd2izopTx26m6C+3ZHtV0yFiBKuGiC+CNQD
tgIJRJOuL75mbB1XQu62UVB0wRX8Tfr/PEo6T3LXwUF2LKG/VqHyzd96dTqNrZc1I1ldwK1au/hi
WoE61609B0apkkV66nKIpjlPUYhddwMRDlc8QuUXLf7ynwcatiaOAmjFakxFkP21dBmNd8l8/Pdv
5JvPqF4e7nCKG0zY51Ykwb4ShCZpKTFgVTvneR1KWGgVm0NUJCsy4XTplMaKjJf4u+Hw/um6lGiT
UnyLIH6cr49IXe6FfrU86e86D7qwPWp803Ffk1/ILrrURTOvMZPkR1mpjgq4jErN0cDIwCOEpdPn
cxQ+AqJ6gwE9H8zjbtKsHCtgnSMMJglL7WIPAibbc5zGEbS0+agMweHbUwPSgbYqKLKb0FYUD06G
bnvDAfuvVjmx2X08SHyvoEAnCY2msfP19q6fLvyVxt5pIvvbR5+0NYEUe4ly0iJug8wzqrw/fPck
3bWtdVODB+k1TVyN5GeFiLvZbfzJfqfAiBwGc3VVpFAza3S9RNV4GkgRmvU4gXgMJ6ppqpAILVCN
2dopUaSYZffQUsVnTMDDnC+VBEtzUmjEMo+HOqdL9tq5Khsef/dYAo1UZuR/TyBSVOGxv+/3lKRM
F6Z4t3q3U4HtUnGhPl69avJpyhHLAlRU1HLVgWEfGrXvoYlZl3dLFcwyUKx3G92rX4/broRJ2SfE
eptEIJzzEcnVSDHAW0s4xrWufRbsHrmubN+v0CRFfMlcpFgrkKAERhxypPJvti++m+XrWcfD0b8x
QmMX0JJIYdUhkTdYgmydneL7U5Rx34Gbmfo0gQknL8nmrLEXpNNcepjP4rWizd0zSQ/gChJFwY5i
ib61pR07hq3XCYRw7Qv035wSwKBAZ0yhynz7JGvN7RFJU80PyuKDVUVZdrhiuWvBouYzBkv+o44M
O2Cn33r3WdoXoHdpkpJcUECBSbqgyHDbEv12HXfK6FiTAa+DWRtdo1B/G2kE1fPi1hFG+ozGezk9
bUFLUzZZNxrmmxs2h91AiM2l4FeXI0xAsarKgqQ31GgXccXaEKXU53G2oc+tTBbG8LpvCRvSY+Ht
NmOIxwAnK5twfmcTQoEySXltrkBLv1N/I68v0mRu7j8L8i+Cn3YZfUVUz1zRunceQYmcZ9VdCq7t
Uhc1X9LENmb91DTS4PZb4Njex2uUZbtqF3Y46J55GeFDotcdCKMRuNlMg9eD097euKN/BbjMDTjb
+nLe9dAgVr0oM1mZdmLvh+ZkIxNWRmSGkgZXY2f1naRs/3BFkqsFmoBr4YETvuqe/6Zo2fCJz6LD
dRexg813j+4fajX9S6MCBXGopruDVqIswTKZltoFl68g2UpJaXCffIbyLA2D8gz+x7O+apOUcnrM
jrrYKYY4F+BYgJvRLxvgYxMYXJ6/vzlnmwhmID4Fv+19kuRrXeeZLUllJX+o0ds2o602V6HN8zdB
GR1P9JhrUUeIIdxVrJGBvMtiWqQIejIoiBXhQEjF8Pgl19cO62fQnPamiTdQ4cuiwMiuEqa/0FDo
ctv61UJUP1e8X9B5bKWp0ioDZt3pcPRvpvF9gRde03mAOZ6sv7Dsr5KUMup3TmskQrLTpLLD4xHj
aQECl5GtKvoAB/Z8DwO1PK8gjoBHAZ0zaMM26luHbKuK+/r18Wzq1gs7zht87ElHtbJctIRBEpdr
LWtpa+elh5hzs8i+qE62VBYlPgFowtjhme/TVVGjwZaSDo0ZoR0nTE8815EZRYAd/zLqbZRy9um0
BoPJXaNmOhDFUkPVHVP0R+eD/fKAWAfOCOD1INxOk8ctJItJLkgDogENdKKrOXZtfgj6DpPSpxw4
dlWAGdpM1d7VIXyasJz1my2/4/Cv0Bq+rZKHy9/pbR+60GIbQB32hFkR18XQnC/HPcNNxkbV8MYi
wR9vi7RYYfQNLeESeJs0ZDyEZk5jY8qIxhW/nQv7WAShsUrudx+RQt8TLA0j+kaAkR5XyFGFjeSc
jtoq+i6mXQFzDE6QeeDyyehDev3cp7JxlUxVw7RpGapC6POTvPv+MnTqtZ6YDCT21D6LXyGD45dA
CfZhL2CoK3uHA7S72QtN0JJWnGAghyhTFLOK4psP5xvWpPZvvqqkzj5nFIDSXy9wIN8bVSdF5gHc
vnN6Ap7eIU7QvFzbV1ERphSHpexodwQDio3gbZdBl70wMiXDPjJSySOoL2hxPUA9cKUC13OHcdBh
8FE/b3NSNTM08aFp/ii/dEiGC2/nXGwa1Qv9KFi55nE7BA0tlmcGYamhZPyAuZVi65Au+VqRMbFT
IxCz2u8UopNpyTk+WiA0fwON5pFb9/6fFPVGxLvYHcpk8/SvFSvkEmbtaWd/dMqsMaBI7eWtzU+R
O8ZTgdMfm6F9G7uwSC9pepHtCjOo9UM+vvK+kKTj25/7SsVrlXntwnYITMWgGpafAlb2mJfx+HSF
cdu8WauANhczhO82BE0CcvA0gJq6ZP6I6ac8wIBlvfot15VNdMAI6SBiwbc6UL+bXwUoE7BakoGj
N/0D9c1ebqbgRwZGFsh04hcsfrzCTXiBp7HyGuwiFDHMlxDxknFZmYBg4BCa6x1oCWbFvfZUkuPl
K4frK1PAcQi1Tq/7sRQUgsLuFI9g74YfF8RR07rP2U0Bd5vQNkYijE/tGrrRXMXeXnu/8rk7aw7B
Qlk3noA6e2G03sVIXumq80/5tNEhvWViYE4KPjGiH7n3iMkze9ZZMjmqSGcqvjaNYtUOd6wsZdlT
Zr73M66Y6WUhqNg8Xe13hG5gVrpTKJ1JSf80fN2SooqOK2yG0r8BTAMo6XkOsU1DVE72BHvT3jPW
bbrA/ULxw9Wy4XI0++spse7gSIqR4xAEfYpkBpOTsHMTG4rLtmRol813yCof/RK3X/2NgXJiw0wT
3emjsnfiJ9S7omA3FZepmC09MV3kBVU5C2vPJCBGcHIzAILUfnV+8M26+LCXk4ts1kjy6bp8u3Fy
phVigM9K0piHoywzBM/mS2/VHfwdXPfi/UGYsHZZmrt8dfBb3HqQLCByF9f72a/ICvwI+FyjRpua
bFyl9KFm0gCuNvV6b0+q2TlsOG3FmjkEvbOaOg3w9DZoaXyOkWXh6NPSHk5Fcxu8bdbaJ6sH8sI/
zXnoKtHWdHvflOHSpfJkRrtXeSxkh7oEks3SfENYhNREDIcNN075i+05SJMLC0d3PL3tBIuf9YBV
5EOs148Qgq7gk/gPia6rUw2cpKKC6F1nWf1JbR6PrICrjooR+oE7KHi0bdhlM7Rl/oIK6wqmVbZm
rnVFQzuHZQQ60jVkDPwJDAbIEgDfcBql/JcBrXEvEwsWA7A63GzZGHVj4rlrIhDW169vJzruxBjF
62sSQ5j7//koySLFS+/pyi31E5qoy9gVXBaDwes2kYb5tlYSsFZtbISDQV3hWIUSr9BjJkZ7XuXP
EBa3TRmCuurQswP820uXhi05BOFhI0X6b0TfF20qU9LB7in8QlIFKxwP32DSjSaluFOx1Kv4Q3OF
bn97UhDuLnRX4PSkzLsQQ8vD2SSQaFU88krMF9uILh6uy+VN7zd0fuqBr9w1PT32xQhOk8lhpGhS
5JrgLoWRImANYVihRddZQmokzG43/dgcCh+TENPLnUG7NNiLDCTtoWbkYrs8XsvfuGjrdQpWdt90
FY623Nkh3ezHr2qhdaf/ndLMfOSkqvCP10Y7PfXwKnFfN+EPzQlGzT435k5G1Y8K91jzOsIoiMLd
eG6qlS/QXFj+4+GgqNByMzqs3ibV4RXc2NIzOkiNABr5T6OtXYECWs5O5ZM0PXsQ7PEbnK6SwkZg
Wjh7fi//cO92qdaceFPnhpPu5v4MjxRaltw7ydeqldNQC+ETYt5ORrVXYHfvpNW0aSOe4yjnrEHp
oudQZsxcaFHdmvMHHDX40YBgFifbwhQT/RiCWKqFe/qjQvDoxT7GjYqqwu3AZgiVIEjbnZUHLKe1
GJHhui6lZHTOnQZVAZ1cHpPwPVEEhH52+dDVsbgNBGDYi5mzFkriVEx7ZzVJ5OvNK9bBizcT8gW9
l5gvjAsIKK8MI8MFYEkLluOzyIpJncCxyT/X7s0eI8MmfF4k0ZB5xDOlCFRikXsm/deU6wAKB8rl
0qUDojx2E5Wd5BSeQlo+4fXRh0LRwwJbVzMXTFF42oi7sK5VNsM/SgyK5G+MXm8lOxpSQOCv9OPy
m4XyymM6LNqHLRaQsbRqQZrA7rFJVSb2AjvDIQ1KnqCADWvMhkyTXFUZQJBxoSKH9RFZERkpH5wS
dDLe1PZAxQKj9BtuWBbm+kJjhOGEobFZ0TpCuGeXYnTmkj2RBVUCgoTnBsSWIgUxnNcSUtJ8tj2T
jJbHqQ8o5DZlqVGkU9GUgpL08mzrwtkw2o3kBpr9VaaiT+YDQIEOdULsv+LywyYUMrI9PfMqEaVB
Kq68crFd/nGukmbiEpfHP2m8ao2a62vf0/pxPIWTX9prpQs3GXXUGeXm2DMItbqScKPoZg1V+1MT
oOM5jogCzUe8vrM1gX8PgYfePvXEEDCPVC0J4arUxn+xnMpOXLFgW651pJGOXlYfLB6fpsLLYujc
hVyQYHUrVCgltXbbtreWUi9vz+UaoGcJuCDbGZlCo9P+WSztYJKErCX61g6ylsevfa+Ym3nDiotZ
oNdKI90AKX05L4gke9ubRtsQ4y6s0V5M1H3w2hpjWS6jWznNsBRpHEZar3KTi8YBeS/UxoKPnu7i
LBHqoz8EjV6NlfwF/2e4gWSDeveicgDXJh6h2n7zvB+cJmMaMEuUeJiABhUfndnM6QoFBBEdsyiL
noRZHKhJo2MOBf9PoiiOZAUN772gLz3jGz8CzUmWbWWJWerjplAfy7OEdu+MU3kNKuxLy+moaHXP
VQvoGEAjF5BXHm6oRg2OxxKM31pDUEUfbdqLUqY1NoTMzq5LYVW5++4Mk/3mNFu4EfjITZV4VLjc
8FrykWHM7RMybwq95Voxsp6oYfrm5N3vuRI4gK/ngCZksbggxHngbAF1iFcaSq549xjLVN5LuJD5
rbkaKPB7RnwwykJpnNXCoBW5bvExAx9C1rbVsjALsZNNdGzNDjmL+vNt60V5gxKeOOi7r78yfapg
AGirZcog/EcTNLL2CBG1nmT1muepvCzN6zWd3lXTLw6A6JnXtoNgIrY3YeIArsDLRIT6HBSlr7bx
RrJHqtwa1b0UQmcQoVuefFywcdsi6+Nosgiegms2ac0/ss0QVOHRw4qc1wGzam06BroNYj0fx83s
OyrUQ4TLUWERj2NOaIGXrpEe29+u2m6yvGRViRe27W9FfBiWunhB1GKd4Wo084z54ykCdXqlzrsA
2vhNVPBMgLFhlNWE5Dq3KaBICWjUIsZc5tmT91mbqx9AM+X2ghqsHoM3c721uTyrdn7Fcy42kMH/
5t2DKlQIhHOXfu5meEKsVMTKfDQqQ0lolGHBoN4T6vY2XIGBXjlfZzdchRIgY7intZzJa6thKmIJ
tyILuFfYqb65RYMY94HRq90/nuRPlJo3oRiWiDOT/C1/HhYhDdNSj2Aa81y0hT7yQtfZmw+l9SHR
mk3ycuTDIrkoyoXImS8ercnmn4UZCEJHi+YL/T3C8KR48PueLlBRWDrL9txgfRuOeY9EVoNo7W1O
4hp8Qg+k2aEA49NR7bzLepM54WvuYyFVw8qLMFzsGZTUdYPfrujgMCPTAnrLxuQmDQA1bKBNPZY+
7RoZfJFkXYL6+bdOt14srFT3Bgbmdf4VGXPli45RR9foxs3x6Ao/HzjP55UuXmVsXgKmU0f7obh0
iSWqSzUMx060Wpgi07ncqZ/Tk/YoShNjTY6a7GaEXI5al8+VsOSzIPgecDOS6nOvzorgYoEuBxj6
siZyYrM+YSYpp+mmMQEoTwY6oeA2LD7DCM530mlQY6McM9+6hqktuwNQ8/ij0HCaP73ZKbx50eZ4
/EJpPingcbD1dosF7QUPdPTIVp3Mlm/Ga14pbg5KC8qlGo0VSQsc79lmmX/BkCV7oRdP/LhplnA4
NBLXjw/ZNUkywHzpDvhBd1Y1X6sVoqRQyi5LHpzYyVwfaYp9cfHTImbkKyXk+RJozrZQDp/nAPAG
4at5JZdHUzrHO6i38rbn1RmlPMjDL+PdHtrlXvLJWakmKzeK50FXwNG4IQu7LKejjllgVAnUPxVk
xAXBytzHSjaVp9C8y3OLVjjhOg1lXCgrmopJb3xUPsx3cMOjdmdni/LlmxauRYq1i86eItDVCYsy
Tpsb46IJBiPgtiZTNB0S+XabomBVqpVgbRtnWgdV6AfBOB7BaV6J7TLPnYUUzVpnzuwAvw5GU9Jk
KPqGNfLDAeHhUfOMmSkwj55k+p2niUZuc6gc2Os5k0iMidrKOIjYHbyN2rSqmjzFz4ULU4PyNHYJ
2jqoG+j13CVJ3u3tcO8jP0khOae6GwsT2bS8oTXYNpefbSu4PVL2HWHFi/j8x23Tnf9TfJtnXDHB
gZjWz9xO2OhzE8cdZkMkL/vhNarGUOA/wNqKRniWD4Cd7lkCDjNDSZihEG7TLEdcndCj4rakikoe
D7/lN+NG7q9DDush323DgZ5AqiqsTLuDoU7nb56P27gGBfWTh4SPFTObXvaevSxyNQvU6veMftns
BZIgFKJoz8djAL2dkeAu96WLoLAAVAdyP28bSA118ll+KsUtvJ4FVqGbaYS8EP/2G0+1qjzb0q57
8rINtqvB3E/JrLFgsckf4J3zMgSYZsuy2uoOpkhsVlQ1cRKfxJvwCrrcp97gK07R7vqMo3TIaJVR
Abigtf7jKCW78Ji7p+8PzPv5AGkMlnrZVan0lKurmYxnKK59po2SXOwk3OaDJElEpoF05KXHbb8w
Dix7Fdpy5d0hTNxZn41umLyHn/q+EP1D5LtYfkoOvThfHovmx+WJ2Aj/bglg2XMz3bAkb7Bx9J2e
pb5XSgWIzM0sRPhKEJ4zatfUl7WhJY6oIraRNu7jM++UAN7/x8FD9ZNiEE/MSl1HjPQB5z/AswYG
aQvmfcxSYM/w0aE/IbIFCXnX+smOpH+Lt+PcVGa7RkjVWKEDJb4Nr6fbXMtNh5jk4H8mzkOKZs3p
7wV3Hbjo5sN6cip1J8HiBnV3gDZpAtYyBd1hq9ECM59E37/QqX9pnSDVopKINKbJKbWpdgPw9kpf
ZQHqSJaas8t7W52eNkf30wFfMvKChHktgnbL/QHyBmCk5ZBjIogfLXxDQcJVFVomR5Z14p3WaaYL
5nm4530ioDoR4Lj/3BAgpM1b70vvWh+Rr+29Zt27cO+9uW80wv+Umix+E8JFw2xqT7olv56/C1p1
6B+B+7BdaRPIT8C2gCXDUAJ6P1VHrJNEZ1YKW4p5wDoAwp0BwYDp1X8aJmFw8WuKRcRly+TiLvtT
LFumot2rBfdUxGU8rgsAk9aaUqbjhUmorkI9AarvPiPTUAPiA4gZvktvtXOZ7C7X9w4OzrxBhO38
7HP/53Iw/k+9E8GC0SBxrkv26euGQaQ4Hv7luPjWtFyyXZNNj2/q+8U0gc10xodEA5/zvxAECtab
YcSVcrlKfet6WpvbVoYh1w6mPDkO4ycUvqNqrmbIobAoHlZrhqCA8rYXLQ1ctSF+O8LGOBnIHmWp
FAg53zQ7AeQp+FE3aqQitnxNP772bjpA1DiJhK52GMUwZtGJ5tkKN6KLotilEM4ryvPKlxH5/xES
ONnvgZOP7nmcvQaUjt7x/SUQmIshQiF/cdy7QdnL7tX/12PJbRkLFFK71V4KAmoSYKJVVTH3143o
Q7aBiSxhrYRlqaf9D+Vq6L51HTEbQvU8tW+Jlia24mNsIECT9V9E4QSMP3V8GWerSef4OSoc5jPI
/mBJmmnxaV1oTBojEOVhmjOIWpQw+3dDEkU8Ei2v6Ec09SqWgx1sP/MTyk71gVNtSO+NG2h+B9yn
rbv52muzOdLTai3swDUoBUuzEpOUNUYAdQVhDTbW0EtJBD1UurYkXSHaPzPNwOLFwhQRg7VcuQfZ
SgqKXezaSQ7m0ll/drtDpZYx4p3i9dHgiSS+RLqsmUm5OQaHXXGG/4DmPxVqo9W0Oy5OOFnMSAcQ
gviVI80MmqXLdA21rCrELB6yNwisJ0TO/uTRRPo2DeFX+qyvyGE7r5sc0mn2udZVT5wGV2oyeENT
rVVzdOFI638DDWgF8IZ+iVb0BWnHTm6qcG1kVG9+YgmyqV+U4eiNF5oW3psLomIkVFbLr0W2vinf
KBZilEla3bDC9IdSc63RgNp0QziHIK+2x+1268tRNhtJrgeFwWKcgrEybVYIPGcduOIcH+WGjlgN
Qpme1OsYg2kVk/w6RTEV6pldT9L0ZxTGccz1Iu1QzAnN9upSh3v6rNbgNV2TGKKH91q5zmdWxelV
2Lo6Adh2Ufy9rt8D6qpENP9UVF7CQ5Lm7p1qEpv3OeYhgzzQMSlptfKCrenXkKfncQwWOOLb0l7d
75/1gxL6IxAmFif+FdLlL8hHP4QE1EZxHjIisjk2+if8GNuJSu9srQ22E02yFkWGGvI4lySyonlA
RC/hQJ1eI80tAOG+1jAJ7WgDiQftyM+/zaV3xSxQH4i8N95VNPHff70MrpXiiFaKmi9vO67pQXVy
JrsdWmu9cAvcbiRdLcfPCa882L/Avv4pIKIZKpAKeQJ2bWrJrrMVdf0BpQft7Li9HhMTOpjPPg17
dWOsv7L3ghh2lrpavPNN5TMDdJBXOrWp4vzHNwtGhF4RGPD5FawavSSa0qCJ4nZ+7TaFlZ8fGOrS
qalfNVEwZh7KaSzLX3emAcG+O6d6GURsHIznexU3kTA4W6YjNgdWcURw96yLU4o6bXEqJKP9roeS
/QjTQSad0YnOTUyavnA2lpHFawPgwh12tQ+uw+AF1H6J9ihA2ooV0JRDbLn4ls/quo5tyFl2hmYI
Vb9+bgLVaTiWW0I/lqwDrtO9A0N71ElMha+vVrF3muZQAgLzeIgjK6AiJPikWZa0mZDa6wdqNNxE
Mlqdbpgr7UpZE3Voo2jPtDl40aQPgRUpHj95XRUTd6J6c7R7AgkuV9R7axEz5deXVnVe7JAjGq2M
BDXbax4Qjg2qR4iq45eEz0/GBWO6fhWZFjcka/bJj8K7anwHKvgwftd+fYf24PvRVlWi+ulVnk8D
GhKY3zrxtzmuxupjiOdPrbUhdcKMfWjLpkodDDl5vkPEuKcrRkOdAN8+0RTltcluAJtQ+ZdtvxTd
BhjCgnvkBjNOAgw4EOj6v6Jmc2E9FabJUfd1/yyMovL+UW8Zb2rQGoAMK3MyoitTpJ7bcPck3Jax
8bqtz6HY5F6iTv2NdFGrhlu6e5XJ04QAw3udDpaxJ0RMKKrQrhtP83/igBi9Dbf7WsQcCbj+aTL2
zdvdMtpDbThpUvGquiEhcY81AFwCsx9SoMWZHWbcBX3SweB7EebZ0GhqTxJ60Z4A+58dA90poVpA
fqJM+AyW0k7+GFHQ3vxL+XFeX+mhJYQSd8Qf1KLn8Cqj6Vt4XYF1fzPy7sVFn5DAzZB8Qj4GIV1+
0Qu7idgjIyok0CtLySfgFXP77WtbsTK4y2QgSA0MMMyiJTomvpNW4TwV2CZi3oYxqaxqf6mXZxNV
rku1lQUgyBLSZR+isQB/Q3RwNEQilGc/jjMdd4qmIt7JNNKNZIYFzLxJwM05up51mqOB9pxdx0El
tK3Dwj+GecWW/MNcdjB2/aDbhkGtEVtQ2GKSLdOhOMvYSmmrHGydf3WRrOiNC5xQ6JK8LyCJUfLQ
zX7sNZQzr3nyHtyoQrGnEAeVfkzI36EKS+rdP+ppY4Smbf9NZtCw8NkWbFlsNfN8WTSsI/ihyUIs
Yy5fgnfRYEhQ6X+F9OorWf4HxIUgNwic++dIxE3mAaQIQjn2DnLuEUOyv7LItt5hTOTj6l5ElpPS
+N4nlzIq4e3TISOuf1Bd4iP117aaqZmduxITI1phGH7Ov7hpHSeAZw5up/6NwDGvMQkvkoxLI0uu
2RNIHuR+0/5aosuaXAgPGB7XoxQAkddR+Cm2HIPR7FR2n94QNasocNCdYDkK3cD5dcLlbk3m9r24
uhwdtmANm1/S3AJTq71Kp6OHi81ItDe6HeA67GTClQBKx515jtE28eLDKup3NCHUTDiaLVwkAJRW
MqJNjRW9Jr+zjRpfC+rwPMdqXhVgLmZleuMgN3bPoB98Ku5Gn8HEh2jB+NdTLTfisPUbibouWoYA
6yw5n7N7fiDCd8c47+QS3+5kqJhChxvMYaAOh/CqRX86DWYQInufjxKQRLn3apY2Uju31GV/EC+c
6SYTW2j4zSlxcWzJhsoT25jE7d1TDMtEsfaYFLQ39YcNQkQ72gkN5FDOi8T3LCsDRgycyTRxZJnF
nr7mDLQinrX71ykseKBJ0wPnJdv3Ee7iDQpMG+svaT2+PC2SRpbLFHWy49yCBr7MDws+Lgh2V7vt
MGeCIBhNYXtoi291EH+c0SsNduyijKKrIvl9JeoHvSw8YGP0Kibv3XpIA4isrVyCMiO8wbMDCFv1
XJrB2sYNHjEsT6MWWymtSfCLSXeC0OluN2V6Itbd3YvLYY7pZai7QbZ+uamD08ENbYS72Kr4qhMK
i36Ri9qQAdYTXd4sANr6H22QyqP5nNT0KIjxK9ohnPMPP1D8dRY33ih63U5y2zMFtaXcMH/239om
tQulNM+w5ijfDZkM8fVP3nyedGnWpY4vz4feesbsQBT6k4Qbes5jtPNw1xqYkYdvWBH2g7qxbgVz
FziNQm0c4DOwNdYi8odnbbZJcszl6B2H4TOzhnsCvoClyAB99MJvzc1sYH3LGwKTzcSOeYOlhwui
qzO/5JWW5QLmISXAoM1YCYP3Y6wQtcakthgBeeZanbnbk9CddITVZW98X9KxcZFZQkl+jNxRQQDi
zl9QPJeoE1HKWJuDx7VN8k97S7dUJ2uuKDMz/ITmfDUiIjXNbAEhhcr9D+KDLb9uz+znF0Rh7kii
Do1dI6fjowB3YRpYeq08W8zyLeuTufhXjBdKAGgJdmYUDctrihJSaaWyVIB2FXD6/hdrE6odECC1
IadaDds81kOIguVMAfB4SiYhRWViXiYWdZQzobi88gg0igMBFd7FnY1LEQc6D6ysci5m1705Igdi
hVHXml9vxxc/e0rhoqgoTRQO3cd87WNsJgri+yYee3ZsgNnfZwyUQmB1QiLuj5i4EQlUMOJwdiol
jSONcQl+TNV7il3KRDARzkZemZFhR5f6CMOps/MF2ygPu9quOF2pv/Qoz/MpdTLoRL16LlZ4FQ/p
NaDih9sqVLFMuW5E5XXCAdZRj8MA7GE6todtUlNKC25t85F+soT4bOmtkBYXoWAiw8In6RIVOHbh
//y4HakNDXyiY4C89HdN6oDzS2qnG/Qc6ad8yhjMTzFeqlAzNd844rE+3PNiiLBX9IDE6vrpCfBb
2I2FQ34fuToOJKlHOM/8wf7KfPFufB/en4G8YYC4xhVsHa7eTHvbh1d1dF5oTYmywrVtVQbEdupO
0P5Pn26sdu5Dc5gYbDJQcozfXKj5VCrPXrf9H///IdYyXpBG65RPSWtlOQXIMMmhyvj0/TEARth6
VmSSgx3YOg2Xx4Fg34cSGlbZP5A1pwitV7/VXsFYUQ4INez7fS4uE0t88P2xC60nvSqp5xvvJDkC
zyVedu1BVJDM9xS+dO2PMCMBgxoG0LVA5HtIAZ9wxAMr70m4BVb2/ORzu2SW1sp3pyXKHtaXVxhk
5VskLAN4KAMQZ7jgTiTxJHKEcusfTFbqgVurWVWrN5swGka367JgHINZ7gncp+5l9HdzH8CF0Ieg
ewxPdTjYXlXTPBQSDb3fvjD7LLmljYaQF1CQCzxJ2T8uFGqsnCCJM7y0FVYMiMKsynJ2UUVCEgnX
MM23QvF2mCSS1aIZ6sYMpu50Xifk8i0jDQh0X51a0qgcywdURQ/+fkBHf0vOnOGfupmLCWTmgLzu
9gXt/dZeuMde2+tC0xVIoDI0fGn3PHpcEueQ52iADKqMHQXVh5KUJ4i4G+t/6s0HESEquqh9Ns+m
c1VNOut9zsGLojpLwSBPnyyPrgGYuPUuqwfmr3EOGnZSgKzGCuG0FPckqGTffPyLtyxz2VvaBYmq
BFD936xgAvMECHDrkRplipdRB6IKmxdWtW2azCKO4zVbxQ0XHfMROJdkolzJynuMgNj1vOxfEuQC
4PxOvkXUs+jzHrl81PB8Uq0g9l8SC3/HJSBj8vpyJNgLG/iezi1P941wuvsodMvwFHxEPtQQ4+HR
U7B1KAEC1lmEkPyfYh24p0PKbMebr2pIwy1xmzp/TLGJcufU93UM6w9X6BbCcFUonJUu09eqeTbU
Wfo8WvN3ClsVsdJLYI6W2ntRxr5cdl4YA9eqccJb1aoPkqcRsDzrxBwhen6n0wfF6+JWXZX87eQv
3sCXaSew4JsHOrVE7TiXqUqfWUjLJpok+SOJRo8CEVFWkKtHN0jeKz9uzHKG9oG/lWFJmJwXWMH/
49NMwuVJ1k1aSA0TtkQiwiLj1hibZedvmObyGzQVovQdTHqVVfyfAmYZH2FMzfmYxt6V1tpDW6E+
bW5+Iz2Ek6gEUNa9TvNKIf4VUImDe4ek+HXoJu4Q3FbTno3F28LPzAUCF1d+r/tmAPuAXfOYn4Oq
iETYWZRSsbcwVCr4dZVt8exZu8Q16nmnspcCfqXyoaB2mH1hDVbRh2rBc0g2ovsJhR5bEXRZmIlL
AQflfSn/vRjiwKlgfxPSDPAkf0ZTD1zvVt4VILR93D8MVwyxnTreDbkPxR6zzOqsYdPFBPJJWYAj
lwWfj9n5jLc7JKWMGgdDKiyVbWYKAZSBoJxMcjjU27UqWwVhTsa2cRLT5IPft+UJX/RTC+KbLScK
MSnZ01gpxXLN1T5dgETvgBcGZogNXhRZXPESvNOhZvgMQY0ip2kSuXLu5tDoXWcpeTfRvo8X+TLi
JIW3bfp6HSfJCP8KIt6C5/DoNWwO5dlrI42cp4EvESygZGbXhPidg8P26VKUsFzYMhUe9+ns9aJU
N0wdpwqC9gJgt4hU/MmgXAdtp9aJnmR4qTUJ7hhNbpSIBTWB+FfIstsKN0AvTEGj7cQJaTaJI+/W
X0HG9I72j/UGFaqADAP7rqY84nEzEUzggdAwIL5MZXPbYqFwbjsYjleE5yYna8QRtbOtOyEJf9HN
rRk+8NGgNOvCaV2crS/hz4aXBEBWgnXlnKUSlDJAFCDDY4mw4KRjGx1CF0CBxGqaEzNW/FlK3lgA
j40mXs9d/MnEtB+ZDEIsX7KzVtpgTqasHBYxl0LTJyQPvQvFsyOALfynHKqcrc/rhEGEkznsvBmR
G5MK0XmsiZecxLgEAq3izoUiDajb9/zYv54iEydV385IiwxuugCwDZ30IXb7ZnchsnGhRIG40N4W
/5GFEArzCuR2SvABkndZ5DrGP1RCNyTzKu+ajsf0PrQQ7gW2EZeXtddlYyY4jiWjEQap27Mipmlj
n/O1cgyI3YDTviQoROiPw0BmoFwDkLqslha/teIuzE+l5G+0HKeRZcp31Wla9iahyleOsenFLWj2
GxP7majWYmNOJIEPF1GGpFPeg4X0WTxtHslGYB29klF2lFgQrdhpFIrtbkit/JSBDzr8EiunMScn
Nq+LP2Pc/KF2yt3L+dQVfdk/FE2YehI20iBi9xnM+f4cv0x2Guq4sDkkSscVtlH0G9a4zi7eXVDV
oyJXEAXULTxlADPJML/j/tFyU3yrmOYlmupaWGK2UawTPzJlHqBCBx/EPj4cZptv0q3rKLMT3tQg
GOc4BAWJDOSEyOZqZTzi6XcVUnA5yk+fh50jGVQcIvVic361Oqv7BqSIDbmM2c/DecqCrWlTC49W
LtLGpS5eihIrof4wzcpDLPbfgtBmAE5Y900NicJnw1npCx2qVKOiPAwn3dUx3MHRTsnXDjkpqO13
ay7rFyOUCuaot0apW8/eC2rorLsyMQgCw/Y+XrmIxvLPJ16y2wH4De0uEnxM92xwkjgcjgs9A1/g
/62IAYgUG+fko9wfpWdDg0XWGjo84ra2CHxxfyC5ZMx4hXxAmVkdX2AlttNXdwQO+7/q6M8u+n3E
hvJapwZLbMwyDEFHV6v6p21acZ42xvYCzvHUCQYjDNWohrKImpc/8asmtSPpOo21bhVswJW4baCx
HqlLuU3G2yWmcvAkqWtrDdJAKM8hVdjDOgI3flF1rcC8ZZlAR2F97mc/BSnBOwqGLZzSwuEnRPkJ
39XIVUW4IQK1G1EDvK6nDtIjxyD4XR+GSN9SGrk7CyI5BaXmROdaoXfXfG1NCKDqVNIYZbBgW68i
6fK89dHVGxYs4+hLrW6aemIOij4UZ59oQO0hnlWMUaP2DiKiXvQZ2R3SwcsCErdq4sEfKyRnDKrl
/4VFmGGJM11Zn18iHoqjlhMokyL2c06wr7aFaqpB2sWnl65fXgU6dphvFqCBa3CB6HdAbol+fDXf
6rHwAjI2700yta/g7mu+1D6M1pQcvEVI4I1V/gZFy5pNSe70FinpxbBzJQNz+9tr46T+dNsnD9iN
rNWJ1ZMpsJ5Z0SO9fY/gR0fntuYtbMHv/gZaJ/pZC0uP5yk7lb+jXGP/j5EybNkuMTVXEKgt3iKG
jxXYc3mZcCBMCAnI/y4BFDauvxv2DkuA/iAheyJcHQD4bLU3Q7eHohRj19fS0kcOcgUY+fYtUtG4
nAcK4m8u4+aPSDsqmand+WQeLbmHCwIDfk40bWaLEbrzMnjUEtFkvGYc9o5gSWNJvIium4eBDWZb
dW3lrKlAawKidrJ3bPHYuAgaQvGSfiqaEH9ktjV2Pl5QVH2hPNRmZbROq0qEplT7bhivKsJUSyZ4
4XB8RxoorWpvzVcivI2juDfG362PP80zMHxuyTn5Y26ek7mTwdfrtCkdc8x5s61YVH511QKXnccb
Za2Vh4IygSSG+/9p9t2BnKz0XLOPUKiKXe/qrSiJqyBRUxDW2y4ITXd/7Z/+e34R0L6uD7Vvidky
IiPEQMpec/DPjKDn3ZgEyV0czZTaLqA8Cu1k82Mm9LAJITHVKPEOeO+4kDfQN4SslnLywCZ2bx8t
seEy5QuZLXp+OOHGVLVLhU6zNROSk2RMZpoMR5qnp4STIwOUOAXx6bKXGZdSQA2U8rSNj9/3cRxB
hYJB/jNbuFk1g8Up9TQhS1+J0RgG83Ll4IpLNeuAOa4/0vbqyiNJ9OqDBsj58/+6Eu7lQ/bvyPT2
J905K0h3Bh9J5rmxPdA7ylT9o5Z3RCNCimrENRrEqo11qxqtHNOSEitMARgwq99vufLnm4Zy+poK
yziYxUxOKPcP+OV6vAYxVnw9QkVCjQLWnuoBnoCjAqMqAEaoiacG98E1hyg8PEZ2M/rVslC3htMZ
m6DRhj6Fu+QEEAbs8ynTrb5ET7UzHoo7lgJisLz8iiqGpdw/wdL2EAy9QDbm+5DqnZMi0+mqy6Nj
1nUtNFxFuzHI3KglYyRWedzyuEOy+t+TjLDPjqZCyava+PI+7M1zhqFcg8U/eRNuuMUatCczj/6l
13bf114tfhepzZVKgSFj8TfLNOUVSHY6pxMCYUnF4CTyI47bn+SRoaBewAy2FYEeCgiu0NjxOqSV
hlPY3kqjW/cP1jUA5eqva3RN0vIIFSBkxLJtD+zEXMF7oA1tyNYXt0LlChmn7jEsP2VhTzvSEMYo
nU2mZ8rCcdBP347PEk6MR00o69nmlz/Yd3YEPKe1FI1NNfRZw9MJi2msSfzeyFHlMw7lWTRnzh9b
ochX26ZyXWxJSPusiR9ILrGXzX8f4NhAxrHeXqouuasn89EwyIRxXUecTtLU3jVw5ELmRMfvEoM1
1+MNPLg8AZpZ/R+oWoqWYnDlN2rZy/q7//N1MGRtiIRqwTHxvMa0eCDKo6wU73rUz2Up6RSo1xnI
eM2QjfpVp613noXZX3rW5Q+E0TnsVJBaK2I2zNHFeTL8ztZKHBPQwX2d7K5jMhDNYRu7J0foCmwu
UYgDBusrnfkySyu4yVnI4kbXj1wM8A6YM1r0A9BZirz0pxyj2DHKOdy1iX8MeBcKHJvuFW8/e6Kr
++vLFKczH+f7tJ9fdc8RqrrgbQBJa01Xpf9KdQ9G3fli6y7Vfq08WEtzbgEOYQ7hJ1YiQ6FHBHNS
XQIcALqXxO1Z5rz2w60IBvZ1B+lKBvoOC+mC6vpQB9rEiGvjV8SJfG8t1VgrrKwrjeezrZQ6MjHZ
/yi2dMRpZ0DrxVwfRDGha8oR4/4E+xYnMbB5TDPpxjWRaLjdQPPmcAOHy6fM8EIt3tENT2RXe3II
1vZX1X4wXdAnQzmRILVebfZiAdiG79q2W57of3CNBiTMwTICtuGtYgXCS8ON7p0BdKWx/kumXehq
ZTjp6ENT/codkMx8Rtx2pFu8KRI09wgDwDmCZ/7jHYaF0tpLBmUt620XQCYeSTUPySCRHI+QMimK
J+w84e0Xm/nXgdMKkw7iDlZAFAz3A6M8B2ToYPvMN8R5AXcEiqzIhYcK5RWFe3uxNvpcJEmgvqkh
/OlPrcg4tr8cP8N4NCtkXUE1WL00sDZT+mwXL022pk8z0HA3Px5CoCzUEAMDC0p5F/SGTxBT5vuC
l2lgyVuN7xGcB7An64wr5ItegjL6lokz2FjWKbfthCixw/WpMy/GE8b13/c5p4yL5k0/bX6S64X7
Ix/8PlLq9NY2bPNdSwqnVbF0FHn8zsuGCaUIQqgQEwHqRCUhz3Qh3W9D4R6lVKqRjECL8OwKXW3g
S+MBX2PoD6LyEUj6dO9A1CB8jCZTY8oTnG8q1X+FCzJmmFLTAFmQtaxoJg5AwIqN/qqN8OmMraef
plRd3xBLO38QNXMhCc4Nb0a6ZX4Wjb8+aKQ6OQLph6OsCpuAGkCu164ZGqn02qkxpoyqdVs8DHgb
Tngv5F+MqBIbweef/cyhX/ylNavuWN+6Sl2yEuxGPAO79cNPPB5FvkUHBotlIYWpD0//r4k1dLvS
heip15QXMgsNk92bJIclk3cjmW0BJiEVtsy/9hG51mZNg62tZV/4HXY9BWrfFu5irf9q+DKtXu5O
XUY3hR5t23Xwnz0UG0rEpW6wWjbsZNubzp+lSYaH2y6+6WA2wEeogect0vNof2By5YMAsHS2je1c
0vpFfOzl2pQQ7FyMCk0+kH2zQgidDal2tIj7Asq1jFOyLoRRIgc+RqLgx0VU6O8ksvkIkaXMLrfx
nvAVd5Y++YDtAMfla4ymBu9ifJ68WVsSsjLcbTuenTeeetEoSANB0DFMxAoCAa4gLVAN0fN11YIR
/h5i/R9lL7wrDnIfIsasw7UDu3oqVLE0zVYvS3mOK+SHSQiMFryZeBOXtIaiyV8ol9mp23YlNWuY
xqourPwiR7o13JmZOultc6+nTI/P8nHhRczKh2fBCZUiOqbyoI+jSIDiR2DleBIH1ny28vl5V/Pg
+eQ5aPgePuUgK15wP8Ms7Z/3AM00Cr54Gm0Ijti/JT1B3xQj9tqnOUyFP31FHp64o8jTJY0NJbr3
eQYjGIRzJnJ04YPGoB11CL+SEDcj1wZqMioRpJEnoh2ckOF9JFFnn2udDB74C2h8XwOZCctHIChN
LRoaMybpi2sYLsH5hjjKoWv9JyqiWNlL7xAYz1Ylk1jrzwBhQAxGa8RlLyDtWTq46gSZIBTy2EeF
Wc3kdS1oeh0JonilYFeO6WyaXLM8BH3pRwNE523vD86rgd3VTWzONL2UKxvIFIDTFunsXLS8B7sW
rcT5c02XNAQZVpia1FZLzX7BfbG/+m1BXLgfZF9UKgawfW2xd1yzU0i+hAEivmrUEJfbY1lDZACM
WbiFXHFgXM0acLiBhXimwJdRn4eb3ablt0j9fD9hdYB3GWo8FJtnLCClFMFuYpEjcGk1P0LOo6+e
dg2hBOHBe2OL2SLl+GbuXV4ThxOEEjg7bIfk0l5ub/mUwvTtLe80I9vk3WcmoBPDGW9c2xLrZycF
+YsEl1YFLO3ZCayx8qI9eV+Nr6rJMpgSlX+04AyxXapmRn3ZdwBcxRITwpiShjoJ7RzsUwhVqEeZ
iZWAf11IxgGksY2tb8u3DM6Adny8YWzf0M3TNDY8A981X/n+TLW6a/Lbc2tqUKyngw6V0zdLgJZw
AK7/sazu/wspJS907Vc23r7RAl95bj2NEDq9dieWTfSDbxtMT9MqA1qEanf11kcZgABbp8lnCN14
GgsPvCBvj+gdtRTOBmpaftvCenRbZucIdOMWh0cNtW3az4KnG3sMt/wnq4LpZM1PsWQMQ4K2lmzx
isEbXGAnMyF6fPChOvPGzpo44B4ZCRuJKmSkkGsSPlE2/TA8bai926aq2BrNFmilxJtakkUQOW4e
NxLb0TvRlpz4icCmE92pygFQshcMwibwH1XwN76SYDnQY1PRhQyqb7KcjPohnOKEOgFqZuskf5n3
wB6GaJ/jWJnNB/hYtd4Ij4KO9j5a6XtAsXcVu2WqWp16u06y9fg8Cnv85iQGvrmP2mQhBiBLnTbw
JuozLG7QsrJbgU+SLx7tZndnJ95nVdWvEtk4ndqU1/UGeUrxEYtOHL9UseLm/nvszDX5uk7T2f6w
yVn86k6yhzlsnZgJSZdZ9M+L2PM0LIf8F6GkAExFJ1aocY/a+gkRn91ZYQAJHbcfezHhrV8a6etd
EmIkIFieiPlEis/rLYeB2/ybC2xLYIg6Ju8RsslEQjcJw0IlMlWU4voE0SeF9C8bYN5wfqCfe5tt
wsJO3FZTrV+4jnxASHXcELZPMmHfDoaxbZh58fJoqvivf9HqcqNOgbbYfbwqesozEnb+9yXhDSX3
cZKuPMLbk3Bv55cmSBs93Fa1amo39R8KNVL/qnfvqgV/Oqgg8FesLJz6yT498NSYk0W1uZGD+Yb7
8cGW2ClfkcM5VZLb46PHsdcw1BbANdgjktoWkS+LGsUBL+nSgr0YAwVzI0shw20D5LrzzV34nmUD
7e/eQ44B/2UwpoHwPXhKHvenMQHtKKM82SajsepoSLOr5qbvTfg7S93oY5aBHSjrY4Ipwim46K5M
uXFlg+K0dpXNB9/qvoTxjzLylggFY1vC/n/NTVfgj+G+zgHEhNRf+H/3eoyk9UCXoSNfUnsjG4g4
HEQw5poat8WYhR4ghO7+dBS1wR8sNaHQrflhnb7bB9P1ptDU85bLNsGW0gjMjTeXFcmDZEYaDp+M
DMt56EFErZ7vX5dI5iEAE47o/1qf7l7Mu8RhUcvdiM4pvJp9H3XHIzP1k47zRtjrpI1sxudCBsTt
+QutbWTegLW+BmkbrGq7hgx7i1lWRZQ7pZEFYhsuC9f0bseipltHJKRxtguOBk6DCdw+boPhUa6z
QN77QU6K7e2m+OxV6CNdKuc7o5vtgQd2Aqk1RHZMbgPrl/Elc6VHmBuZFGKZqsjLsFsgy0DfxFht
8jDKehT0Qs71Yx6oQEgnS37iDxHkGs3YzpHKY7wN+6vlpkSKy8stGI9FgDg5kFHFrEPnZlLfXIqY
6mh4uOFD0sHPEL7dyTJT8SbaoS7C5xPKUGitkCH+g59vaW2HEC6bJQHWc2ovl8NLXC6XcIq9xsGp
G179ufwFMEbGpnhMvilz0wzS/0wcurweoyO4o/9rLCMMqq3IwyT7Vtq2W+knGxzZ7sP7tsUXJIJY
vFgoPKDMWBC7EvYCDCQDv9t5vK5Pgev4Bi2at6GolcXl3KWwu4u6RUzAKIL9CUJvlDx2gSKAdfPJ
KlHqH7Bo2HcrwLC1CMAbyAIaK9pWrEx0rzKh4CW1MYja+Qib3LbCJ9PebQD/NzmYsOna/Tlzcw9V
55Bryw13q4WSKYMk0vGGQ7P1Tjp17CGFwo9dttnNIP6DgOGVydCSAsf7uiCYVANfwur9r0RZtrNQ
DqheJPyGJ6giv9UH9E/NjwZ13oQjR/VThZ6pI+ENbOSUI57HBzL9wZGu9m+gwqEMJ/IRVE7V262a
xUFXdjko+osR3Lduwj2PG59895QoWAy7kan6tar/oP7lLiqSEZUIu5MFkGlVk9FZx1CY0PecUqXn
MPLIZqcwOLAtd07OWBfkbzzRjf6/YpVYqJ9+0jwV8mwHGnLjQU4Lx8xF1f2+uZtVBZMCzY2IsLYP
XavLSw6V8KnFuu5GzB961hRiIkFKAZIqdbzG6CTPK9UVdMvD3FR0S8decGlTIt7XAJlGnazAwx+G
W/tvEuwOHoNJhRczVNaHkYsLHOhwMG6ad4OUkWOXk1xiLocCE9w5uOdE3hyy0HkDv+dehssC3LrD
ytnefwntDpcdg6Xe9oN9ccbyO/6fk+0Ii2D3BJ4heZhWIhNdHxMwd8zwwppCtsRnLGf4EcQd8CzK
DUGvZC3MweQWLcR7SR4K7qWZwnvjuV5w5ZzVYiDU7GmH6Hcl79jXfjPUbp0Egcy3XyTym0GI6wZh
l4kLve3d8/jRbeXaCMP9LNulR6jtm6SYQtvf8T8AfITLBwyhRDP4P1Dd3e5AwjefppDICQdTYzzW
XI8g9de98BTaoxBjHLyQer5Ae52+dBP+qZHbiFOCT4x3k5ejiuHAY7qvUd9CzpY4VuAnIVXypNTB
bahJ6OGWqCBo/z5sS+AoKb9hYveMgEtDigtQMnxOzlSyaNXcg9dRSf4L+eDNzM9ack3vgeFSS7SN
g/aI38IvCoAwHsDSawJWs2fw1WTKS2u9hVUxn035donirwzBCIzmuk7nVq0jLUPuMrL0rbIkmOfP
MoXtovAFum2XGpS2gjc1LGIC5TAij+pCdAg/yZLWeHBEljvqGOZ9hgZ6Ke/pd0bMiE0nxxIVCGmf
9rFEj2wtC/nPvkBlrr2SXa74k3jXTnw9QfdPpSkMH87zFA8WqQtGeLUIqi5aYaB0CWsk0DK44RnN
ThCCD+y1+PVHgKgJ1Jj0SxXOCQI5AXk4J9h/Pcdl0K6MQ/xXDs2Lo4E/hla6QlFk0uxuhlvdutAn
T0QrZvmJloEfyFcZtfp6k8NpO3VlG/RuMYowVJlfnBD4w/vN7LVQAN1cGuy20Oye2c3LvxtJ5gaS
OryC3u8RaygdVoCTSKDZhLpqAiOWnr4e6eyC8HABHo9pYYZ84zPQ+zDD2e1j+Kp6kvtP/SEfCas3
K967RQyPDjZMsEqzXXacCRHuvj0ktpx5yMrbbNQtUcFO0T1x/pDV3kboSi3U7CcKMPKeLF05NH1E
SZJ2b+Ak7rianni+O0wIdDNG4YmBHQIAS9LLU25gkIHxULcj5QLPNPPSYdOdLojvINWCnsfrLCy2
Cb7inMHbmaUhCKJY5bIoPPNocBf+b4lMZJFNtQ9gq89AYuA+CgpQSaiLq12cvStXEbFl5ejGGkmn
qqkkrtG7qiXgdVusjQYcicARO0geOGxukS6dksVc1y0fa3OYeA7DUq3aguUZxlZbYMq2QkAEQri5
71FXtfACgTWw5TDLfri8R+93nYTtDqU7oHSOfZ86dFmzDMrR73rFtCzWd6FAbEB7myFj9VmHiulh
njlu0ozoUYINxXoUxx5spIl5oZ6ueAwg0S/D7b9NZO2B5nVJIG3oJ0eovUweFf21q3mHT0/yD9IX
nlvSiKjkJVFIE6qwj+0FvYli9/8iZ+VPJe1zVbF1aGyJNMui8e/slLAK7Q+2N8zWeLPtRSMLR9Ba
WyYIHzR/Yp0TOgPM59etKfNBFjnDokMb4kzTlX0os9yDSRt8VG82FuuFM1Ej9AJgaWuwjaVsU81c
gLKUsisyG9G833NEhBMqI99tXlQNSVjdR5dT5ngJmhbm4HgjFVDwqaIcmuhkTUnH/2fqd29LuIpi
nliswlT8FEiS1h9sm55gN0sfQTjKAulq+qKGXNGHx1HtYXtiwkOwocYNmd4eqTO0LlvX1wjBZ8/P
0fqu9fFUHPOEJk5wWXPXoegYzECfQ3J2NsAS7Vf0PqkBnSJwwgD5+iq1SkRiR4hCuoBVr/FGGAoa
9sIwnbHR/WISSvRFu9gwkrHbhd6g9NoonO+LBXIkCD60JvgdiBPyIk4WiFQE0rwCQ+aJeYHhbeby
jmaWHItn/Dxl32UV3bfgEqBoKY7EiIUUKDFf1Hof0+LCyXpUwjzh7dlMWFqtUeHJvV5IBbk0WlPL
5vRBXDWs+8DLF0jOLzv2qnzE4Ej6ig44nYpY68HPwZTCseW8S01zOoSGd6NfgZYOUvvccLK/xXxj
wmPXivxI1pDBUTnGzgeT+7cja6EVJfjWYG/JbrVzaucF7OHxLKH3NSUbtDcgUtKuZ95q+iw2Hwhi
0DtfJeD6Oz7B1eAErUp32q2LsrQdgCCnXxO3oy098hoW8bwrCHQvvy6KtdauXure5VFHfkSFq5L0
Blh7CgP2xrW9YHyEQzEGC3Amuj+Dmh2NPK7nA8k5HmOH9n+H7MTXVdkUQCaLJyDEfDBpbeCJWy1r
9xh3lTF4L0dYxA5s3VJrOKoMuWUNrTOjhwreFiDDtJSO8gK59ap/PzB+jCBNCR+rQL4pe0sRp29p
eIHjffgfXnePyVr4ZIw18/cAP47y1ksYnOFBjCsP4XB5+4bG0SIWCq2Aij2oeh1LXs/eeD54Hut2
mfD+F/bqIukTHCixOKUmFS6E+6Se3pDkXtNLgKqlGnqPxiyDkVNXibFVGWV/nVlB2yT77h9RViDA
iGg0SNbcMtR5qKoVPWf3O8NG2gfyvqUtBIglh47peCgAlcwtC/Fp9JHNL6okO7ashyuguwYJPXte
TrYI8ODOzRv9hf2zOsUrERiUDK1If3CO5eIYI+FSpSr9zzmiNSV9GG/wyJTsB7DtK0YUMSwPu3yW
CvxY/dI8JvgYcAT2q3P3CJ7pIO8MgIxpfZGVRf1pBVsdC/wjrn7B0u3Vu7RCQbUnhHE792JwSQ3p
OM6Tymz4Ob8sl6Gy9afJnZYP4VKYsvx6gTOpz+OuCOz4/2nsIAD/gK4mPA6GzfiBUaCQbpyCAJGX
EHeA8onYyj5NLBHWNaN2111sNeNi/u9o9thOuHcR3puz6ySeu/P6H275keaWGYLOCP8OKQHFUdT3
z4zntzLNeIzZ0Ny1ONFv1b8tn9UpP8w2JyBMImM8D64nGAKiK/jXVLDwzjSiAQPpgZvsy5BP1Mc4
p+EsFyYI4j+hChUpxpJQ2Ngo9dHJtT50CMIjo2k1Mi0tKD1cl8HknFr6SJ1dWTv6/AV+CrXsIi0K
BXrE6gR3YCaXPPaY3Nrc2R27oSuB1s/YG0ulVO/o77/VRyk++jjvQqhGNJ18HJfK5Us65EMzxAqJ
qBrOImL3haaqdw39sdMrxXyngEHIUyZ7iAulGZ385cG2VC88oLD1Pss8y9+nEDn2oyyN9Z94W2NT
JMFQSG0CenYuH35qfUNeUKDcGdT037w7xgbzrAQD0iKOdGw9hsS0+2P3PUsiqjtQPIZp2z+fHhFq
dALdMfc80Q2Vb65q5ik3PcdDhas8NladkhNJIY6/kaw8x01uEdlaUF+l31NnQhPty2YptHuLr9rL
2k+Do98or49Y9qwq7mJDTKxqbMHUnRlczO62bvqmyS+kKGEXX06ePWaKpg8r/XfK65VKxgiFNaHj
l2af7E4HpY3CH5cfJ1+fFq2wwlJse/GwO7vWTn/xd30tAVX44S96MPvoB3C2d2zB1Fl6EOZ94Slq
4HlxeZh45tp01kvMdXc3x+5fvJUcka+jDci58F5croJUw0zGVqCDHTfAQAGwUH2BE2LrvHPWxJ5l
CnoNh+6DvqAEtdiDTba43uiDhpSGbF8/t2v27kEQRTNUuKs8C3NNVYzQ/lT7AxXUFgrlhOF1vD9b
+SWtYCxKbUMQ3lyDAFubzm1SRdw5eg1mcenlAnxKsZJ1gRtp/kjdghe9Nc4si8tNN3GHO0s9+QNh
fUYbcVE9QvLspzfy0hVsefjjSpY31H5EDMMZP0MMxrQKEMBpfObznSYSUYwAdYFyHnaKzG5VDvCL
g72c2lcNP+QhBdQtAAxPgyrerA4rc1RhOmMsTB0M7P7MuHKkdc/VrxpMTFWGhdwhVHOlk5Abt6YI
59eo/+JSTK2k0Lj3//YVxXw8wIJpkudqDn9HGseKhz1+FxQny0NdibujLYpXOZ0vJR/ipq2To7dV
hrrNNYeayA4ZHSu2wjjV9ZSzw2xUIfIhZhbWTYqX04DtqjEpOY44QPbxAg37YMbRWzHp5hCPAamB
OFDY0G2lxFbt2jzQVYjfCAEYc7ZdmyFeEs16hYggqft97pX8SWWfz19zKXLcFkFuptfY7RkMP87F
eciWCwpvoBHlZfXmHdG4a2qNsDf+ha6QI5kjnqHFYb78dbEAahQ2FoNdDurbrM87hNGDSyhhtWL9
DlV+8Z56Val5lMapf1Yu1whYJUCyhI3fjbQPv6rcAFsGZUeG2FkQToLmjMtOAeMFXwNEMNpIZ+4E
eDH36Z8iCobpmyskBEd/am/gCNys5h12Tu4ngZSUDOKiqar7PR6YMF75AoTqqmXfh1CokJr9KRyX
AUlEy0TgGN84FioeTyR4QHlE3ZXtPzBTg84J01wtlz2DIX6ija47jiJDc3SW7ui3XmcHFkD487kl
yBo2XoMJOdbXpWR+XNEx73ecEzWaAV2Zuf8hlEWvbLiKhO6yWD5LRxhbjhIouoWoljHO2NGSNm2Y
wU0qq5dKIXIdTZVV/d5WgE8oiGJ//d7dXbZ7jldQHLg9SgKM2nFNCjff10O6/RZYFOdtoTQ9Lf30
JWsThxi//CEO+nL16Q0m83if3Gr5GSokYKAYqPVFpAKs+WTxse3azFotMxAaOT1wyDhp+hSsBy1N
N62vVQw+nfaVP2M07M7I071R4tWsg//bdLZgt910ocwLaEqiAOTEWuuv46CIKfcJmFZ+xTyuSWox
vq2rZpxO+7lnD1BSNoyxG9j+o8Vj4CMUivggzrG/Nv8gHgHwq4w1Nm+m9MUunAJgPpuqUNlO16/P
zAF7mVBycPamNNkRtXLyWa7jR5YumFdPJ4ZTCjJwaU4hOKLTWSfSZ2cnDlUWdOzsilGvbYb0fzf7
u21ah+sMuJcCXUcKSSg2HGI89CRPMipxWby8uA/o0Z9mL6TLIyUbaTKcyHZZEHTvRoyl6mVr8Oi+
JSbTe35cSma7cPAvXW+QXEeC2A313s/E09SqyQsnXttMqmYMiR4mJhAdopOd4XQ9H4tHwZTio26Y
wgskzXGSYAeSmPQbOFsEmfN1wUrsqEuGs+Bu+rYs/i/dMwiO8BOtOLLKSPBjfZNG7Yb/V4Y3bF6s
aZQHEDsZkeKMk9FHg3g9x3Zx+y6XWgngD+8P5GY5tuQzQww9SyeEM3wBnw9MgRs7nsMBYPlrBqvG
knXMA+TDFJOy5/y+MNQTwKH60Cki5EDJ4QXkcStOhWefYQMYowtkfKO6L4yuzupGhGGVRuYdEfGo
N9BAl/OMhiV1Y5i5uIVqfMIzYt9ByUAWDbVAYMI+yaxeR6Eqlku9ydDadchxFcxpixqVF4fTtJwq
WQm+UfYjYzBdrwaHlSW3IVcvP8DaxGSTYKqdt+vcvFHfNqXjFJE/JGfFe0OyhIAXjUhTja05J9LP
Y2twvN8Tp5VUmClVNFBcRE1hNTjvoDeB0UOkSVOf/h1qqxFlOzGBeWAgPD8XaStsfOnRFggudEJl
vbYGUvQ1V2CPaWUcXvgddnuIkRITV/GYS5R9hZA0RbkQ1O148lCKK5NQfYqOqyj3IL4PPBdI0YXu
mKtFTSk63wHkZxcvVBxjJdrN6oBGTULRZ+ln8efKbSTC05d4I8T47mFeAKBU88OnMLzfqlO+vET1
VTeV0U4PlDwR49tsUojQ7pnpph48gYk24MRqr1P4Y4Kbrb6oLMIw/LULhCSPThor5SnRemOUL469
ocXARJKvRMnGxXSHiLGFxFRukCQmUK0/2jTgXfhnH+FLQu6l5AhbkFcq/GNzh+CVUcwpbnCd4umE
7LDXE09WdN8anP2Dvb3OQ96ghei0O1oulXfFy1cpYU76S6xYc0b5LlIqKDba++6sx7FSq3oBmW2y
zP47yGR+iVYXyV/R0XDtOxnXX4lkzFTKtwy5CkI8fo5eaNaX2TkAbgCl02Sw8Tao8zTxkfzApKy0
Gf5slN0gTYhnfkXuz6CCCR8P29FRf7i1ftsaua2690eUypw+tCIUx8i0dwz5+cmaT5oGPRh4nFIF
kkFoXNtpzoBBieVhaSAQY10rgYwsHgKoFkDy/gv2bdHnVKNGGGVFSUI1/d9GzZKIHH9hWsUE0RKv
7cBdTa7AW+9THi9Dh+EReoYo6TjCrqpw280nEDAf6WqAqReAqBGEdTLu5jNpxsRB5O8FNakk6Efn
4NNPydlKS/2SYXBiCmMYyd/mJFhx0lhKLvK+Oyt8uzT4z5KGrZNqEmZP5ucoyEHRX+Juk76sKf27
8EHxmc687bxLPV2iB2L5ojRD55wp6DVzIQMiH9D7EXUK5mqdMFkGLJs7QQaASk9xmFpJKl8yskrQ
IjpXUQYcQ5UIUnR0ZojGu7DzXbcRXGW+9uyxdeWKWWerDMxp4LN8m7QLhSm1tyw/2CNVXo41qNl3
+7nfpJqzdnKQpq2xTgx+56nEJ2iANoJzkDotmqwhZO3WpJ04dRN67gIU7nqkENWeh8SyAsEnFxjo
/Iiw1CADrkJrzb5TVey3UUiM4L1/t/GsqHRdTM/OKV9FhqWGlpQkDoFhDNWO4RCvBOvRcUt9HYpC
6whJPqes5B/GuK6a6keaENX6tZ952gzhT2WcbCMhKfwujlwuMRFQD9yNw1GZ3c8FvAb9UmZgjaYB
KHMJdeMuKt40RBzuvPyAxZZL387xo2yCzzA8j0Z5j59VaGAOzbhtBeXamZkQcchdd9lERPu1Yhkh
2uJbHGrVB0IAk8BhQnk2ZFa1mVhrpVkgN1WV8045a9JEp/r2WdYtJpINe0stZVY59/6U6YVErVIX
EkBwfmh/XfMYlqIzozIHOupFG+9w+aZ6c5WsrD9xjFQwsV6GFBBjQTA5ekaT8cSeNz2oGq+ykQBh
9JRekpWvaMGUMB1Izak2njeP2fG11zmfWav6cXSk/mh2fvU0MHrJ1umaoSyd4arJ8GdMdPh3KudM
Dko0w9bMlFiLOOHVgYmElLK8GwvjcxXwrNPxeLHsKTeXWfECit0mvtO32AwEcqADfKyzTDp7xXMh
jVVDlVnzancK1IQsBj8FAdQK7Y8QknUXZGNHF2AZhh4GAXkaqc8zJ41qS7YaGS4ttkj+mZ+lZHMM
uxGQEPtx9tG8d6+ylw5Dj6C10Y2E+rNm23FrabcaeDFi2aAf2JGBC4/WF+CzWq+m69/EZ7cg/xwP
pPgOADTm4B6bMHy+/mG/9DMiNW1NPExvx0dS9CjPk+5E8G/K1BkWgtWXGkoUv8z9SYmnhUVDKlOr
niYVL9keeu8Zl7wJedweJC7M6K4ZWtXblk0T1WIfJ2/hETVshwbPaYGzuIyvNCe+5lefo8CDjT84
qTrkeOH7O96icd3Cn+YsCXQggE15pZCvTPhAWpErAujc5zJiux/IpVDy/ZI1Or2gBQYdA5Ha3np4
mTQbJGj/RuAAOOrg6mxUK8KrrLp+GBbKvbotAQRzvdDRJahfl8wGpBeEu+QFz/Qh2V7VPTjWuJf+
6CDTdnp1Pwg+IZSn2UMMNg/KseqZdhJTu5jXTEw7JZQzGRmek6RQesVBseaPosSFLxr5+Q23L00o
LhxmqsMYmLSUKtUmc5/vlaTsKbFMB48oTLckzNtnxWbyUu20LpGOL1hbSFZH07q10jArVLf60/Tx
9OEpLyyBrwRCkt9toySBpVpKgvTCs2SF+ytgaWXfTf/9GWuVEhKgAzoCi41/04wNjiAnbBr+c1dq
MtrYAx2l6oOhti5/KOj9IPb0r0IkLm2WYxs1HeGyuC+iBng6L9XjkYlgxQdEoeg/H5ZxqBEaci+T
ssTzvz8i6TVtvv7YADBhSA3gF7dzvBXEzxNw8DvvkQbWsNKVzLpwoj+gy26eiUHLLy8sW1exeBhY
zPszErED+x01ankcxykWWLneCni05erTF9nHKET+23D6TWwlu2SgRAVmQvPogJAWfQcOH0xiH9tE
98ZPSl2sacYQuS0fCCaq4HH6zy0VM9uucnl1V+GRJiWaeHuxF4x5ewvEnXW6t9dfMnjN5RTwB7+I
oYcET33ZlCBPI1iHTiwAnlUEc4x7VdFqH3G4S3ptsIM4XVEf9VqvAXutl5lp8+9+lKtO3nUddWpe
2YsaAUhXTzLfmBnnYIbujXMWYBzhTTRPNoJ52MKJQEcpoLdNZQF8FUx6i9zyTK811ppIPGRhSimV
7Z8ssaqf//G+iG0kMSQu0MYfTypVCooXvut6jSRvomJpWwRTHps5njRaWoFfegYAfjt6W/HoLz4h
+lmmySJi8zAX8MVvlTNTthV0oyfJ7thRV0lHh4q6MDUm4//53FuFR7ehOp6PITW675s+0KF9YcWR
rlYvQdDFTptk70nUgt+QgUvNmVWMYU0PUtrEKsEqFmfPHYUXcGDhMue+/Y5jgTAxxstv3YMpact1
FYe+5hzv9IdFNVIqnDH01zNe++umvIOgl0Qlxl0iA9Q8bgFSe36CXadHrsHRqYqTXtfT6O7+phGL
Ph8UO02R8pGULIvsogeq8KMOM8AUghS/v7u9g0i3MQnxpQCp8h7Akjw+NV807jr1Uf568gGdIxLu
0+zvsKDhKZdaqAUkq9jARVhDFq7qnxL2l4Cmnze+wMNccTDQa2aUFdYacW3DGjQ5aERuhoStaQet
UJcuU2QTqxT5nRSxj54rWD6/proDyRajjb8IeLTiI8XnBlytDnJtlsEJOa3l/POCWiWy8d3qW1tR
tFqKxvF5J5bmqpO2TExrsf5bxJgpth8hZGEdIdxOA9dzjoyhaK8GCMwXCbt3LB+F2d44/TisUciM
u/zeJ/bfUbvS3X0WMYOPUDoERhIzBX/CmvbVMVnkcICncRkPf2C8vsNlZfK+j8FO9ZSoQ8vOYuaV
BQG1y4QEs3AtEjw6g7gj3OzLshCqq2U7xH1kWug22RrLBB3yJCneZ3PYfoCl8X7ADZyvzZ7upK91
OmzAE192iv5aB508gmni4tpd7sXAE50R6WrMNi3b3TFaT+d2qokbWkJ6QQx4o6JIbRlnspZq6SHs
GXxARjwXloKhWDEzeYbyVeg0+UqrPo0TbaBcA0YpCMPpyMOVfKjNa3NPJRfyFekJGjvgEiAvsyLJ
VXvKcRXLp3hnUMIlKQ5vzCjI9sWID89wLLu+UWU8+5rgvz2GyKJHITbsKXqpypQbnF3KzzFHmJXZ
yuuhSaJ9W4zly9adoqmn27NKfEFp6L+0O+rSIwRitDg7VEqxHZJhxRDFAAFUayhaqVd/nyDhUCVn
NLVI3Utln7D7O5yWaqT4lnfci/VTYz6Ge0g55yQCPlUGuBsjxwxl+FIhwZ+WSCblLiJ9FssGscPy
K3gTwPBpt28MeWbwvZNDJlhq8Y7w7bbtES/DuWz8UpPe1T2H4dEOs8a4/5sLmtbMJdSDAyob8StP
J2kVO4/EjINvsOHG7ivNfmp0XVZuMyTGaA8LRM1wCepLff4SGVyxlrqJ0M71uxxANRMSF+0Hv85k
njpYkS+eWU+f8nX4f09k2lsA4ZUqVVztsNaehXzdH11ce59SCumhc+wgw7RgvmzmEqgjzwA+M8LQ
wEsawgUhJfEcDscybIBwYLilhfm4um4VKC5gRZKPqLTIdrmOFrD5kJA5nzi3Rz32rs8qR4aVVsiB
qp2KqwXl3lPucR7SU6eTzmK59Fi8GiM2GISWshqUiAIDNRWDYR5cCMo2oGlXrZ0a5ziUiqwOjOq/
D2UsB0gxx3wSODZco8uSlqelCUscAjjb7D0HShpLSoXNwUUEqJvG5LKO1Z97PQ9qRI6UMlk7URyK
EBgR5zV5gNT+J/0nU4FhAr/N/Xx0w45Vx8nSMDo8WIH9AkZPCMJmDqNOLhA1V7eutcMpE/EbgaI0
GR7oIk8NqPnSahetmTdamBnCuSEq43noNXEnrDk4i06NKpkSGtvyE1tKctGUh0N9Xy8BD4nWF0eD
IBGRBla/wn6ebY8uBYIPRvhGqPOWJKj3g/8fI6b6VwedvhsMkF/CBa/X5/DZWbyHxKblATHAdwqW
9e2epODY/OMJgdta2+TN5s7Ecdu8e7AAn1N/TDvEjBHNLJiZbCN3PdDXBKaG3vXy4NetZ0tdTk5C
gTVaH/xKSHN/2f25q7CqxgV/NHeYgRHBQkVw9/oJlkQLzhij6RVTiBM6kxfFMC1RXM6ELUTrQnko
5SmlfyYQ15HK+mUFbr4IUkiXCycMYTJolBVPg8tqQLnn/6sQFGlRZPrzul1jpSNYnGVSpesGQbfM
Z74m3e8UHZbqWZaLDje3JmP2JXbdxq69GEvQ//ehAPqn64JJ80m5dUE3bD4T4kS/Pn6KVMuJc5+M
VCUTfq5yhGMZ6fFqgAYpRM0etpeA4fEGuGVJsMnyZX3r+ahUCX9m7NaotRTRkcbdCZUV8cj6ERfc
DfT9su/9qXpaKerl7VSEWTn47Qp+2D2mxAT+cyKVtdZDHrAxrZftqxImTDBkYZSKK1van/Nr0pnK
4j0KXFC5L1dYvIXAccAn1JaewiIH2iSwnXiJijPaSwKE9E+g7sZpb1LGO6jLbKpzldhlsJkGhdYG
Ehh1ZxsUL66ae24iBp3HQdmdgRYKhLi4aq+qM/R2EYuFZi8yqIuNcL345naEfZGOxpNUrjhUgWrI
fc5TEt+lQw2cJ1l93RNEeDPITVP1kJoIoPAXH1PYhtwOoRGlg4VIx/UVg8UbFL/UweLGMbQWATul
XIDPcp8MJwTHpwXuMHo4NrGqvLAQ5C9uVT9zmNkMO/CjaNyJ6XkZvW8+8SaYeNea/xOnfEFRdquF
xSwqbWBgpwNN40KCyeYGE/5coWNEfLd8xk51W0bJ7X9EM7EG++fVILBBrfaHO2HT+YytJpXBQT1x
5ERKBOzvPVreLFSKCfk1lMb06G8+i2UOXPhwaHPhqiI8BrrcSAVlvyNz3NWpLkgiEGt4Mt90uKly
AAY3KNOMe8/r0/WdfNjrXB3EttxHpR/9+8NJQvORSufykWbN9VhA5PVKjB88uytQ51l76ChotvLq
VBHiScXe9KDjRJ1CqQR/4QsI82EyyfF+wD15AKRkVDGtBzNcQrjaEBq0DJWLfQ76lGq9gU6433+2
C99rYAG/SyOsObsbaCMTKF2BBBvrwCPigv2pR109z+L/9swFv60zwscY2uWKvq9HfKroko+/UMrF
JhNJKy1N4Z94zGxMzY2DTQp/hrVFeAQeSxAYjbAmUkfKfjlUgP1N6Lf7E7cfB2J9C0W8bzP6WiVq
3Yk4aKPYcJ2zkelmuZBlni44a+afrmF4zrg3hMv0sYmXRhdtxiul5ESzUulsYFlKwxXLaxSOoE5B
vZxT52vIGOWHMDmBLexDfkVOjgVcpuSU6eoSZ/kw+5KVP5/pgKuCCJ0X5h8OHVQm265LG+L0oADN
VnUIlxAkIonGPHb3AJvSL//HVmoA5W1UX4gHIQxFNa9wWUAWhy6CxWvT15djQGQOWsgv2dw9Vwx5
/+jro42cVjWhi6UclDPlaWTbUPh7SVS9ackPAs52TqcHjeOmlyO2WwcYXH8tGnbI8ExxxPNsop7Y
hbqc8MYdNQLkdeeQFTO6iz82nQNfqa3SntTlVdGVow9U8Mv+aYPz2nmUXMciQnMbtmXb6k5F5Ygu
c4D38jKnbnJY9YMFaa4oqjrqWqgbx+lbuezyqFZu9ttGDdPfmJ1Jkq8Kj2gFxjh2FgLTDZZB66+W
hyPIPwMbjCEqFmp9UTXWqqEHJ0pfg27TmGZtJ4ctXjXU96PCNAAVvq9P+Nve7nSLBRKJNFRXOJyN
mVTBPtBB75cWFmTWNQYGj3qzUFHzk+ptoZdW+Q0Vtf8ZGIigF99DdgzzXsOcp433HbdMaD1B5Xnd
ClimhwJy2B0pcKQ8dYdf64ZleBS8QYAO7s+fpHEO0/NHVWE3wbPfrfsrErcnM/eSrjwGrxRnG3yP
VHv2frQekOgvqU7EkCgcou4dRtB7Z4tzYchwWvb3UHSn5jxXDjO8cNuOyOpCDwH73t71OjdxuOJq
JiSnbqvizdAE5jVqRCa1BZWNqqwr7yyVkFw7jtm2jzJm1foQp9BLRTIgTUxd3gXIIv9O0dmnXL7p
qd6Om3ngAjHo3/N3JsXx5MF8X/4zzGMxMqnhQ8sIIjM2ambV7Fve0QMOv8imcnj3m846NVVNs4qT
Pnti3x5gsYuqNBWBVsNDXNKBZug7TWcBlM08uCG5XmBypdHclaE67k9Cp1xZmwtGqzlL+a7fJbkV
6g8WeVsXUKuvDozQ4IESNVMXlNkRpGsDOVuJVzpd8LOdB5gOruF3frmI2Zj7CeWHKDgL0qsGFMzi
vI0w6o0GmhcmEr9MMivCw7OIHeXz3kKf4Ar7edWJZ5L+JZ/ewmr+odNUpgxFebzGowCgt3A/jrx5
Zbq6vX+x8orDF0fEn405qV/jI7gWgz4x4BRf4WOw7jUdmux5y/DrV2RCJ/LL7KX8o5G6HmZa0BTM
Nhwk1/zJ1BFqaBkLmU2l0fZPtFuqB1n2ukYyPZF+65ZABmsLAeQgK/Eb4XXgJGycCTOP8KDvtQPi
uH0LAois275pw0eFe51ZKpkYGHOr+k9Gsr3MAD+k69pLzNAJGwKAi8glQrfRrQr5NoUxpvzpv51F
KdY1RuyFvDUzB/HU0up96T+JnICURh5xaRf+RQnfIN7VMSZkLKnnJqQ3HHCHDdEwsY3iRe74MOYz
KAeXgahtckmcV6dxI/GrmZQkpDHdkFEtaImfnOTp9pQsy9D6NPsFro8Jc6JJGEdUH0o3FoQt9H8E
BcHFlKOWivolQpraTrLdv6t9evboRFS4Lhj126UWThYE6GNvknMf6eyNI8m9rljxoA5OPJnKqb3a
wLJeT9/rIU/xgMC/BhRxAvfoGx/MANd2LiEbl33TKy7r7aYNY51B51IVNZwIFsCaSJdxUDpRDonn
NBOyrFKK3nrdf+k443tjPu59jSREwXiu1viVUmZkZM+6rH8NWQF4VoJ282pZjjVRvWe160WSHkZO
gNdJMhx5sMVGTMX46oEzolYvvB644Av2Dkqo0gB2Tc1e9o0uc/NNAY/epbbyEMDvDdGkg/MdBfrX
mna2ID7ORRIL9ALAfINrgsqFuVACYcqshrSQuHCImNBGahHqv9/nqq1oKI+XWbbgj0+3kr1m4223
O9ghy4v01Xn/fZ3lgdPKLUvPCmchpXnAkMxRDwCBhvyOThLsXdTaymOJSHcW+xBtNhi/lmf36OLo
btfzM1K+cTWMtw8EpOIqr9rGOmgYoCD5M/HK9bjZJ/L6xa8zn9fHVAlIcmJV68qjFzJX8m9wvcZa
uTC27yeJpSE+nx5l30XaQ4TsiRphRyAmHGEwcd6gkeAT+DFnV8vUzcPCUgoiaqZeFzLvujxHF0ga
V33HQwjF/l2rb07Cb8mw100eFrLRBEIW6fBF2nCTV9Swqg1NKREcn5l/TjygcHAdKg6Vy+flNXsP
E+J3j3F4B9RXoIJAczyrZT66hbwnIcx84HtuO+d3kPU6Glbu9EYkBF+0tCFBONSqMetwl5klDvqi
WBfofjmPLK8KXqkN7utGyUmvFcMSTIMDIAt1PlZC/7E0p101wGQCfhXqdbWisL/M24AiKoGfpv6h
KuoUrKeakT6pebpjDh2Nr1pgs+QVGhWeLbt0X/YGLqc/CBAab+Gt3rZViiQnJ+CsTxZRer6NXJ1/
yoh5+yYc8gXvbYjET5evBAyHbPTLTZcKMUGkeGlOV2xZN6WkbJTnG9BWOVWgshgqLh63ZW7Ykk6E
4F7LdY7+ibl3faJ33ztGakLDdHckNjxGOkMU0wv+U/R1fx2Ju+wiCJ5MELqcoL7dkdHoxl1OemV6
CsqEKJo5Q3oi4lE6NDRzVslIG+VuMNG9ZLTYOdX57t3oCkYlAqOhyIz3nCbFrUOGjKO7/FEU9W1Y
15idUN/XEB0A0dFzWag365kAww1Od2DTrQadzhiAX2tkyWsVL61TNZ8UG0691X0ED5VuhI6BmqtI
8DRxpl7bWLZi4k/jiBveGqD6GdrZEsMWQMaj444+lsgWcgRqkUlnKa2OXLCsa+PrKrl8O3nnAr5C
N3oAuIbZQIw2NgE2Ufkp0nWJj2LeLzQQwr7lej0Wwwe3MOodQFgULaCjqYpDCY6cJEBL3TTnJvhi
6zEA6CsALQYXXw7xhTYl4IYoZyBZlbLu5zH4qkrFd2GwkEQbjJl5sGdsETVZ0bIzHkczSzOrrR05
srQpMzaz99EwA3PL47uX40DuJ8ouEoj2yeCh3zHSDructI8aLg10xJA3HqiD9Bg0CzVzeUBw152D
hmy9OqKuj0yAd5pVxR1bIPlrPS5g2y61HU5HY7xASeUTfJ5u/6/qy8mHIRBR1lJ+Z4M3Sh0OqGbl
mexTZSeXUd+pIhSGbsbTrLQqjUPGbHJcjj8j+pwVZL2iG3WB3kptvFxVDUwqgE04zkXelYJ0NVkg
+BBM4w4wfOf9xVXcW7fEijSTrUsOSt117yoERthvHsjLr1xtvpbaaHiDph/TrHBolfG6lrq8KQZk
eAmDpIq4wQOLQqQi/AqKrjanx4SZ55Szzi1iDQIuwXb8qgovy2edCobamyyvQpsLMfy7YPw+kn5c
JwiTr0qhPSisGRemQYI7fm6VfNjd3ZJqJTUYQJfA1fcAOcx62Kc2UqIr1aNElLd+pUmE72wI4FcK
+uWdxSNwe7gINQGWPog63ftzzJPYnMFug6n7rdq946+ALNfQOzhSlV9b7f7Xl7Nfj42fsz0s0Mib
anom2ysHCUDexbaKfWot46jhHQ0X8y/cWa49a1Qbpa80R0vio9af8Jk9FpaTbepMLJ6e/vDhTGjt
oe8/eVbGFzpq+AojQr63CAmnNd/0BqC9Y5RtrsCOjIgXdi8e+jemTsCFfCTxNKVEe5wvSgHYIv0R
4eV5GV9x+XxsCDgbwZ+ZxMaZdKafNGCOtbLWrd4bh52qvszw+sQkYijh/16i3OmRNGM1arZ0Nc2M
HP1Xk8G313kksQ3eMoafYGilsHd+7MrA+DNkBYnFTxD2biTAilHHBWbN2+NcVaOaAIoxO/E3nt99
WZCqPshmPIp9GwBa7rfAcQUx21grUPJCA9p0jHiS+hUW2rBwhPAKWlvZAG3BtGPbS1mj+MRLO9FS
hfAokEFIaeNfAmpYO/7vNQahJADBPEiA7UsZFQiR/qxqI87QOB5F8Jm6YjQ7Szx0yYw2Gf5aBHFl
YLnBMNx1TC4lxXPP1t1K1DfkbLjhJVpfs9dDDgObR9DLwjGSZhp2OGz26yAWgJd0GPvg/qnLGQHr
J9Ryjiwq8JJQUkn7pNzuWJP8HJx+NKXeMsK8ZYqm2nPWqZ1BkfTM9jm58+rQFC8TYxgAr5Duymdh
5MDIoBRAPTUVTiggQ76twikNN+XlfyNjp5GdFdit+taknrU4Kh3aeFBiAuQHooK7AthkNRlYc8e5
0sZz41Vr0CySvFf0s/cscljUF9BmmFxs5YXJL288iQWZb45FYHr7Q3mafxeP9kuAnjvE5YbMXg+M
YJ3v3Taa8gydQaGk62RT0OYibEAvguzVexCdYBpV9aWjX/k/xIkBsGoEUzVb6NNjPeSHvnMiOlv9
k5oKybZpBS19rMOWE7MQ/o7SO1ZlG9Z2siSXSmNV7dye2jz1wAV9U9Wht0+EKbPmWttO0ctoGQja
bGQ5HqS+nN29K+9BOdSUdslWObJYW16XEPFOl7L0gqDKzuodYFnlvW3DgKaydqjJqGbtPv+ohA5n
NYEgSY58y6TAOlP2niYe7sPrWLzp1qH2F0NOIEZ++/Mg0e3LeO9+jRmwn1OBh8fIcQJP1yScPo39
BRrn9fBRCBJNwp9uwQJMCDXLIAbnJXZ2afB4q923rxduT5WoOYHwZFx7fR45bzy74AJlh9BySZGd
yN3qYRolwkGzaMtsuvnKF2BaDhC9YASdxaZHyTGlmARgyk5KCM/98mXtjdzc2B9Esu5Ab3oMOtri
WWN1f16q15EMdxhGyyMswVen8r88RcC9eRZVzeSrdiDCYUbB6SoWq5lOVVxp4XxidVTV4+iVuKPu
SlLrd9KfsagwwFAfnLEm+Y9148LPH7HeVMAxIHzwXz8SxIgeffuLgmB/8kkSQ3Xn//OjpfowLP6c
wND1JT4BIRmbeRO4LAIaIT4wKGQysPm4BAEfG/Pjm9mUu0W0MuWxD/B2EV6AfIMreeIce7hs+Uq4
yXBd4IG0YINsDYTZztMeOrki9YFM+S9vI7zdlGSwPAvt9jsoOzyYNK3zQyv3M9P+dF2/M4wHsl6a
JG+6YRp1Cumg7rM2lRkxLursHbvKOsUijTR3bkHQ0A9bKuJl3AzgDwyhdEmh+Kopy3BqVEZBxwSZ
kSCxYCm9UZflcb95Vz2upvN8m7CDTOxr6gw3Lz7vSSfGZpeMpJJAoB2qK/wqN1IDjAcg/m66f1nQ
BesvD7sqPk0NDpXDDBJnLHNcAMmpidrWlXlDxvURFepgdO3+389nbM7n8cCSC/POjdH3u9ZvrlpU
jzA7fhk1wimYqChLYmQMi5NsVP5wo+BFlO2YnuA6tTACh1wsoStJyNJNotNf+1u0JXQGDYQngx2T
ebXWdQJ8SYQ1egb4EF8q9A3A32tDgCPOP6WMhpJwG4ZZj9pLSdqCaX5ozDZeyH5bZYMLhfJubPGy
z0HBSq11Lxaug2JnUeRPaqBYHC4us0WoN5FS3vmcFlUXkFz+7Jit2CX0xUKPElfLOUMsYt4WZOt2
j8tZvKzDq+5ky88w+cenf3fuasYOVf3pFU5nKCNzv/k6f3NchLyRStJlddcmHtfEVv5cN21nfArB
NM7UakBCcK9eJYZgu61Uv+WzCBFtl5LjLhRkW5WkaF50pb+Mfhg94F6+Pbk0R7VRJglEFs4+7L7L
IpEaUIAL+H67KuasRZMWGJNHSWDLolPO6AVPTzCPwwtGxezEWGDeKjDvuvKWmPh83THmoTrlmDlx
6VzSE24LYT5igwWtRwaA4znvVR+uhCn+N6CFoDdglMuZspy0WW4gMYSqpID9c9ivq+KCImUa9hIn
BTHoXSQaG5rJ8GuGaPCyTmRZ0THVKIXsMA/W4prSqBxYHrChJ4+Pp9x09Goml0AL/POer3iZRWjv
rZCUDeV2ZbGiHQ2415C2D50Pba5tD0IW+rR8szWUqRQKQy2cTrY9U4Tz/1xsudPQZfXjC4MKg85z
Rz4hZloYgT6JkwfRSLCU2++bTFZ1InaKkNkURHKxJ3HiA9e7WERdVKQOb+Eqlt0Iq+69W6VLaspc
TfSRDf9LiwTcyDD6XQ0IDDwJZmGptZ5tZZ3Hip22yeal+42v7XdCgPn7dB966zLrunQmiHuuvlRz
9pFtgnQzgOljowCTcoz3Mp/qIZg8IlZ3V1WKEZAlqLPsEa+QIzBTi4PBXTz8AD3W2uRE7xctfbz1
sN0wgn97LtPh1YW51TMxe4oCdPofsBPmeu8lbqG+wEuAxKSJ1f6vz5KuaFIayYp+5RhTOd7/889Y
0E/1tgHJrzzghh2QoidJoO2iXaBsutCYk2bg0SlgC02LaG1D6FApI77wPzfISAid5K7cPhP/Z60+
h2QbTHYRs/nxdJCtbZ5fMZImdYVQ/T9yBFUp64kjZdEVa/KgCqslsfDzRjkYfhdabve2XxUAMeDm
qjDLfYc/16jKC/Pitqiqcj1y+bahPhTjIf2AvmYsUrgHaUsArxEZaeCzKMwpn/rbxevxQSv8jV7r
l5j7CUQUSBcnMzTmwigUL5dTpP6JLopzrZHLNiOYezST7doQvs+LqK422HVuuPbTyiXfQj2/QQ9B
O3linM16kgR7ULKhA5wiwSQV9P7RBboxdwKYJokdRHGqfIBHeaLgFZuozjFvJSw0Ty6KQVDsWwHg
ULbYgqCb+c0wRdojtya1elzCyZfzU6JeFRbgbTiGpOKvWu/w2bCU0gIBf27/wIWKtap+tT8QEgqU
X0KioGGQdt89qNEl2nssCeuJVl4Ky/njBzGdZuMr/Ls/InsJlb7pFiUlv/LUWNa70UjghtNuG8T2
SZ068MvqmeyKGQTsbKpHcW7ar726653wNWZb6Rlziux6+cLZwXQ5hoWugWDF0E5hWHm2E2mUTxIp
Wuds+ZVsS4MOoZJCsMS9Lrq7xGoVeKWfG6hCbq82ga7VJbESdek4l44yxR+mq/MAJD1/LYCzrYir
/uOQN/5Cjeex+qCOUUpYKOSnUc+c7l3bpwr8LcLE7RJt5RCrmDDCWSooAdHafQFy4wpCaAftSBdg
BB+kila2JdRlEW+3oDS3XuO5YfKqmkBsvBSa8D67rq5cOL8OsGdwXrMTE+kbjN9K12w9jg7eVVqg
iDSsm/ZM7JlkGsrroMMZbkZmZnWVMDi9rprBMmSkvTraecYwVjCHvlmVop51p1CdeK2DJ+Z5V7Ln
V9XHTwAinvUuyXiXBInG5txzL+ODQEkWexUlv69LuiYZKXhqQJmB/Z80gGv2k6XizhVf6yyKhCTb
CT6XvO8WefrFU2H6Slf6oG0K8iAVTwSWXB5d446YYhqNc5D9n8Pb5pwxzCWaMtVwzXCWLShO3eas
wliuqLYLLooqFCAmu/I/GRBlb4gWoJe6I7WFVHbnVG70pQkV6Jdlyr5T7aU7cGBtoAW9rn3n3az0
xBp2+plkcqMEuZLPtCQaV7eCBGQjizUzvdXCpeoCwdfDHVv6QCYKpF5cgUoVBX7v8wVfocdRd61c
vmDShC0jSwVHzcTFflLt9gUNK9D4hhxi8v5klNZFnhgEYymjWFQJlDaxTgDDL+XOwNFadKa8xv4W
KZ6kdrt2mR2p5HnuWIqPeH/2ChzwGXONSNEzbNDcwpPi0eM8tZUZglRCEiI9CCCCD729ZtXzGLU7
pLuvhq6MhMn9ttFtVjfSb3JZ+x41uQopC/x/hazcTRhxIqtqAE7O2UNyfZGpc96PfKJ1azROYAOi
C2TAXmZPOT0jFQWswVGtfqg5XhhZmBqdFTuKX90GEAXsjmJLA08BgCnhwajW4xA7OBnsq7oD/RHI
YGxVKPZAAu4+jbOeZzha2sy+97SULqYM+ZKCSGLkMUDRiYwM+1D6LackbbxbmYO3X8dSLLFaPOWX
IK3XWmQnxJwvZd+aeJ4y8CPWus/th9Q3JV5vAITCvSGtuEivg2SJE53UF4D75a1xMZYTqmD1yJfR
DGH0EfJbkDLm1VwaIKTrwuQXs6zTkov2jdEgpGFe/IP57Pa2BwuYj2W2n2fyfGnjixejSUcHhkgr
Q8JpaSRlBqWrCrucIUi26EEMpGU8Qbz9dx66wEkBt2PK2mvjIXTFe9qmRPZ2F5a6hWel+mEFcH6X
YisK8Jb6UItV5H8OiQpnsy2hXuir9lsQWLhxafinOIyDtPs0Ypkgr+cftav+YSvRq8NO+07g2aNH
mDhnr6tSjpBCJDjZD/ZLRSNwPjJsaFEwKlZ6qZJAho/APoicOwRb5DcTXxbD0m3DXLr3FcP3fzr3
Gt6yxudUVcgRLT67wMZVQBx/Th3ddnLd8TVla1Gj960Bz+RHBIWeAOp/SnDedYHisO9wI0XPA2MU
RAyWobVQQaxnTCnoGQnma5Fh+8wPNp0Fr+UFD3CU+sLLlgLvoWa6rAaQHcE2J2rLkwhgJz/i1c2v
z7EcYqheNrwAZ1HCM68Kh0ZJf+HTI6G9sNpvLqE+j/7Zt5KNt/1bgwAacUiKmybyHFXzx1WvYshi
qQP4afshuAExhVD3NP2zOvxL6J0X+0iiyHQQgOK5nry/+bSqGUxSq6qO0PAESUzxSjDHBy/gVyJJ
Pr7OJhX9FMYFUTrRz+cxgr0NlQw6hGUnVlGl4c2jj+vzU8DPjZml9FnvPcdj6dDnTXw5kmu5KRbU
O7454fAbchf6/mtx51MYHwjfiDJeBbCK7mKm4+S4vB/GDBky6RISYSLNdSqP5DDHXpy1qIIJ6fWr
3cv/pGZ0/jCJi/ydYBCw97ArhWUhthV10vC+Qts3NOahFdJ6lMc3mZtBoMwZmFn38alS8BX8hA8j
I4a+ueOAMf6dkKN/hFu1yedob67HUP17L+y6oufRHgmu0EFV8Os5esXaxJFIcU2T7q0VSBQmmtPg
fpYwtG28aGQQ+eWHCvL8TIIrg1pibyGw6XCXx6mPAlm6gaqbELWA6EgZDHAB45b2P3DqJtmgxhUp
ci1VACE2qI6j0wR4l+fpP81eSDZID8h17deQvVxwuqqsSbUzlZR9ii/uoimwpChFcCTA2nY8uiFn
tMQkCsm9IL0u8i09DiFoesYEKk6TP5uvqxh6Z15nFalEhs/Znlk87wwEj7MPwCCu3Y4TcMvIPxj9
kFllJbYn20+FQeLIox3Zt99b96F+vOoRjkHUGaIELwg5NLTvX9MVURFXBPmjzoLUAhGfbIFXzT0Z
emCTvK5rjiLi3ZBQko/gmflPdUI5i60wdL6UbPsp5Tn1caUQ/8g+oQarOzbg8QYbpxX5Ttd30uzi
lax87Zojl/68sXPR/OmZlL2YOQ59M4s8nxWTPRrZmfsXoFz2Wtfq1MPYRWFSL0SLmheQ1kP3Yq5t
w0HmleDkCbv/5hxJvzB+u/hKSSxmzC7PxgO2g8nNxPqHwqPQwAAvRsOfFZWaMo0RWyQ5zKRDPbSJ
NggIiqUM4SgB3LT2yf5dSaJFTv1r2tW1+0CPLKd1TaXzA+O0/+YyTJ2Woa+RqziayYy1xQlMSKpT
uPRUmnR1prZxqRs2QbHyMfWvKRlyLC8vtkEUlfm4fUmxl7zhFV7zOo1vuFXePZBZrpkGlGVAh/oV
7KTFkhxazNxnPEYVNEcO5AKOzNjykxoYVdjcsw/TOyEDBq7w0p/+Qi7cu/iSiI/2K+Ka5SFK2okb
xW7vbJi0PaIH327H/7mKVrSeeqlKW2yghkBp/oGYogWDV70pzhuZcwM4bjcaYPW3sDwwFzTCkjPM
B7AZUAI/8zQ9geMkQ9x/744bWyaHvpFWFdhO2t5xNEiu/AD8pbTafJETyKQBfdi+oc1aG2RHC7UV
F778rAZT5bmvpv7etEJ64eNNmKfzb/fxypLYPcl+R40J0j02j68YLiOeGtGIREWcSLtcIGTL5Dc8
Ka/fEDs6akAiQGX37u7w5yE15ENXyP8ywd3xqAHoTI5fM4m5jkWbnvn5dzzMoKQq+s5boQOXZzIG
CPaMfKzXW+gFU7Gr3Uds+/GpnqgoBp9hVtwDtWjaOyIDh9iAEa4CxHPwbswvtMLiRIrk07kItiBG
3ISaJD0TiRmThHDAqS/Nf4b7CtTQ6PrAQjfwUXRSyxq+gl/tG8v8WPxFLI9BLwS0db1ghXv71BCf
G8BZwj75MjvZHskC1SOSbxCTSs4qVVLm+yqwPFFYOZB4WkcY8JSrQYo8Eabdi0n/XD673Wi3vFBL
nqx6gdhyy420EmxX8yRfCS0A+kDkLMnljO8PSRfIMBJrXiSW5rnvSYfq2N1noY97/cP13/Ov5TJW
vAQHND/f3hEQN5LtEY5Z2uDra6aCTHB0huP5iUIEZRCw2B3k6UWyKruHxAaCsB6ZM066CbPhxOSP
STohY9S4XHZn4ekxFtNRXcYMe4PN5DH33Hd2MJa9rPnDyynw6+uuLg/SFu9Ek0GKDNL23mZetr3i
zn9Iuhcd8xrVJDbBLxGYKDi82fKfqI4iiW7zcR/KHyZR/WqLWkSaSEGCKSFqloyAb/mF3yqSKiv+
wn8Sj11Bk9Shyu/jhb7UBWy6ljCzVMlwJg0iVLKORp9VqK4GAQTNV5ik7tkafYvZ3YdYKm4OOad1
944mUDvRUC/BvQPCaEnhMyy/z5t6RlM91ShZ2mImBrCH8fi4VNt/YUIvn6K/7t0JtJyrXVlbter1
gN5HhUtcDldxN7f5A68sPNheFF0pVHbAUnQcrTMOYJzqV4J+YwRTxZTSR/mOionQKxPDmwuTlr08
d7qR4vgT6txL9oJVAtEkUCQRJG0NXtEHCtXdTfvWrclGC6kkn6Mm0CVPQfH20jgTV25YSQipVzBR
Iwf/fujbQ1+At8s7yWH3Y3R9V7wFWj3Hqgzg6Pd8NOaLwIYXjyoq8d7q+llpxKV+qBXrUM9/1hJQ
Esm8eBvr5CmZnU6JXNN8LO24j4HRLK613hzLjijIDkaL5on9Pvr7t12GBRM3qeJHzvGxK3A0I6nT
Dvp8mqO/4hcuS4qRwZ20/iJy/sKjssdnlYiwcvQN6rr87YEokj178mYRzJ6q26fyH6GLX2//cXoP
/mBwplex57e/1ZlJKshBBImzjPts7DzA5ZAkkCBVdZIX+QwyXxT16leQeBiCBE7gTlkKM4VoMB04
Gz8iFgKRZok1Qs94RJA4BSoBNcAxgfDihv3cGmBkEzMlMoND/KUlwpquSQ5nZ3SB7r7i8HQIlN0i
Pn6HeAI5bIGQtMCPh4iyFRUlHUPQJ8SSNHIHhuds6YchQcAk6mHVN3j4alf2XFmTqm1OKgjVZtwH
+8cX+hhkOzK02zRyfLBsJ8Ch0R51en3ZWDCWBdrYFLZz+qUa9vk4grEAbAiDg0RfEjqkAOeGWn7F
Tw0zCybkxvMGOFdZj/Sm5DsNO7mMqjGLOT+7bALEj09VHjjHEXGo7aG3JCiO3AjpmKmri7QbKAx+
Cr2+jdKPcYu3YZ1dzIorJAyVNkxHCRHkCs2luCRyZfYpHBix2r3NkrNZkrInI3vsMIT4UC+NQbJe
sZPVXOZ6jiL2kB5MwuSS11A8eFq+NxUA6Bveyoo19IULuCcTwC97Bhc2IWTZUOQjRt8dfVciZzQ2
o4KXMEfRYLFSVI2BLKt45zlOy/Cmm6jW3w1W8rUpKGze0FSyJSc6uTMIxfzPEHuaLQESGXhBmn6Q
ok4hXtOR7lwV5QqnlimyscD32LZHmwKNX0Ztg9OWGPIL5Qg7sLZ3+Mj/t1w2WutAZqrpJss7QhpZ
0SeXkIGUjrXWJyt1rakWNopPdQ10C9Mcia66tzZbpLE+Lt4x5eRF3BTcnrzRtpQ0JVSaXu67viVS
4zob3Lg92HlRSVNp17qpuusbxya1lxI+8Y8dEGflpSEED20UQB/pKG4ZO65nyQeoY+pfCqA3cClb
ZPRPArAN7mwWl9UZY+5ZcKEgt7+/4210b4jrEB8FOx+Q4KinWB6tdlNmatNhPiq+k+tMbgN2rxoi
gYUF0cueClHysgQ9mSksRCy/7neHircTxHJfKaFr8jZ2ASfEvcUkkWflzXlWdAMZEBu6irGA/H//
0nPFMW5ENTlIaUM35H7VD2yJ7ZaooJSbFBQlbK/DfiFKtUK+IpPPKuqdo0tuuSFLoQ1QdG8nEIaF
LRXB2KritgfOUxwIMK1Jy/XTt42qJpYAnHlts3et8t/xp2D/5IOflvT4PXgW8P4bGnruCAGJv639
cVfI6k+PcTiswuFdL3O76ZNdAQ7ShqqjC++kyxNKIeDoCd98ej7sn40gpo8O/JHv63hjsF9QHzpm
7V3Dpj71dfDBk2WlWXRC9hG0bLjmX7i+ndEzkZbT/d1ykH5Lo35SPq7SgDgzKv5zNuCyELp6gmW2
9WakmFYUnOfO+WKyVxHpxwqkOiRAWyOxv+tuMdLJ4+TAyM7mg3iyci2H5hYtrngn8gR7VCHGAjNR
VmEFPWHtxpISjrBiA9JtMsPnewQM2oe+8cIQlrBWYOnufEJmMdE5VBrAWFNer8OWHLWF+4z/4jQi
NnVpNOmThg3IK7okda9/B3LzXb1+4J5G1HEwb4Tijr2YTYvsqw6yxRdaPrzLNnp3vUL2U6EkhnvW
XDuL2kj9PehljD8CTTTsOsu9TwzSV8TJgbPL58/EUaekf4lGyZLhFa7pxPaWnNwupxl5DYMHExoq
35VJAEBKrJc5ZjTJjtFBx6oRgqmm1URsUkovXYYW6wNqepvaBCIn5J5k0juWFxeqomoElDPXe+vE
rZ/kBuM9XA6NL9dTP77K3iK7ivbTQnWP3PG2xM9a0GgHhJeQ4SfHc3hDPf1jDHOkvU7wEJlwGuW8
MFu0Dkkl0RHdj64t6eglnIEpIZ0umPIPoMMCUp5KJlexugTzbcPKFQImKTnO6+a3+aFstxr+6Rqt
wXSCYbfeqZLWTML4jDV2ykMD5EIAPcolqy3n2iXUvQrqxhnlKk0EPq599Xy4nX7Yqf1LCKRKjn41
MZDduYHsebDZ0BFv18JeZQOJQDOb6+zET2YXgPobGATqoXAoIBG2RAd5A7wre789QQjXZDdlE8Qe
73vvuNv7l6cR0yUiirhj7oa1SKBjuMA88Ov9ZgMdH1Vz5rCUyv/6eyRYZgC0eFWijuav0iHYctEC
Sb9GPbKfkzY1LTYPRvr28KLzHFe7tEsYY1Mm1H+cYzQQdBv68TRWuYrER9rB3M0PbTeEVdjuo36f
DmVln/3QxiL7WIzCFSPaA9NSAm5PKNt+ptsb8Kn6SYMDu2CJ8mUY6ytx0uUWvF9M4FW5MfMDM3gf
MrVKADm681NoAthB1dzuP7adIqr7eOkIerxUqPK1h34aBKDG41fOwISudA9zPVAekOMX+SrIctqo
+V71NjWDtBZWLiyRhJdfeIWqWqxZb1OugV2KbQQU/WSz/+dH8yFhQgVxwsexFInEgnFKSv3+kOKW
+i/0VH1PUX0+t4LjAMNJmCYx/EXEcn7AsmrnAjweVRNLnAo/lcCWF+rDbwrguIYAxOD9gwuLd+eN
r/8EjAMUWPV1VXaOQX8La0n9IqyLnQYQriDNlWYoIsZgK/AymN+14hE4/ePie24McMQwi0P+kKVV
sTuQtZHbEgyb8/k6/ACexIOz8Ya+2+449Pz17ojPKj1GARHdy3JV0Eewc+oQI11fZ37Lsryem84f
qPlD1XIFZKk3rQ2lhhIVSJs7XNEAKO7viu6xlGyZRAwOGet4/GvUaef4F3mL4mXGxoDN0TTv1MVj
Xrz1RA90K5zURvwdX8Kw8lXBJVbE8EaDlFuIlX0owS1QjOSsMKshpXRNVpk2RcQkKCuNpKnl9egu
n22hM7E3+a10BQNJpkY3Rrnfc4cLjF5hnLRThtdLz90B4+dOgCX7XysL7UZJJmWoPNprOdEZzd31
tMJwxXYV4gUrzeHbDM4BHLAzjrNefWnkRc2badWTwWjKp1Y5Gop+4HJfPcVCBQyWshPOf9ao7SL4
JGdKrzWr/BMXMzZBfjNE5TGGXw7tlU6ComAfzjGtLdbXlnEHFl0EJQOVVhDYDFhOt4SZ1h5DQdrp
sAJwCjSIysdilZCqSCDThr+ItbL6VlZhAX/wVqxYwjiGv1Xqacf8/nAKZV7GlVUzXstZnbBntYyU
DCJdZFSTStgu2eVlyoXS0RPglXfNulMIWZPI/ghX/lyGvCrLY1yZ2l02s3AFcG1ry8wnwfZvYIau
AjIvKZn/jrLVGCOoVtNQYmASJcki/sOvaT7vc12xjNyZ8FobSIUnR9TbNdPYhGrdJU7ZLI74Ma7b
ClPgt4k6iiztWzfclMSbouP6uqmT7KG4tmXAXP9b8y08QuEG+CzD+WQcaap0VAeGbgHZWYV4sxEJ
c6y3hrQ6tEqkkPtjADwTljVV+mprFE8yRd7U3PJQmVf6dhiT8HKVV0hfD64DYEa6b7RZg1Gzlnht
bRrpPWLJxK1uMPNNXvzlB3GZqdx+EbB+FMcm9n4q8JF7eOjo5IAc6wlRnO6/lK8PMmZMyDCenpN2
8WxQ8DlWbVYyIOwvnp8guAmTdzDDhI2Qc/t/0vzLrjE8uC6LIRMji2eR+9weDOUUVbPaX34S1Yk4
ptunJ66KBYGl2qbDuykgp6cQ4Pntoq2ERm1V+ocTjpmnnEDvVCHuGl/Md1MrCrRGPITvw/ZV/djZ
yvNN7yDkobFoy3zpJDS7GVzgYX8JUJY08Lu1X7mzb7ocJ738ZiQmm5516XYXT8mDeeRbzqPEVQ9h
TFFQ5CeReloRWkuqUB6rGQ5anJac2U0e37bPEbtc1tulUkMaWs3SHR4y6rIMWW+ojsgeLME/04bB
0WwCiYXlMCf3Ov3AYkjHvSVqaL5NwihtVlBya3iKSoaLHVEUOAr6AM0jJ+spyKlg46nrTOLDIFgn
qbATvYsKC41auxbGQ93FnTB+jzyOePIldWdmhCmkICdS1aJJg0vveeJm8nCUJxeQz0nPlHSjRJg7
5jn0OqwXl7dsKFrLBWurSB8wAFAkoDWu8Ctx+2Br5NAP+hdBd1A7vbyNhn8ED+oEvuJzc69shwyL
PMJ+j/1TGnCYQCZmbGcTYiexZ5CQeLA2G074e3DK25igEZfIkOF9M8MYvpF3o1d97XBRxfrWcTID
8poioRCqHANxxUOnXgrngF4jdaTaBzTDNdrNd0hQU2K+2MypYjCF0mTnQ30DUiquTYmA+TUNoYmn
h06KAZHefsyWi3VOdYhtcw2UrUyRN6ywYzYBpYlVac8v3o8DyHclGNEG7VYYJL41/yvKVAn+O4/V
PHhnmFq6JPGiAnIzZcWQsrr5xAUe8i1/QmjeABscsqnLRlHPDEggI7eVHZ8h0wiXO63BCoiD5JbT
pPjsWaDfYMhXWbsUagyrAhwbBV8f7IxQhoKBmYcVka+sU8OcfNl5adOjO86imL61Yf8RMafzGcCA
0MzD5G5xCxamzgnJv2YJUyQgBBaOU0oY5z4JnsLLogTeYdvCtDRldNC6Dk9MX3N5GP7Ruuoiw69V
R54MUYu4IAgg7bwHlRHqzVHXrNh8oGgIOgfe3SeymSIuv3Wi588MvQc3Ykl5xAUyOeo3zgSgu3Qo
wmeckouLT/mIu7F2ZWM1mFl99zP3GvJ9SJpY8f4xKlKuyTEgLnu7ET8lBDI/Vh78hVLY72vX+yl+
ZKNoZ39aBmdO3JSFxftckIqnX1hqgRFvs22fRyaIgACVvp9Sw7bFDyr0CGNWh+yw1rdAA2C2L96H
Axtqb9mOqfJ+5xsKLLm5E0V49DOrvkzlj9RyjXKKHLnXWNKn8pNtuel2u/+xZviYZitE5s66O8YD
Va7wyCiZ5y01+hI0Zf0AhiEYa8R+unY589ZWgubZRoOmGk2RY9CVlKJGUT39ws+NGffbK9DC2okn
fDYXFnzLEjLcG2Zx1erdxq8W8NtYVVNlWJ5X7Gf/1pLh2upc2MAvjI+hTFz8hUsKGoNgBFXq+bdH
YoLZxLRpEGQkn5m+OaJTGPFB7NLJjjmNBNgtdCUjN+zsQjqnLNm3FUvJnwAn7ypfoL9uHmzLNpz0
92zzazmvNVNmmsFYEiFt07OrRkJQTNdUVa33CapXTrd29CJrxJNa94jKyaPlqmH5s6k+W/vy6tSd
iDENh9jtuuv18C0s2TXsHpD8fuw78ReURt3L/1ejwJ+jpXnhmPdHTHy5MAZJhIEgZmGrK5S8ELZg
FBPopCAmMvxcBqGKpcF8MDBD1LLkGUrFJ5/Uc8bq+GVAPOnwaTa483jnnRDfqzufGZ3jxIxGPEGO
nopnYI1zn298E5RQ4jBiBFf/ISoMrrkyqEE4AzD5BRDhNua+Xml9qSrtRJ3uChVdiVkmzYnh6b8L
DxIuklCuV6nNL4HNl0u9/nhL1xnZO95ShF/8h0A2+QgkXNeP0cSw6CP0z9EBxZ8LX3dpVA3i9rRG
t1sRI0nROoreeTiVXzG9jMUL7DJNTL/DmEb1PnTSCDlbksNI6poeLRinmoj79GdbmhMiqLPsaEku
Eil987bPoupEQ9Oh1NpeMH12MIjk0tAjpJao9IL1GnGsV7XR4O4Aj68mQuftwZkrbUVet6kw4neE
pUWRWi2YpS59G64Oz/mlbwUI+IXPIDXbQAys5dDXOf+A8lnPMwdWzS0kYqID5e3GnUYCLugowp25
On8NmBiEP6OF1bxcUi1tujUzs+7CQMyjjJApCTTLtJKBK6HzaJqOjrl+aOdGDdIRdd8NB6/dIENq
06IHFM7De2E6chKLRLdZxdjZBXwUyJN1eB9PutxQReIejzTBDYn2gMm5SYG2oAJrz5XD2LFvM4zV
pME4S+m2NLoAO9Q7FjBZLAsOCefK+WF850pveWrMDcCCObcU6Q7SAo2fjncYBtSbjTspep5Tp6nJ
0umXkmw5c8Q7gkzOe6o5xhqgMgmMU6RJo/8gr/IN0B8wCfPOxdhUnN2mGeAEcAMi0NMCwMDwnP8S
D6bGTxMT+eE3aF40WDriYafajNjjTgnxha5edk2imbPdlQVNKjvv93vbvhjUFHhy4eGH7mBw3KQb
XNpSCi+bKxwFMoyYpiP8JsV4H5vaEqRHc4SBp9mUlcx9CvIQmf0AdUpzMmoYMrb4N+wkq9sNtDsN
gX9FCm8bf5qpCDBANUv69gIJLDaM5jpxjJ6HVeEuRSSToCk3hiZwzfzB17Yo5t0zfA1bjggGDNGK
yrBIkHK+S8bMkQmjP+E+ms3sdt0AiF/+DRXEwvag3PPh1o3fvWJa0DstCqE9oCEWq9RZFodYGjAn
AIG2kPktX2b3HueS34Vesz+DVB++7vUw8af3PKx+3EXEHt4YZeen3c3ajM4XvDIhol6Oiyb6UpLW
hdFhUEBsGJ03E4vKGmKapWCDB6XiycHHw+OeoQM9bSRSSMHeLwb9NCz1ypzJPzZSwnA9WqxToUnR
4Z9adJYApXjKJky+u0XOmkdzz/IsjOGgpTZDQxXZiVjwkexbbSRXmhXramS3ry0pjOjuGwhfcHwc
0A6zOSF0vQXsVU+c3se79Cb/fVOegUndmDv6pVEDy58sEaRPqNGjXUW8RahyzXApEOsHZFMCbuss
u5qPXHffCFRok9alUqFNa2Kx5xh0zc/uw9pmjJgS4kWwsNgBaFDr/fCLuyBwqAIDWkyG+U3F947g
G6TsM+qlNhEOIt2DomRloE9nih5uuQ5TcgHJYAJYznI/gqJtNOOyDfMuBDyecwyQ/u11fB2c7S1a
x1CHX/OThVMIvs6/KLIYfe9rg86FFMk7nLlFHC2/UrRux7wLkDM3alP30oDv/3jgnLawPj2MF+8i
89BNYnoqH3yC4tPcIA0okfbBO80cQyB9xPYEp8TTERtGRFLPf0lMrAmXf8/TOPKopscAk9Jofb0n
k5NOg6tkZcd+8UGsQFM0y/ltglQPEdWmo8F8LdzV1zE0sLa5AkBIavvZrNyva3n8qLI3AmjGM9iL
a2TcNchkULJufti5WRmlImUfR3DET24AwlaKON4cHLawdzQEMI/dPjAujT3rtaBqz1JifwldYz+U
ol3jEcgIMSrOxaX9li+PnQfDWoy1Pb2MkZXYymcNRNf3sFBJwc1k7RlWy5RJSehiIVoP665OuuqU
szpgvXOgoYyziwb41juVf951irkQCie/VsbzZL1/WVcQdvRF+sy61sRMdYhMMDHeII3+Z1L/3IJF
AeTOmScoKmrmte2Fkt69GQKsXaX2vF4FMau6Kj99es6qhSbnl4oGCDUYgx4AYH8VqmQ9vdzFEjlo
pG07ImWEOEe1ie+pQsyj9sGcq8DkWRaR7ET6/5+f+UDjp/byFayFe0ewUZ1wPCAOyiOVAHWrRYO1
PiSLt5lHFQGcLOBWfabR//+kkI78FkVMmOc8qIHkNDcOuqV6rw1p7JBGxDzLc1ndNL/D2XzuHMmA
i3bNPyqglp6hvJbgMOiHuDJEV38BuZHMefe0QNbJzpjEULM6RgDIQ5wu86rXskWO3LM0hlfXoAih
6UW81dAoELgkjfEw9aP9sQLZpNSjEjUjV1hhAUHb1Hyqf0JonmRIzqQNg2HPL+E8tcUbUplKz7x1
3ZUue1PbMNhGKXWWaM1XUuXV9IfXWQEBWhbmB6lDzSuV8vcaCvRI+RecSd7/C72CuX0FgC6OFqTr
hHetbQYfhziswwVQxAeQvElX6bPh7rTK/MnlYrNUYrxYpWxUaagK1fWzCGnlb8JBKd8uVw1giBDa
tkTohvS0L/9AR3gMqARip1BiEnPheA/ptwN1CoER+SgCMC6ix6594MKUrwG9ZBZ/69j9oNQNJyhK
PD0kMI1QUpUfl2rYo5kqJxYo2XWBYOLb3fBO6mxaLXW8JuUxURPaZlRH7u8ZI6hnlml/IY7SQu6R
dl6/4+C4g7uU2l7GQaAD/uDl3fjGmZYbSPVqpA753y1Zk20bQIh2F+rElhSX6IqCCynaBo0NHiZb
IMBm21JZzZW1dpBmjuEAnexR4InBY9PJ7b0gcQrC/yeW61NPC6lI2WZ9QoVl2v7aHJ5oBDwSUP5G
TDppCpVa+DrOYOU5DsqzdRinc39h1t+IWH2AaJA0scohVlSHrGPLhQF0JZ3UcJKN3J19h1Gpb/34
sXbe7Iwnjd8vQXxfP/Ch4TIX0sq7zURI8BRCgrBzz4oUl3rcN+ozjJuuI47vAIn797T51a2Hr3ii
a3S3SnCDWw+v8OIlwuRmuddA3QSar/AhzB3U5JAaSlgANOQcqhubPKRwaRVfoPvhT1fDvlBWxJYM
PpT/dkQJEtLNALhmn2m10VCm4KhrFFLbT9AicPedLkPux7m9EOalugwbo9kxqzJzruRk1Qw+9v6D
xDB32IgElXpJfDG8mI1x5rPnayX1+sGRP9MZmMbOxY2GKoO5C8ozMHodqBfKbdvVvl4BTB0ZqiW/
OLudh4IG4Zg07g0nifrOmmomT8Bswgbsp0shMs6BjGck3+SpX4UomWfjWB56pLiP7iYReE6rItTL
m567aYpYXNG+3woHYxWD7NbFNIuHT6/BRI7XTQIydNlREd3P8KEgKsfLgdS1Id036e+uHfUaZThw
IF+BwjIozWB3q99NTDoa1gU1EzDoZp7RShj+IXjh7Z+PcLp5EQ+cmD7Z6vQXsfe7mR1Z/hc6wT5+
qeH6rtGyIFeyE+6vRDTtqOiD5oylitLQfpeWlBcBe0huIxsm9eACH0epXGcr8ctuVc39jvKWd2+x
n+bYHU9sItKacLvw+0hLKJxusiOjlc5jm4a7Y5govqtRCmHWR7n4t3zkR5xORaUyf+NCemJNvjEW
AFm31nVrNIQz1E4lP9X0F9ICjl2haxyAB64SAAKJvMB/71lm1RUqRklOvzTi5zxHR2Jysgo82e58
nlvWsg87wfWO4XPhmX1gaLoL0H38ZcbkajVHumH2q5eHC1p5PS4kGw4QDybqbMFQ+nKRtZ0idvrw
oSXpN9eD2q/xxCwGiHy2uereu/KX854VicJjC+hK4mzM4XScgXbvve+9X2XP1WN6gRlpe3iB/AiV
KHhglJInVzbTPF8IfIvKKqIPs3TVdXLmA5+YU2qRM7OY4r0C4mqEvJymqy3JEp5odrIpWCR20iP2
VWdwRE7Fc0R19/6b7AhqBw8NyHYzsRnQdUUlhNQHBRGlm2yWJbksOJsQqPpXTr9/rkX5qMjyb0wa
8JKyYzAamVOM32YGLW+PTpaluTJ1zLjfld3K8rG6IDdjfP2GDyIwhaWFE5J8/jNcqWsbkCaxi0ix
BmZbiYdENep7bXooQgZcqDXv50Su5fZ+eGyLJyNRRVwQhIDHh6rdx+EogSZqcKvkR/9g75iBnTGW
gf6N3+poKUPNYHZ7aJs+Hlwr4f0y4HsNqW2O9+cIZ6VP68muGuRE2TnBTzgXMcTZiyye52ZH35uk
23daDiUNCRdzECeXIabQlHG+gTMR7+EjROHk1/PwY3HdG9pJkJV0hq1CBQANYAKNc76NyTFa817F
GTAcOsTfWxO4Oi4FXIEebynhGyJW1Vj+eH3xXWCcpNXTT4+6sWh9bCcIm9r9hofCvoxigHHDvW7x
WoZnA9ZfW35zIcR6gYeslqYwO47TsJj3tX9ghTHQCVmoYazDmC6MZswg+tF2yNLJhjGRSxViB6pM
P1tIoAApwDT19mVNVBlYUpN3c13ESsl55vA3grZO2qnCUJIp7cKQWKqhssQvt1QHopj3YYcu/7hY
VkyQXFYwbddlp/tVxt8h8TPluDto+NHCLPSFfrCvt46YkMPCsCj6s+26Ez8w+mKRdXIKGoMnwEDv
X+RDcubcIpFJ3Y3UKQ0Nra4d9For2ObsdezM4xVduDUqMY6Wy0j/6MO6/JBt25ZW5e3zVumbsLAn
oHgPLBbfVi99rcf/AJAidqd2e4G/Nr6nHsfpu+bqQR4bgs+NSbgOGTQE8sNj+sOBnzaFi0vgjquR
0IrS9kz9J2KvcSgs+OSl9t3BVcb/eWReBiCZTtK1Gy8yWHU2J3r2L6JGwKIDEMfHQ1OqezXkmVaB
lc+C4GRq7gMTzQJsw6jEBIrv1GjFt+BV0G7uXyyKaBsguIv60V79W51+uFoF87gJjgLA4G5g+GVi
mk6xNu4KsPhThSCB5zzX639k5APKI5As4ubARNh+7bnJk2I30uHDoflBpu1yeEaIHDOLcnZir5N9
fbY9vOMQfU2tAKKUWaMCzMGGCjapfRvzQUmdpbb9ziEeaFDxJHmI2wJTMFcM2ODDeohwhlUSGC33
Ljqy7SWRm2YKG+8aIIO8cltbHTXYRWVaceIrmLHWDOrZvGrEBREoIP6rb4RKmlpOn7/+SdOoLxvx
mwREZHIirbUG1xbsuY0qBUONoy7Pd6pKwpOG7d9w+wez4zTN7LRnEn8Tljz420nzcdKW+SzHkNTZ
wJ+nCwhwdSxmUX+XuPP8LhubpQG/FKoBVKnkFBEC1OCZYrXDy81acHAsqqSMYFLuCdvnoQrH4FXF
u8o7yNkh/pNaQ1vc5GnCd9O5Ffwg/S8nrwsDXy6EIrMxKEfOiyBn8HYWHndsqZgds7sK2q+HdHqM
59c7/SM9rXeHMZFi5YeurpwwpwjLpjoNQs3+jFlNCc2vYhCSyAUJ2330SmPih49MgoFlyaO4xd/I
bV+B+moGREwQ2AgdLB1p4ELAaFTkK8iOz+Xgarh6/KfsPTCIQI9GDWXZBu7GC7Oht2vkyagq9s1T
9n6iaRek9GsI9JsNBVzeNYaAZ79wYABlk3NMUlvQLP14uIy0REjzjsIkLgcfott2yziF2XzwLMUR
bBfWt3mfStIFEGNnYKLf5c8IDpyv/wWDlCrlroUDr+zKIUbftiRXRfnfoJxKOayU9PSzJ0QK4/G8
EkhafWtqDRa9qjhTP7apA6yp6KUJ0MHetbQEbM/zXaEpru9aY1UuCWKVbthnM9puiONk8JtkZuU6
/esYNzd4/y/KHjzH97rLkvVhEstODxDGt2T042OeG6yTOnmX5SRRDHEwE2FY1FJYafKYroXGQ5tA
ETqTmJyBRgGrnAEubHU5PcXxy8nrIDN2bFhBOLPGwgZvNZgXtOgA0SpcD+Y6Vi/A98o59xWlKU2k
PABHWugvpzsT7V8E640JFX79SzQA69XcMRpqjw3YKO2zlrd2LN0vxvuOtCQTV4KPYepJ1np+IaGR
iVF2LtaLOJNzneETzFpG/YSrQ+xEgV1EBbF7E+GbygVomH9i1CdF/3flLafjFHl7Yt7Z/6G4VMWb
FVbzV9q8r7hVBB3Kvg3h5MW/EmLqxIQIF4F9XsuPKccT6Q7AxF0ZZuw1Lz3DWKA/K0E9NcBQOevu
YWTPn4bx3ZhatyP0d4FvBfpqI9Om6TFfylVwe6MU4Z5hmte0JplDUrbFNvO0DsfzX2oensfvPqbl
2u4idJsMPUfu1XJ9Ghxt4xqTenuKshveJ7w4dWDV1hewYUtws3U8XQRaPoRVWN7BVxhIuUCDh1Np
nkUS16gjmu30PRd2swpnpxoXs5ncDsl516O4hI2tpq/XvxOrrg8OYyay+I6hBrrFi4AhtyfmpWAL
ZFD+9nm/Nm1tOHJ/82RMV5AmfDNOXvPEEniwIJGJY7+PVyISPKsROxgIcZhuY0RSzk1sgHz/6/Q/
EGU8ZGkaZA9c5ncjhVPKJQAKCXotTOVu4M3mrw/cjV2rMnbMQvuLbwS2YyiCrjANlsiLYRDvbxXQ
M6UazaHpA5MugK+zOtJmbJGc7Io877YzZF8s7OOmgniyK5OwxQatlM+3jsxtyV06Bqt6V2cS2vYG
kQaMaJJ1ZrTwvCOa+1hZSgqk/6HQYLktB2fwwOvBJJGSS1yGATuckcc11VvDHS7FPa/6CEIgUElz
lB/nnovaRdV9hVgvWlm6yyh3SK8HqVqeB7ytRkMQ0RjaAdTub5eD5MXJTjbw6W8aFJxqHmaYJ9hQ
AiR2ADY7mUlgpaARMezXZK1vxhAYx8Hwbg1EswNHHrEDThxKAbxhMkBLhU3of7q14y3BtklpPnVR
2YyFXAV2A0KQhxVKt+8X91d4VXT6mTo4pIbZx9zjVjhk9CUuXGIT5xobi1zUNBqvg8Dwju+iI0Zv
eOC9JManjsr0oj95ZAWA73aRH8a2lej29tNYNTpzejpCFK66NNA3vHkf5dyg4zg37fl2zgOY7+Xj
XoD/+2njqwBl6TmjVGQmzFpFIZJgsUtvl2YTNR3gMaFTIKS2c+vGzKAcUpufStsTqVZDy4iFk/b5
nORC/5Bv3ycREBpW12XSzMqqjzsj02NAy9eIlVn8LaTaNUtwRqj5Be1DrRnXZGLUGb8J9HzstamT
H4jVyTJ8ILVgksnnqw0ok7ryicKo4wu7Emz75TiAEww7MU8uNsYdd1Gy1cZiDhugnMso2/XZ6ku+
f0yq4f+s9tIk31hncwqUgn36iU8ui+z45gbIyV+3Vz0i9rkkebxz0OCDorgXxhXb/lL27SURAmfw
XuWJV9EhAWyTIAgxxjmkdJ1opLnn3Sh+Vl3MRzpPeGWLRX3//MfNPILv9VL99RbrsqXr7pk2/G3Q
4rxaKOcsW04dMePxtWwotmx9hQz1OYp/VtUpt5aqF8Alqb53+vJAXb+1OUJOq+qN1ykQQyYxIgCx
r0zj6QvV+1+qnau2zR2tX2EPKcmAvUjM4XnyU7UouIVrnIs0r+1m6kUALM/EN4OsoQNvmHCw55LW
l8DEBiYNmoGWksFFS0r3ruLi4uhfC9b29i9Z8fYTAUyRGS4r6qQBkgfhSl26Vfn0kaOZ+ZSYZXhS
eD5B7u+hO36rMEcmDhstv4eVpBSvmeouT8YBEDhhlhdacnzMGnMCIXnWfJX5UwQBGurE4k+bbGcI
Qm3GwJoDHuOzV+cI7zjjAfqnsxxR8tWGVbjM37c1GJIaUr9tThEQ+cVL1FanQvXajVMmGJu0wqTT
2ao8Hj4RlWUurloo4VYe7Buyg6GAg7PPo6kDmWJyH48AB1HclsKBPEKy5RA+2HqP6cUFMTeICzVk
DXW/6nVWMUnJITjvSE8NFZUkRuZorGEb8QAlSpl9+5vnXLTzhEA1cdcVlciGx9PVd0ybtsDl5zJ1
ajl8WREspEZvsNwF1pJJfIv9OH3+y2jUNnOJIleDK8PPcbqEZV5TuiEH5S5q40MREVdgGwOLyRej
hO3+RLk5rPg3Lc0QzGVRTXxmshdlJexl0gZ8WguGcHW9nSU0Sahe8AgVZGj48bzfpsQagqQvDLSx
WM89bUoxv7+jBKHZJNsOhe9hyckmNtIuWiV6XV4jTAxPQgUVay1zfAak0YPD/SJO5hFYWnQad3aa
tR4MAaAr04Dpk5M2WeJdIjHlcEZvVC3NYTBFaGU0n1KQcHYd/MSBQMFTWcV0hw6bu3zX0AxjyX4m
ISaFY18dmyCgA2guf4P+Qb/hgNhDaYkKFghpLr2oZiibUVlBO0MLtxATlZYDyum2LVbWJth2rdzh
GcPbvL7J6G0+fKDLpbZTGKaSNnrom7rwdx9dCNvThIsf3sezFhzlcmutSSDSABNhPQdUL45G2Hna
P8Yzfkr6PSle+eVbYBPKZtpRXT22MIHQN4yG6nsb1TeV297fDVMXMzf2sM8Y1/cRIiZFVh3D24i2
Q6Mj2JAx/GlegfzzzVwba2WzySvbpgKTPrG4q8/2tD8Sx3yFJDqUvEq7sronQOsNUr7wfwvBNSjt
TmDgJoKpiAOZ3IeHkO4iNW/QrF5sf9sBilHhTE0lz4FhkqwkvZq/jDuReKUv6o3f+RLqG5rR3Zgb
pRsOyuLrfLlHoy2SVrLgPDtPmRevHYp9PuKYs11cWt/llFVoNcxfMvJEGD4bexVw7SJnfV26lLFl
S0R/ojwZYZBbw5SBk0uAuiqM+IAlEuRcbLzzGBVlwaomwLsbctJ96exZX7RRCB14l2fbBvOGsgTu
7x6cW9zTNJBBJYDMHfvZ82KUy+4/m4XLOo2fVUu7/hU5e3067VwRO38e9SO1qRrKUs01kn+nz6b3
aZMjmcpYcNy5J5/c3oaI0a5EvNG1D1yDzVIagz9f/NnNYFVNiMMFhfbq4DC24oBMm95pbhML/E8W
6GYcu3YUNDQbqCG5hyn6MI5TsIyzgEZ+HMjm1xo2DPr3gFkUgtpM9hKuiWA7rB1jPa87cmSVzAYU
7fUjmJfzXGXxc0KHW080aORjUZq2/RkPogaYTX1t0myLGjrynh2jpTXBIdcvRrChrYZXKMq1Eavl
MPNZomuoG/EchobTcC08pv1HsTU/ucro6/0DIA1bFeUIs1uHzjpU56+L0uNAdBPpx/O7UUEy+rkP
EZq7IOPOfYQQvl+Q2ZlJQjgV9cA0jm1o0oxdmRIdjG9rcf9TlsYvo8uu0wnccsxQ8fjyTdc1UNlA
tGaaw/23I1HrxG3dIE70prc0e62dPts5miNkUp+gnnQHzFb2SLdHbSrr+kIZ1E3Ua4IXATqk/7b9
Sg4BwholaomDvzFcQ0nfy0HK84O1VIxQ4sVfiZJivMnpD8sXbS5Baha/Fr+PZsPEkHvsmQ4eNo5p
qNlL+3eCaaiT8OgzGMw9RnMNmjvhzfr0YRAaftdJf9+WFildUrFukI53CZefs1eD/OEPjltO5yyH
jTA55WIeDqT60l0SjCNHgA/qT/2hoAwVWe+uE9aVfFZH+Jiui8KbNrWXYcvRk2286WUqgtzFwV6m
lKyJrzwFx/tfEo/sNOkKKYAwSlykS36d50oneOm0K3HRIiFHu8es0BE/0toLVGHXFVq+L8pz7Rbd
NZD4FPCdD5WDb5IA0uuca/miex7HxEt6HuAjwjcyRumV65JglZZNqk6EM9X/KW8h/wlJUNgEINaJ
498N13WEmx2KpAxx0Gs6PTiW/B3j2xrhfn0HX7p171nH0ldqitJXuoHlWtDd2gqrP5dIG+0VwXh+
vDDbjfhzOrjMttFlR1ugvq/OQzwohAjmkM2CczFZ6Mg8IPQPaLsf1wuInEN4/QacpxQGQwMWFus3
ZEoZ0CfSckNYAcZ8ZrkOnrqGZCZyKB+G5ZTyChf93XHSTaMHu8nFlljlCRp4kEI+5tg8telMNbD/
2ghEuTI+7b5X5cyKm2kp0MPfYHvbdYipqB9O9rJk6ka50ZBxhtWBs8j3akKuXcTE0qKl1a3ZX3/c
urYquk7lx/dmG9IfcT2WJ7sR+YT0s/fKVpIqK/iR8VeBZCD8720gEYTCutyBG6o50VXS4Ma1u63L
ZeudBK7pOQAZguNc7IvODBEksPbzxDBCoIB0S24K0vglNffU6vHH76xzhJue7OPpIlmC9UIGe0qk
CNNGAvY1z2AiI3VFmyVlgKoB+pL0vTTXa/Iresmznxvv3mITTHQRSL0CIPnywEMQFGMlpvYiNxaN
QSomNi4kprpSbDbU8V4Kn/9d9TrtxjW1NnQk5MKPGg5oKtnh9diAY3Lxhk90Q2WbquDhmmkEJW+0
Q0QENNZMZfqr3F6SumeUDmnYy0p45wbmVdcuynPfkHjmTwFOn9AnBcxCoxrLYM0OUPhL4q66m2kW
0ZkARLtprdVfRbO+Omn4532OOtDwa4vicV8+bufwmSWFY6t2PAgJxoRL0zmRMAT+O6yk6406tptH
N8YhcrpKNrQHK472RStocK/3Tf2Rc2IAaggOus67mUQw7hov+7xrR0pgNmT+5uvPsFmPbxyKht6v
sp8bIStQWyFPNw1mUxnQYf89ZTyqjkpYs6venYnE8cOVS/tZNpTcESEPqi+hiRFFQdMft8LvI5iS
qcybZxB/wc1vZT0v3wLSsbye1xfcHAkCzEUyH085ZHlGXtPE75WB81k1euNFAZzQ5PTYVioSstXI
tnvwUHaSa6jAbnATF+L9qS5ewXE5mAueai1sX3wq361aQkIGAq9N1iNaHexDNrb8/Vq4zidwl5i0
f1pugQfcz6p9d3iKeRJcX728z7uWqXyNk6id8yFVjIS5rHQaONrlb+DjqgmSG9MnHurSWpoz6exU
uN8etxOBJAjUKVkUk5nov3ZqLEhP7yhe6H40oWlMCGURvh7XsG3LIqbxxfJudNwN/6NfYoHAsMdZ
ZBDqxK9TFdk/Dr+zzUheuCmtF+So3IV5u/0I4BB8VcgfVE/+SABqq2SKTuz3cFuxjrsTnHQPZ90R
FXld23WPAuPMDH+91hlo6jgHO9eArzPi3qmt/pqaKKqd/4yWkF5Q7P3FfmCykpPaaUc2SwFT/jcY
9IICy3OfefrhMZEO4dtwSAvG+A/sI7kr7nfFWjulAIl+WT6w1Zy0tJroK80Q9/ZkeGhQuz6Xch9J
+zzqqd7maOsb5tSA1zbMJQO/yDBLlgmoPL+lywu4YHZbm+Ny7EJEZif2Y+hzVcJUES2I+IfhKxoK
V1HoDtcytxw9V8F1PzpTlsbfzY+1Esk1VZLALz/ztbUu0n5y6NbbdI/Uoj9jWWfbf8n4gJ+pAxr7
lgoNpROCwqXnHTbGqwgU/xU8CxHi9srljy+qtbUhj4W36isOeE+aawLjDeqOXUq0ARXUQtzx6ZPP
Yye6aMNDcyohNQTRStI2QrzbtQ0s/mpRb2ujEvWuic051hWFs7rNHD4vAbUlbcYRwbzZikNRErJJ
jMmYnNSMfGvxr0euGowQHSr9Se5plWtu7jaZRJj/jIYrstqdtbQr7dsCK6+r12dCNc8gTaYa9Avt
5D54olIYshNxoYaOoLVOU/WzcwefJ1goG5LOYGQrT+dAy6nMyTA0gFpexC25O3vBVMeIjUsCPu6J
EAYx0vyFSoIP0ojm6oGBUdWyLXs2saK7gaEOtVSqE09HtlY9gH9C7ql9Q1szsOK+v0LC87TFMq0Y
FEKu1IkW56SHjZ/SPQ+UZSIlKUPER4sfKNIXk+ky4FZV9TM/tNQJh1FxKfAe/iHRhjCcQYajDXrj
i95uDwUNOJVTH8nxxGmyboiG8x46U+NQKBshF7RpwhkkmvMjlw2PiZtK8sk4/pSlyAQnNcfVzj6g
1KS3mVz7R0cQJHdWntsze/K7hqTEKRpGTPR2ISSfbPg9QIy1XQRnHtiGeVu0u/Ae1Y1vrLRJFypj
dp+vxdIo5SHfhrXaq0X9/XgivPZOPYIXRq2IZFWOtQWiup5yiPPBY7j8JdNQHvOORyHpAXakYDbt
HEdBQfHmnxkrkTTHWDfABDk61Ol93MWGzxtHtU96GpmxwdK8PacLEth/I1zS5zKHvtPvxb6sDuPt
EGJ8k6iKAJOFQBY7UlZTFGjfI4Mt/oBwpsRL4ZKJBrt4eSjFP/fQsf0PgbqnqRkbXBln5XBtJCyP
2QDU8Loyq/zBKiF+hvgU8vdxzAhS+QCylrBE753NnnPmc53F+GgZG4HFq7mD01U9gKIN2PZj2xsQ
7HMqoshMtfLXL/ABrkViujajrXDGVme8UIJQXMAhiZNM86TQMmREQ6ZM9e3jY5AiEWtxZ5seYwcW
/EcPY9orYPhbeq5s7H8ANFPElluLjW/dwDP9FCU3XTvxCNmyzkIMqzIfofH2DEIDEDsYoE3XeVAL
n8/us6D3SuKEL7vL+q1kfZ/U8r3zJde8TBDltX1pFJMhBsu9Xzwxfmy8Lie11XjAJL36lBnPAPHF
FCk8EX7hLmaGo0IUbtZA3838fzPPZoN2oFLM7KertdFUQJgUA34d8M0ps+EzVOuvTObv31UqEAwB
U5z8OYqdmHx3rJbqO+yJecWcCYtEgRz13ZKN6ZdgaCqRf3TgPI3uQUi6v5NcHEvvhP2rn90H5pqt
f3hZtPKk072nZdDm/2wTvcGPiZMcg5eWCOKgsqjr2ua+zeFbfxkXBq51AC05oGLIZriAMYJh+UNO
pndh+YZ6VzUcS6SSFtLkpUwLoc44hHRMIxt25Lm+kcuf5YOoAYHt12402wjARv7cMJgsfYOLo9ud
zZfN+SzLeFzGjm7Xzc1LmA63F4TLxwQOsO3b1KqA+DaKUBRl8oUzNNNQSuRZDBIbrwuciZvL38P8
cn6l4a2fXbvB/S6mjJZ547TebzeCYioZ4iTATpe7skhvaGmhwhu5CqM7mCqVH/dDvpBzw8UPWzZV
cc68yOdANQggDMxUilAUue921ZGV0koce1Pl/pUhYE1aNQMBFEJ8DN9Q7fISIj/M7XU3ZdfIR4Be
LZkzJMJpLoqmXxuWOm0ACBuj3yygr36T0LTebVnq2L1voupM/QaIZuToSez239uRllJRxzJKIwDo
7yOjcKzlPyxeS8UkmAfBNj7fKnXoFPBr5EebQca9+bedNGRvoK5x5FRS2FlfAQGPE7fFDaZJAYD/
HTeXDFeJDyVL5iWFGBs9qCVCIl4k1no3RAM868jtWUhkSqDwyhRNbH69duvjB2+D+Pdo1FVvv3mG
gOSsNuXR0aH/2j6+Ci5YluzpooEiw+y/fBNj1AwImUdqu0zvtTQVs9KW9UfsO6UDY+ISXZznSqcG
7EvfTgRcL2RpPy6ApgBJysXrOdGRU7QHvdYk8dd1ipv3AhUlIP/pLEI33pSrTEmSRFNfy/kvUZaB
7FTVifdi0awz/xcxr9Piblmp/WdI9zHAPHSoP8g1/HzkbiH8uTaKjRZvSPuXqXPnjgdGX+dbkflv
2eZX933K5TFYXmSvvvW0/FTh4n5x2HWUOZlmzSBP06TM4ctzHYzPGE252+0aEKWv6tmwgCkgncRz
e1/Gu5N122cF99ZWBb7zPM2i766Ge8SvYV2wAIMMNjZuZj0BOsC8ZQAAqgYxAIJUIxisS1eMK50o
KMH9Vho/3GA3CHMWOge9m5bakE3mXpFeqjHno+HR678uVpYCHxyFCz3U+Rhq/vC3YrDPSJN2CqM5
de9HLifQRnBE4Bx/RTkqisGl1/jQtvemXIz9CwvxqDQ7BizwswjgxPcbcIPvJ2zD7HtR7W+R67Ze
F9p7mS8FiEskdZVjH+sstLs8ONeKBSU6POqp+ia456Nwe2spc/aoV8agroHSOG3UoqOgONZbFEUl
JJiqF1DB3vkFIvDxDxa58cktVwL1CCx7oVVPiC7/GHbVJhr1Rr74g9/lFF5e1SDXMNNfV2evcmZ+
flmfdzin7tB4vUjrnUie0E9ziQvuQQlRsaLOkFqabso+2Pkrkp8RO9U3KGSSzzqWsZHwUeg0/295
IID2QhK6Y9iYNLuZvD0UiOf+FeqvtPw1+cCvgL4MgL+JS7N0eFirLIEj24Ic0EX4l950c9yjIpoQ
/IsgliXI0E19nf3b2RcEXsSZYTO/FOmZ02jCV4TwUBGSVt2cjBrNsAEVTxD0sXhIdsIXTPs5adM/
/k9Wd/RqORgal/xxmeX+Xc/UneFikKNz9P2QK7n26ejTQ3idcRC6oUgNWYeN3Bq6J3IN7GLhar2v
ynsc+omr9mGKv6kJHw59lKEWNU93c1xBPpjo+ykDupa4m/Wdg1NF67axdzJaSk2NLbmxLVos8Jgh
WX8R6R9trWoMgipWsPirsII9ZIsabTX+6sY7qKIx4Eo2BpjpRQwdw7Gmo2GsL4fUczQzS2sIkYFK
yQeSJrL4gySbc7pfrVx9fma9nJ1iwhe4VQ8LbOFXKbzH+BWnZnSmV4xHBTOCKwhcHy6qjTz4AgYf
piSuGiAMqe6NuatddPsc1SyaUi6h5vtaeQBFZ+L/sxPr7HhxRRk+vQV7OCw2zLw1XPquvl5qTdbQ
QbT3gk7fppCT95uMn9AWR0S6Y+kCIGhxNkds+RH7FNnwkm1hMwau/pjdvv9lYGllbMSshPnGBKZD
JtfMfyI6pQ7e8qSY6xUx2jQOVdPhouFioxHjJeOaVozyRa8baWAzOctE5cK/onjiJt5Rd9/KYKko
9UE7xk4RIlEQtLKoN4SY3eIIF8GHBOMzh4jV/w9vVH8hUwjZ9KybIrPbbYUx/ZCjphiE+Uh/UGu1
sKrHX6k9zKjQNZl+7FrvtX+/rL0/JhpHJrclpQT2nrr4yK+o0/QQXFjxNY/YXL7Ql0d9ev/myQm4
7pzyhAzaDpvRV1IPsCq/Yt/TpLSRxY6Z8gZx+5DvbLn93rkewK6Odh/6KQBqKnIfbJDI/NlpOHWP
Nd73V9QgxgzKWpVWtGb0Y5aJ0duob9Z3VBE9oQcY372DfAaUjt5ceifWNWEpnbAOJ0KzRqbEk7HZ
sHR5EgporYFprmqrTDg3LofD2jCLwkVEz2xeQz/e6+gnCOGepXcRYkqxDVNe/JYcLclzQG+S1HlT
JVC49DkwLZB0hZ5Ez1kVn61+pYU7cLVmU1bo4hCiCMcmK7qMZhjs9buwt4KOXrumrM4KZmyp6vaX
FjQ/dgDdzLM1p0HvK+gJH05QKTyLq08UJzElDiXgP9KtB8UH3cgyyXZO3x2UVxCWDxayhQKNJp4t
oK3QSIW/j4sLZu92lw2m57Q6eFHEBF2AkAXj6yPnTHhMN8DKPAORXT1dQFXorzmsIxatcndqWjYe
jWGpgzVyzA5Xsl/DswzHlp7X8qoKb5C2LYQ0+nkRHSJCQz66jIvU78anj7FV4v+xRbUllClzLBas
i8Tq0ZHBPZVu/Z2cXzvausFPlva8x5UXp509GoWmZPjmh65x+8j3ZQC8DyKiyDfBu6toqziKoyKa
i9b+7rB91o9rPOA/bWoD3+lF9R4lx4Tike+3ezXSJJATfvXA2MkQ5qVTT+t5KNJTVqtGmI84+KP2
Ni9qWh/FcjOzDjvcHKleSnZKuF0Db7AjyQTMs2rmJNgpASIlIHMPA04bQVOejh4uFSDUsJvdamn1
AygkJikn5RhPpGUiTq5Kt8diMfbuIXj5eLS0ANmm5gWcjnvGbMExLru+FF0n7kx4wLvhDTS0Genr
r+MeVmPGbFKGDpQgN7GoxrlJRoV0dsAx0oMeDRdUQgnJLbcBi3uUhYhjE7paPW/YD58zU4Hbg0zM
RN79RGU1jcJvH/1VvspJODvEQ9WZRIy530zduerlABZB5H8B/U68/7K9/LC3VmDUSZ7xDxp050i9
S33y4clcmkIVfVYSMTfvimtjlWkAFUmSEkb7cLcc6BYb9pjeVZksEC9LdUWrssgDmWcwMgMSOOkJ
d2X99/7q77s8QVr4FdMvLYLxDaDZaqk0U9llBrR12inyEts0ngXh7RlD4kzGyvbbTMKawoi7GmZk
LK9EJ26yyQ5m0XDftGoTxhF2NGT7uS0DEK8QdCIP1ZaQshrqptigAytos7ZLUkUc0djDA82uGVBv
dY3ys4edN+0Et0X4iqh3C99OwIlU+scLsUwoCQoRNj6Wr7KLsELjOA8DYmdGA7kC1bDiSijqpmxv
W5x8Mrhl8fK9mVH3V0Wwx2ehwEn9TEf9RbRWUZvXn1PsckIDrtC/A6I7ZcK36RqHNm3NexfgFGzo
cQn2hb7I+N6PFQ2wkFBFoxd5rDlcIIW/pFWUuTm+T40sfutHz3j/ci5utlm/sY2Mq0VPjnMKgCfW
RIcS7jcCMncSjp7Hl2WYmEEn1j1susgSNKNnMY6Ni8IuekNIeg0Fa4ebdzbV14s+A1C47s7Lw+bN
ncR+oWmQRAPtHxGZwC4ufrMw/ca+ssiDxftqEPjHOIt5BCrmozRqj69cW8DPFUapWNgAZ9ZUQuXI
TcZTisL9TARv2+PaFZKP8uMK258R2CBLITHN2G5ADBVJUgRGw1vpmiThlc4wjwu1UcXmusJDIDCN
xEZeWC6mNGX7WR0Fi3udx9FP/PR+ZAYUzoVGsQRte4zqw77veDYVma/wHwOnPUjo/0u8nbuV3ief
IasD1YvwcOsysEvCQJnCUROi9JuYiHRU6xzsY+lYWni8j5o+G+BRA/U4qaxt+8rvr9Ax5DMRuU75
ThNPCXTKJfrPmLn4ERzc68RUPLhhIrlEKI+8guQqbB6GtlBmSKi4tY+vJSN4lpmtrwbWPm5t0KE1
7RpwiBYosvr694RZD98jRZjhzc/HwIsud38wcOnT7Su7Ms47xWkxgpS64XpxcNw1kN7BJQlW6iKi
6m4R/uLYSWxPWTxMcM/5ZOMsrTwhNgM71ZDhLiOGKRdYqiH6+pTCbieTLX2k+X7vDcc3LtWT4d6s
v9s2G3mK9jlkVfr1gwhnBN8NfM2qcqlDvOA4ui7hj+q3yueW8pqd95nGBepM49SoAezrVNpyZW0r
t2oJOE55agKlYpOHhM/LGSIVQJcZyhKMkqAnQQtw9KrZR48rjcNEQQfK9sVEGT8dYysYdht8bpkf
TU1mucbQpeRo9M5Vjw7JNcoqcyKqY51gR0CGFClzts3K52MNvUfQqmpOJplzaEsO+95mS2dwjuoB
56QEkCaJY1B4MzcRwf74I9fGNjePUNVz92DSU1USb5FhO4x0SK9Qv7jSzbBzaaP9+r8WjIOtFo0/
AvtldfTf0OqxboNgfkMAVEtHTPjMj0+GawNiFNyI1OwhxoBHWE4QXINo1EKZua52kfxTNAaI5d5Q
vLNoOzgykZ0J+Cfbtif/3Dj24I1nHuQDjqji8TrYQ7L0IY+EsksS/RX9dTPsR6THl9jtDuoBMX6y
FiYy5GpV5foUz0Qz8XuMnpWHAt9liMa9XhOPBrUeai4sZw3K2I2ISQXlZ35nmWR5YBAHHHoHUrzr
LsHg7uUrsHUi6mb56xR9NLGyAm+Mrj4oW7ZR9l/mtqSHCmvYnFAgeuFU54TCS6yOEuDcMbbNOYzx
UL1Kg3q638FSCCDvkzfUcE5vBC21ya4gK7EwtWMLX2/BwHkXlHGJgf4qFU+CtKTLr8bPq0BQO5uu
uKi4hL7dj/+z/UknrJUGpvnDF9LvMP8tX4U4ES/zt4P4inQrSldvfM2lgPTu8gsupo/d2NhR/nsi
6Et6tx6t8HpB9yW3faX1ZupyL6dW5+G09oH6uoGHTI6ShNNMGFhFL283soaY/bZL4kpji2oqdWlh
9YQViVpHLwmQprV7Cdx9IPpuqB+qnM11AvgvPGKkd2Bxn+1PYe5nQl5Gt8OD/vd+aSJB2UggitwZ
JmilCvuXsjE6mjWPOyKoowss5dWoi79LynHvjZDvueON4rpP5p2nzUukrMd8VhNDfNB27V/4WJQw
m+IMwBUauOO1Xjb/7npcRmn0XYIP7KUoj2bfh2LmeZ9s3WPvBTTpG1Q9ZQZbpRWjBSNqS45HQlrd
494Uv370uiAEvpjDiLM7u10MliAtcbd1Moo3/jHluWbxONR5NzL6nB0yreM3GJq8d5PYOchx6S9E
T/rOSsnXy+ZyCpO3VlBJK79kkJOk5iscsf2z1K9xftkRjohVzSwPCZLIlEJ4scyDP4Nd5INAMadi
tGwL5Dv1wygnYZM4/GkfLo62AIFjhhG7P5/cNwa87XkRYeCHBXNYfdVo3FVk9pYZWvAAlooCDKwY
cYFwQQwMrIW+hwUoKOs0vdbGQBQa0FaEAaAsseRmOLAwpuU8bwEXmuNNEepus9xYPXCcXtDY7TOY
daiSLyvTd4EilQgcOrdxS8saRZz3ceIIVd88WFT76rG9AT1gbpyqGV+C/0kofZZvaeBBgg3DX4mG
p5/2en6I+gqr3H129v5oGs+ilSo7yn1bqDpx21N9gQMODiB7ke6URTfrvFnINAKk8JnYnPB5jZeb
ad792o8mJ0+8o6xBrHhb7OdiWq9araTLGP98KRrIs4GaJtZ9dDLLvmphAaWoDCaxtplXKwwINMlw
dkuLGGCBYtRqCJ5frYi6k/zm729jHUYhXsYHZGv25ufYY4y7s9KXL3W/ZK19ZP3nHEMkzSrRbhs4
526/C4akjyMGLxvFUmnjH4CWT+ZwaTNlMvqXvg4VSkb5HltSUi+cnYuMbfWSkBPMHsc49mq8s9Qw
Qd1tz+CLUkMR8vJdIHtujTWPL6pnyWMiiY0ArMU1jg5LXI1/9mnKV+SjSuk4+8yn9vu5s74oK6tn
ddyVgdWHeJe9K74UhaJIWTvN6QO0lo8dv1DoRLBKlm8eGbMS+fjVDrkbkiUDijlmfn8ulOR4DlSS
KHhpJIn9+0EvwSQEA5I4t4feHfLNXAzcTxUfRy+gVsVpfrJiwYEQNlRYMJ3sS+CsiTfPPF2Sj1CU
ALD7WiLLAbu+nYCjChbEv1X66xLXs44GW+3kpwQk/l6K6SnmOqgOMsppLODjyowaDSr7/+Dvn7BT
DhWl6QKldyG7mAFrn1iMFWQGwOQsgJIZECAhhsfNsbtxWfSUV3uJPEKA5qio6N0wdq6voOapbRrX
x0oVHIcipw40Ckg1ABniC5+tsIMQaCPs58wlkDVAacI6QrVMcbU+q2OIx8hUnavFncZ7OXQPopi/
jHdGdfezRQou5fY8sW4pKW0RXlM54nAC32xsO1+/yQd3ekLzb2QpDtklUa+djeQyxvEb8msLybXr
UApmKrUZ2byZg6+I3vq9P7SqyHuqid6Sjyk81Hw3DoWUN8qkE+p2hv+w+tOVIil6LZzgngbwmR/A
8Jevm8xndMNLfSGUisFLtpW4FXy8YKN30nxaMLKfab5Xue4ABYALowrrUmMhwYVrdjpyDxoGhIPZ
/sm3PFFWaC6EBaGbzOkBP5vYKzCtwblEdZwanjrwt6tWXMA58pka4d0c0jVl2P9nwkIP5WM+5Ekb
xp/U3IssQc/wWqgwdMMxgeS3sGeOZtr+IoEFCXNauEcCNX1EFmSoZNeWqmXJgvRTZbPt/QP1LsuV
Rmn5PhynENjfGvIcBKmC6BQftu/vp0XZdTMS8T69rjrxFQvvcQvWy8A0q9s60tXovgc58T/5+QIQ
dTqNleHI9riXbkFlGobwUx1aGcaaSJCT1NwG6iCOkrdTOQiypTs9X42+EdgKi9ob/7cSyRASywcn
ybk2kvKTVvDm9I5Ck5/J9BflG7RGYFEP6IbC83eEwQcRevlbWr+hgYZE483TyguNIZxiUxN180Fd
9gzXYHFViJsuO6O2nalQfnN2CwQpz5O9tTHNH3gEtMqepA6la6qbC1jX9RxbTjFJswSvIDD9J7tB
lSxdKiCZy/KzguCtiurjUAyQV/mxmcYJOHV5GRZz4AHdnMHa3TJecoMga6A5Sq+6tGUfch2vtAX4
j2+t1VRyWVVohohwY+paxK3W7WGMm6ouAaT1vRYBFCsbjP2iqsXmyduuSjYCkVKbrnhgNff0GC12
hxPcEMbATB+aXM6wfKB1lscrzOgPYKKnchQMVj9wwD/jPUVxqN39ltbnHnBP2MbBaGs9KxJxRxds
6x7muhNCKOKOUjfJwHvem2h6SnoEDOcOkS0jXaDv6Z73dObPEXWTZHklQfJU714zcnt8JkRtsC/9
7nfPsFSPDNmEdYl94sNM9uWYeIOIFx0MeSvAm7wlGpRiYCK2HDdPhVrlrFZZaWVbGX/nyl38OpAP
Mu/HC6z6KMcXLtBI8CHI1bpedDNXEDe07oJbsMXEyFONb4/4hZ54pbScYWtjmlFfEqTsoDdU+c3X
0gjeeybXygjGn85wNuA7PL7yN6UHYjAwNtKcogavxOwbQ+5nJ7dJx4pLzduIgErUAQ3akzHTgfY2
wEpkXfsbx6ILDIBiLHj/F8RvLnbjL50wLvadWjNkOdWoEOJ2snpW2pqWOz2W71bY+SNzUh7n6yLp
cO9sx/OewMGhko21D3wYWESG9+YK+XrosGF106cFsHZU9HR5JBUIVuL3Wk1BG3eW4/hdDEAjy2Zv
2ZEQ/m0CiUI2oks3yFbHkKkfxiDxDXhU5LXhY2t+AhWHwnOXbH4wRiC36TK/Y6dU1V1f1q84LuwJ
5YmL0mbFPMiCEK+KUpN15KObD9hbuk4flezxbeD45evPGAO+oqw6Kyxx+/zBKO4JKMG5pX2e6ibD
YNxuwGwe6fkWUWHsa/usyjLyhlrsFKSEOXLG/YqsEl4x12KPtayC0OC+bYe4+Ibp/Rem8GlJK03B
oQIgXtFNcwkVyYvtR07nr66a4lOgpXdymHgYh1ca0f+lRWYf1AC9NaBuCeL0/D+6Mff4vfGYXUtb
mNB3gSb3FEns77uz0d+I+0vSMIF+itnpjc4AhPelkzuJKwPHk2GKdzessbD1vbOcPei6eDt84akA
G44slSF2wZbVAwLCdLxY3KQWdYjdca+GiJuBla54UWPZU/bxSGAN0UciHObKIEPaDwuqISnrC+Jj
jGkhC6YM+azj/lotFys/xT/DXxkGSYKbODPvps62dhu+OjPLBhqxDehXojNNjc4Ife5Ieg26SIVt
H4o1GwxTdOfsEWZiPbONWEnX8/4exy9cfPCNiQZx0qBbGf80IyCLi2Kw8SSUobFi7SDwIvGul3tC
ZCHt1Gsaaaw6p4MJkuBxErIb3h5HSceV0p+ew+zH/Mjxo5KWww4LvE+VVs3qQluTkVCyn8vmE6iZ
UbtiQXXEqtfADzwTGVd8+Nqep3jj8sJNWI7IYpLFdQ+I4ddTssVZrXrRcnC13Slm9wLX2p0Tj8AC
dPsusj53iOZnC2VOwO29aF2huFlFE6ru7R2DDT6KMijwm9yBiY5X7NTCDRJgOTpfqt7wEUnqk6KY
c9HRUUFCPFngs3+7+tqOqhnSlCE8MMstPU4FCIYxT/3Y34991MTgPgmUrnG70DHZ3xY1yamDtbC2
NBRgBeGBKmrKO6RnVtCQkXsfaAM7V0k8C6I90K0mOYv/fj9tvOzdN69767cJzPuNi3oAxmH1e0ON
1E72RybJWxmdGL07yKHir9I3c/XogiXO0OR4nSr0a4ls6xmoTgvQKIOT8Ma3KWyiBz8FWWs5zRMe
g63SafXdDqFm43vk3MiIGm7aY58X2ycDtUSF2h0wlVHbnZwBPUy+nIwF1w3TqyKJQzF0F/Uhv2Sc
3+E2Q4HM8Vsp8f3jT67gVbjadOiCNJjglcrZYHE6V8VzzDDC2a2pWmAvP3a3mIPMF7wZzoXRlsOH
T5KqX2htj4QCIfyKd1TXKHUGnAxaSj6Ra6ne9PPjscF6MWsjZcizstm1LLTcjGI6LSmacX2MgJ/h
om5y0w8Td0vX4Azjmg01S/ustef37YAdRylG1mBzIeepE3py+6+PA/DXjkFwMCmcy7krIu66VE9q
Pw69CzjJ/CJ3GacpxZ8bHDI5MctHS6/iTgkL0z53d+44TGyIK9+k0HijQCxxgzapxh9ruiZlbSkm
0bovtXQC9MdZm7PDA5gudDLEdPKB1Q1RYntQzSP/m5vtD4fx/n9q2HXERZebaC6XXFmCa7mya+K/
MYNmGmue/PpXvb7Narc4VWqDC/vVFUMaL+Z0USUdhpsxZ+gT8V6wcYZEOAfhn7PhhIQB9MMCyO2a
DUCSuTiI75qIANWy/8GlMLTB40n8iV/kQytdjKspAJcFhT0FelR1NgdUdT7FuXIzTJcHezWWvZXI
0NS+qW2esphDRxQY6FgfzvjZeJXX3sN84wF/KBsUo2y3ovqz76x3uCuU1SrKbhm1kwCYqcyxubqq
ZIrOwciw3sNEr/n5Tq4+XjV6yZyW3cOi/Tsft2bGgM1xwaR122Og+jfqVnXxMWvD57F2doGR5Vs2
n13xWMmf4d66A5949RGvBb9hjBH3oLhh0I3DCXO9RIJ+WP972E4vtNo4yrzN8hCUBVk0Y0kUJTTD
pJYvwmimASGO08XSr8rp6D1Bzm7krtf7G03jeH8EMJmI13yxxMI6k9X3Hv7id11tJAxAojEC2FNJ
Ezkm+dOpWbJS8PNg7W4kPhxrblB50hQxNEgeHkC1/G+7Alzmev0XoyjosvVDSFaRK/Efu606pMaz
CtVdMWXJoZz4LlWJhlKfRAJPZwxzqsobnH4X5agutXweSDqajf+Rv5Aw67XpjLitqz7l/TViESvx
iYbVTvoDg3f2Mb6DvIB74SMA6qTW3TK5mQ/Py6X8OZunqDsc1rlXao6L62qAmTeXHIgqI3XfoZpV
uhuD3R9SzBWQR+S5AauzfNa8+fYKgqzoYYYb5Zr6VRbjpUyZhSk98K8NCQIwWY16fN+J5VxKqk0m
sWh277XhYzngdUEYW7XkdngI+nRWkhIqsPjNT3ljGXuLDMicLpjFfTgxluW0hD3IuIeDls3q+Jsl
fLDebWIjyiyE0W/HsIvm1XkHnHhqTlbIAZneAIPaPqTCS20m/GOCZ7l1J5YHPRHT48Iqw2OunYf3
9LtRnWXKL8Aq8awThu5tNK1CmHekhDnFd7reyI8upwTt3LuIo9nH9GvgrzkROT9X51IcCge+7k5M
jPihIUI23N/aBhR4OUER5E84aW5QMenmm5w5j0jfWGdCWqSeXq3FWL9ELa02b2AxApU9xURYJlH5
zuRkqI2uY18rlykURCHT7XyjOJrOXevrqPbiw4sR0r8EWLeONUFdrqTxbaBqarp35LtGydFyhRx4
z+x23PUJp3MIaEHFKnImfp5WwHKUSC9uJ+nR0co28LuHNNPuT4ENfqd94Y+pSZNNwCmcRa0C1+iQ
Fgv7CSHGLhCNoc6vn8WR31rvfoKBeimiAwTdWPAso8mnAg2GTRRQUo+EkoK33Ubv0avSLrn3N2Y9
jMxL6EUv50fJ3C61DBeTiMA68wcvj587d1TXECYuq5ycPYejnKW61m940n3H4SDxb0fjRlUtQ8hp
CS4kQtN4tCQc4nVkHpeCQ2WRXQ/b7moqnqwkRs9Ts5RWazbhlX2BHUcb6eOholrDYHDZj1Fr+h0V
cevJThXZxtZ1fb0DYlk8kPW36vRGpHihmhuBahqTvPlEEDPB6GjHRvpDFIrBVCXi66e1hgx/Xdtu
BMPFkufr0i6lAyb2WTMwBVJD6Nklr5/FuSwzuz6CdOH9grrn9PxGfYdCJkrOyzyyin2lEdi33s9e
jlf31IpSH8L612L42KQWh5W1sGfInkFbxbFlfPBw7qL0aUzoHMEkWYoRqRmmwZi1mI7Z5xGYIQOy
bGiZ3YtLTMtynl7EATcvC7DCgweQCYsTo9Wogbp++9MUVXsCjcDozU2onhJrMEYohu8/ebopUTjK
EZkvFbukX103XjSlZqUw6BtB2Y/nZ2QZ09m8f/GgQ/bo9sBr7/Z2oE38QcU9Qndhg+dNBa+/4ZGf
htyAEzG6xHsB6ERmGXXwyde5yLzvRKnwL6LNeUF2yJ8LBhlhpt5log7iB6WBxif9DMABtrclGCCe
BZG4ta83giM+4bKAHbbdhdrQ26pW3Bl3wdGLlcLWD1013gnajE82oaGqr+vh9rILnw5/aUzyr0w2
RALsmv64lTjzRJAwwxdeuuiMQFNK4f13Bc6mJj36c1FBjpG3cQOt3trJIr3l8/RdZLNfjvL6zznr
GkFWRsAj6H0u0vHPjR3EGcPO9fT8h4ATBgniotv/KhUWwOIdIwKjK5a48nejmI/ZneJ9EysY2ljw
n+L+xZl/Ttg+a87Tf3V188dZphDYYop7D8AtcSipoWGVgF35XYiiz0BArhN6/TllJlupnQaNXSOs
uklPCj5gKhSSKS42yDidYuNMLfFtGxPy/NmD0f/aTAw8aPOnKptwsZVWIvKWOckLVYRZV8yb1Iyl
sTRTy8kXknYAyNYeVVBQF2Dgfk8k/KiiYZkE6K4NXlHdE/c2wFgYZzK2HdzekAJEmpjVkEmNaFwp
mMXSBwqJMezS01haUODfe3aVAXuPpPi2M/NBCdgDNWaduF8TSYO+w8Kkaae7cIoQTr0zBnYJ169j
txYt/3JzCp6P9jDf+X7u2LfEYBG2K7/+YeuBhr4ZqWKEgl15SDtE21dCMkt+llqM6OmQ5pqNujAO
9n41GpoAA5ncxyk7teeJe1IwlwtAKwVqfPFXzpLGJUD9ztgoYx3Cx9aLQZg5GFZtGONlkHguhdNu
WXCdYsouG0GJlElKTmCybLv2m9Uz9pD4mw5ckZ02MdBB5xHgkqjaR1gkYyAR6EHNjBAd2LyyR99Z
oFpzvzYVEAUNE1dVMocKS+zei/lEQ2cWSpexE7Kn37V1COpQrzqNb7RpRqaQOLe2BmD4T+jKSExo
g7XvQhOG51S4Kl3wtUxqgyshByRImfmEobDjfa/knbQvu2xT4f6A3Kgwp+hwWZY6IaOa9rma3Gt+
m33Gs3F3dSatb8Ojmniwr3n5+h6DCSnn5tnSZz7dZYmOGN0AUJTb1TE8BhnmSPam4E7atjhUUZI1
u9+upHPdva9BMfVSnfm6Zc4aqFz342uRplCIUoy4cQqIuJZpIPm7OVTCorqpMHRqCFVAX6GR/4ip
rbqfwC4u6N2Xp0Z/RCMRWOxV36FqRFjgjPmpv1WBv/zSRkCg9OeP1CIIgZrJzFlvsDODLpR24ybP
NdgxRVNtF6T6tr6wCrnlI1KZM4pvbaGK5G674DrLyBbR2iClRfCjcMDndGjU6i2j4ji6ewq34TxL
n+9jIavnIZlSi+A/kgCLQY4MEmfqFCHuksVOL2tRv9WUmWAG12jisLOm9w4g/RuMSGkQOz2Si+lZ
MpHhHeYsdZJJcU2rk9wEIiRko9DoQICYi00/exCm0smCJxoyUjkz23jfaSspmEgQSHCncUjiv4d5
lYkpZFyP2kH55XSl20Iob2F5Il81pzgM23btt3FyImmCtmJZsc7MGs5uYr8sG6ln7EnHr9jFEalJ
n5lacCySD2wkWDx8MAu44oZyTTMqSVhUgnZf6KwUS9K7vMYy4YBebdqNSk0wa/qCx4ADN+VqZtOr
FKSQsKc91hVR8ya93+mobnwHd81jumLN5KgVwS2PwXqWTvbBmt5Bmu7YY9J3aDEzFvOF6lLRpohN
k2TtrhGMYd4B/dsxyzK4WHxRNSEVieNgukXrQJmeUC2mPA4c4pEmbMSGNStQSFiOdHisTxE5+h5t
ccF7I+ZCmE7S3PoDmHtJTZMzoyL/Zz1omsplX1a9luuLDQERyldL1C7jSAjhsBJ6jNv3cKS723mh
feqiimMK+oYfwvNThERZS2ysTqSErAp0n6Sv52rhKZXPh2UIX2vkBd3qCoU2PUL/vhtk++/a622s
gBIAG4dz1Xn/1KzcpIkGMNx+1euuR20pol6leNGFYTH+hsV4vwmMJmyv9ypVJXGejH1GHtFS48yU
KHT41qXc+6TBK67UDt5kEjeBgPtuj2pIHU2CTNf0bpFcGJ+JrS3e4kzUfhS5ixbYzfKG8M2iRTDD
YCttyAiy/aBvRFaP6tPSoqWW1X/qCqIsq6Wb7wY/EVO0K1ybXEPqGUE7fWz9KLngl4TqXqbr8Qm4
ayaqe69yZmPRgREL+9fmhDY+ez+st+HcPfOcb1lFswZIzYKZ405YHRsISroXzpO86YnHCvafLbXe
3YoeA3i8HZCrgSWNdQPlqGTFydnt7W5qAyMSFLeph2qK7+yl5swXb8X7XxTVv9WvZJIL1LPBXy0i
W2DjeaJ3UnjCSt6vYQKaQ5yUmz9wmeODTACw/YxtOqH5OTH1AAJFvMebv0/R7Prox9GBirBTdUxY
WzOU0+1IuMjcdqAGiIV3aKwOWgwrBu+tuTDfilLeAr7ZvR4MAtD5Nkhu7QDLgc4Pg0ymlKbYog0Z
Tj2PDqWF5TabnJItxza+mgCYmnke84EAPeWOuoV62aic5XyfYx5Vx42UrftYGsqLwh6oFh9/U34a
uKkeo6gliSuprY8Vc3d1LcZLmbStuAlVeShZ570FcEDUhBig/lU02vLZ1hQqQ0rpkU+Pklw3Xwvp
I0nCM36br7OjJ4kU6y9dOCYVf3fdqTuyLtWqTnvLqV2laGlB45D24e3WuxGCjVEKKowFLB9kRSqb
/K6NW1g9Hz3ruH0a/ZTqPpsOjXagd6Qbtol5pO+SG9vMhxAviuCRoWnGygA40rDvrdSb4l4UOL//
d4fof4ea4VrdQYzZd2Tbqy5ifFuSmtgiRxfTJQvt906UAxGqquJzPrZlpETTnmPNG21P+qepNrzl
vR8dOk2DZ4UcaNyGiANqoJOAxGI8HJZSApRwi1p9b6fnI1LK5Co1duv9IH6AIcCEjdDHO9i87b0R
H6j7iwi6QhOMxVuYi7iksIMu3sOCU+h3O7HH2ZupsAW30J9GOoQ6BCWdM9hvfM2oAX+aRt6sN/uB
Mzkk8U4KLm/Q3vKXlP/EQDuVCYCV+ZzK0xdhz5Y2KyfGs7yVyHyTqstkg+6Flh0XoPpR33sJEiHF
nN4+hBY1eVTkMIy8t+ULqb5Boo1vJNmAhVJq+X56qm4lRg+SxQV0532BkqQCI5m8DWSp8BS8T0eW
VPozX/Gmb3gAFxI7FqkaVvo1j0oC0l42l6TVGdvUvoXiYz4Sh24YbNK+3i71gPEYfuodR0G1kKO9
O/lWqsUvv6MyxeucFSLGuG1Ezrg0MGYBV/JFModAcwjUAAyRMMFqS2MmLvZX/e/Q09/sAQInI+Wz
UknAAq7wun5iaWKmuDZ/mxEyx82oKG+dJ1rv/5ocuzcsCnrd/+6v80vpAOR6Yb573Hja/QCgjj+F
Wx6svKX0sFNVLjPK21VEI5DU+Rx++gPisVDxSOcfzzxotR/NB1lolQypcwMkZr2fcFC6UhrsZJvw
8L5GokD8AbiZW8KX0Faw9YdNYUgeVyJXOc7tVA4DzBPEp7Cd/IVdR+xgwneTKU8na1WssgvJzM6c
BCfe0wmNgQLhikStFBRF96uGrvUZzYJ9z4sVBR7a0k29es0D1fPEMzCTtHUDJyk0QHSnvDfTVR7K
FsJIbs7EfJsxpCs977g4I0tQW3gclGsNnb6p0lBP3pP8B9XFPphNbCygYAfQAWSfHdd4cpd8YjkD
+zHDKwG7SmZva6LBUd3U+rCgbOpkY7dWJ2yIcGhw9CrLHj6qPfQi5bFlydKxU8RPLbRnLZTtBD0j
+aUsecJJDINc/VMtCKDGrCdcdaEZw7gLhTIWpEug8GiwfdJO37r+liInYhLWOW4B0nxDv74uo4my
uLyPJ5bPNMozZseial0FgoVWro2hHnknAh2hkwGpn2G2WukrKeY9luCI5FEdvJMdL4C6z9nIsoHU
z3ncbpFpOKFFu7sicqqIBDQUWKlW9mWN0OL6uXNB0eb8VwIiJUxC86iZiCuiC48ZfZkSPkBtfn8Z
j2RfYloB1bGGJSEGfCMbagnDE6vjpAyzdWniCGaN7AbHGuKSKzrCHI33bZIPcORX56SjeWGRyS+G
Qe3tDxeeyk5oEY3kEtDdhgSKHxme0z78YKt5rOcDWlkx8MAEX0QPBTRHviSrFSONfT0YeP/kD37/
mHrC3qmn3dSWBdcpEYlyJtSnKhyi9HbiJ8/sDqS2LU1fvy8q9TReZ+y/LIa3Vz14BnnjJ+bKyVF2
YPTOJru8cLTrXkmZqaqFnF15ZxWCeceAB5n/SSZi2OjkEPcJlmimMFPmrButzMd7w4aR7N2I57eI
oYBaGM/it9RdhZX+r6At+tNKV7oP09GkO1CGimMXTLCIUsHJbkEP7YIuZgz/OHxXWV93FegBR6CP
ildzB4RX9IXoDYxcrDM1+BJPJWcc/zEQMzWJhWBGZacM9CWtHG5aNKNy+kvjtbm09UR+LshEdAb8
ZRUMim4nZHJ8JXZzOmhrWq12R05Pw9XqD7se/m0OQr1ZlF1Qu+z7MXPrWujuSVJ6qrTswFZrkHG0
2WHS5zq3coFT9H2B4CRQNKtusHaHjips9Yrh06ZMbvdLuA13rAZBh0KroMq/EuSSss9TSuYqTEWW
nWt6HT/HxDHP57Pz0Ijd+TqNoaJvZ3pkzjdm3pr5fqR9Re2tAD9wdXED0EQUhcM6R1ct6Tg5FfBE
zTrQXIe9C6j/O/PCLRvJzglkaX6Bl5UO9yLSBa20KYwKfNuN9u4aNH2UGPbANlgOBb44CLZhMi2e
b+77pzs4LRS8H2ewjhgKZQxzQzonqrRSYR4MkWBWosxBmyoS2dzsJZGoZeFoVRi5WKaElnl9p8OV
3Q631q1I2ZAfzHHa+zR4wxqoyCLlxCS2Fskdk4qsPoy2hO7mip/NJmyCGIpscCLl8pV3S5RYGxk3
iRE/1jP7dTRG3Mfe0lXLnhxQ1xLUgw93IbRlK+or+VwNNVKtApfabW3AvT9XR+fc94+pQU46QPQy
F+JhERESX1JJp+/SDmRxRj/zDA+izLNF16aLDqJQEybmyT9BJpPuAqmbQZZWHU6F91Vdixiaeany
zUX9ZqzSVU95rWq8zH7yEQLzVv9/B0bTHzm2V5tZbiCzoyQ6RM2+vtQ4ueFovXIfFoe8kkkAR8h/
KV+jq9VlyClocHsawUTJDX8D1t8cA4TThdpQqKrrM9LFESf97LVZ16q+d3HiVxd5PhUBqn2W5Zpf
kdYZmD+Ms10P5mhi1SKF6HiqM+i44m6S1bNzy8T6jHYaRRpI7lI6g67CwWrJ1KLT7cLs3K+Bem8t
9bVN9qFvpDiAwkBFD5LYoMHCWyggh8ur+Kg9aBPLHo/lmxlxDUzeHVk8NJ/C9LdMvIts+c8Ym+JF
FMjuJqs+WTmMO7akhRq7ZTFOfRgU1OZRt8kTxusmdMvIImcL454Ckpli4uKi+n/v8bK3stCFWWbw
Pj7JtGDrPKlhdADosYneG4N9C7aRjSvNRIHzDp4zpM7mgpmKWmNj7AudGon1U3ftcKJobZBnGmyb
6Wv4sWYiiwnbEuCgDulbLcPAQvpYCHyfMF3xYiDICyk+fayAa6WaWcqYzjYx56FAOQzgV7m+f2O8
fWzRTtSmfb4LPZzNWK0P2huE1rurc3yfnE8WazozWPimErIVs01rvei16d9AvnDlq8OWKm10vIcj
xKL2JpYvK/ZlZQ4nWpAy0jx1Sy1yyFTErLYaMMQZ7XCZqG7av0qJtN1GXApCjc9qyXuu/IBkmw/D
fPoKDSq7tYuuKj2RW627ORtHj4YOHvAbf7gY52dGYx/bdVka3w6yMIqpXJ8jltMnMuhZg+Iaj6eu
tgKCB5VbO8FRh+pwc6H2gT1K/ZTPNSOt+MF12ojNOgsLzrEOGTQoZLEwVx8azmWP1jrCDDyTBjMj
R01VwFHZsOLpjBo07cdxxR1LkTCLGMTuINnsxqKdVXQMNY21JFUM9WlJQOvFbr9r4p2Bb5g0gh5x
Or3RtrWfpE2cvEddRqptu0s+303+6FdOGTvSOEa94XTZ0GGbG3DbT+CRggIlnJlFN2GvzuNXrskW
IAmIylwVq4E5zQ98KR02YJIv1nL8uzP0ojltGQzQD/vIgS5d14+UDmLuysWviWIzUe5DlnHF+Oys
LywHDNAkhKpenxdz4070BbO5WaAP4K1isagcGPPidzzwWaHVayX4R0q64ryAyH8nJPtF/Jdlu5OA
6YJ9IIiVyAR9lH66V0GfTX73I8GM9aj25r1sGOS8SvlbTWh+yhuWz7dOFMJB7XsIwH/TdhqXT4el
4hrG+/3Aon+utOXLksmbgZ8vdxEunshJyl80/IEd4X/Th8baWTJHhx0UZ648ADPyyE2SdsrqzSoN
QPhoig9aaDvBOdXXwZNEyx+cVI6pf6tYylqQo+N68XP7tRxLfsMTYsTU88sTNC8Z+8z/20Is1IFP
kjHLRrAUT4djlazqvXZHWrag6CI5cL49r94Fr2KLJVYWBdCyHWtlckIYERHFIEsUEuGI+EhT+i89
wMDmkRLD8HN3DkWS4775GtMf2QFiUWt/T8E5JST9+xzHUOftjOtPwg4OCNNn8lh2V3S4/sBzC5nQ
Z+AR483Fmz9Q0KbeqME0DMB641DjwqIwQFc5O14yeZNsqNBOcmvLXLgET1UHJpwYyE8S7vdqsEu/
KrKpMuaWXd0CzB5t3BYdSqm/DxPM0Xn714SsurGDWDe1pmfEGSQXzjRugW1vbVVwmv8/bB2ysmp3
7WavI0Tjlod6ARJExIpVbufifsPVEaNGGoDo2qQXdhqf/UAryJpPiyYEGS4aLrnlgtrsgwoWPuWF
WRuh6E9XpOTZeiujAOrXly4Q2iUv2X+9gfQPdACy8C5DojgU7JAcc8rYAmeS2aM1f/bajN07rACZ
CTgVw0ZSLUgRLcanIjls2HcGUuboEf1A3EsHyzNUT3Bvv2rU8nGFqDh7RF0yt0j0HpgKthuGZqdb
XHAYcFJ5rrJW9L1cIJjA0q33hqfDn2Mtp/Nto4la28W/QP3ad7awu4mVezinl3G+iodWwtYRc/9Q
U/JQrKZgSRezM3JrsmQKhjckYkVKfEZ5cnbHsg5hnBbe1BFYgjd/+sqWSAV5f+8413e8c/ZtLMj8
0M/KPwfRud+TgQ/Tz1DAf5J8g4K3wtKiDD2XVjPxQVCy1XvUw66iSXHtUV73quMkWni9gipf0ORK
rAA3tx+PbYbYK2A7xpjob+kbhbmvGLk3LVRlxCWluhgNN6d9DfVBXu0XSXOmZ3KbnzsIWaHT78DP
kj0OFkXgEsyrm7uY/qedF7xFOdh9oh+zaiNsgMq6qiuzUdjSsYpTMR6hCnKPyXej2c5L3GjKcGHl
5khXUDqoZUK/ciD9I93wzmWAwIxNhpvpdnwL8ESOFt7GBWmjnt59fCx2qDzzqS8px0CnmG29dWtJ
W5wmtF+zUnurdHP1lGolaI7zocCk+vHtT/YHr2MPbZLGo9Oh9Z2jEFm7vvD3LRJGLLuYI1r6Gf4Q
4qkK4yRnTVtGOn9DkeXwlAt68imWimO3AP9It7dwAj80LOP7w5/4dvyFaBE/77Rdjom8Jb6Zy5Hp
q1G4mH4zUEItUz7/PNpqer33vf1fIETyMY9mtEI5AmrX10zaZBUSsrb3vgfh8HDRwPRsNvzNKtg5
uuviYP3kS2y2DVfMpdKFi2QMpkpnbjNrg6F28pqUcOyX/5hGQ7/03RzYLHd8A5N9lU4/XRWjB4qT
qwIa+yii5aCTCGxHBM0XUEhrfB5qzvr/D0kzyYOXEuA1FV5zqVrzdlOb2b96q54G7eW2UcX3E5MY
skdgRBVVX/d1NuYC/7buycTQ0w8dKEAoWwOIEXorAeFjh+KSDha372dY3wfFs+OKE3NFsH+WBGT5
eVYtrPH2/9GsE59QrhOM0tiZQHSadGFzeCh0xp55N/f1AA/J2h8FlSnl00iOAHBCBpsewcDTFv37
QXdI8+awD664SwO8QrrzBC42AiN2h5J08gZD/pct3lJlOD+Q2kVvtD1q+8bcIO/+Yy+1sN1KL4fr
/BXIVGjR9YwJ/2YJatQm8tpUPnipS1KAh75SR16iTYZkOR5insnrlC8ZSQLh079DWCHl4badRNIG
4fLMwKWKO/oqEZBFmJktxfVZu7iEsfk3suLm6GMyBv2SdOg1X/LlScg6aQnrS4MuyqSbpD8mrZc4
DEPv2H/ltQcid3CBJzvvZ3+jLS2PuWzfeE18yurIwWPrJ0/yBfBJe+2OSHmtzHwvgn9ESGG79z0v
YkpD97lV5oIr9AQiWX8AY2VhYkMGVbaa8TaCm9wvdcLo6fIMvz+MZQv5pwagc/tgzUrJsvNi2Kvw
VFd3vyHygUoM0KON/loOoCV8a9NY7uitsNUmm+/zYCngmgaCn5V9gxypg6FFw1TkAfo0sFXKJIIe
b/Kpq6wOC5mR9iGKnSjQi56NXrkwDJgVQZcAn44TWthSbH7PBEBHfIImGx1bGZDwD1cukgoX6Yl6
1ydQ55/cSfsVAWgeMO0j4KkqfGz8qwdmYlW1HlnoO6k+nJYfBuAR72K4d9R9QGSpv3HzrOhfHMT3
BaGJ1z6EbxRnGeAyHvttYdh1fUNy8lzvAGkIvEhh1NIqxEJbfRkTNsOtys9mb9S9F4gldZgVWG8b
Lm5w1qGsG1arx4llUh0HnJ5XGkY8i874aYL/dfFWicQYn7QTIQ/x+C/9vgR3AFwQrUslIfck9ODi
QhNCoSvGK1w4UTUMT4fIJ5nOT6nlquprW8LTo0GmHUD8kiLGGAzsBDeLB9k2etXvKgbWqRv9l0uZ
Ec3GV5Z9tmeAq7gRK2UiDwvwNo6lmqQNBI9+OuBRmohGP4aDPlcOVZzmdH3xRWOQUTLDdsS4cL7+
zjue/z+eYDMLKmCwcU8dpOLspAIT47cq96T0X1KC1bZfE/LwUGqsX/w0AW5vQ9FuXzEowZK3ZXQj
OrLOA1O25IKInV4nV1l7XnSxQgMSD8xkQbfImtEzjA62wc4NJzQblQWPxjl6dWt92SbmIUZlyvXK
IOVIvrCVP4OijXGn3pXqam4Ix/s8sDTRD+OebOT3ZKVX59mPV+mlFH3QUahSng8keXwfwoJwBz0T
SgFKTa+uo5BPT8eW7VmxsTxTcyLaUqj5hJjAQT6qX5+MEdw+/sbpzfX2uiywaZZQL2RDWNvrMI9y
AiHeNX2SOuOPTmql4p6snAyO4KFfAg7e7xJJMG9fl77gBtFQfaF6CsbZ8L+sMiiDPkLAgMaOv4FP
k0m3lEm681h8roZUEvjIp0IKi1TVg82g+JOCJMNry7sfggDa5eP2lz2pD8U0IA6DYxi1nW0cCBRu
myiAyvI8lpgdS6o6ZaJDNnf8rca5IXEr9bvewjBfPbQBUnP64/WzoGFtdZ/rK1o1IxBgTcYHyKSV
BJNe47hA7svaw+DYGr0Dxeh8Ux1GYZUkNZUPL2eZw74yLJBQd37jeZ49kIgvmPBFoUbUqWYDUEws
i0+Ye8p78t+OMKkQnegbhPngtgEOvIwXEr9eoNaI6jSCsqpoahFfzQJujr8CdETSn2wBePy8Mtep
5YC14zbgQ3bt4CqP7pHRF/0UOSB4jpLzDq2BZyxBsL1gBW+YQJszAHqpJFp1Dupfb8gJNpJvEgaA
90lAyZ+Pz40SaMtJna/O8YL76+Undx1/acxMWYPdqCxQXKYWRTbii2NWY8pQ4D+TF065pMjLYFL3
/56/nxjymihG60weNQ4/2oxqSnuOrTxiCxQ9YcC28quKpmutEne4pxKKB+hl5+Q9Ba+dUucsJ6Oq
ccfZOQ/U9Z17xykyBZDIL44RvyXvlvtM+NT7gvMmaCVkf7bYgGSAzy+BS+U0QGv44UPiEGXF5bg9
S0JRpLTvSpOLb85iRG7rS1bpTBE7nPCjG/EO27L0COXM+sV54CxibIwjWAdmPVPjL+Wa5FYssryT
6seiaKMEv+rXc2OiFE9k47ggvYZbsyNz/1hf+j5+NRVArcoLGn/mkUuS2e3O01bW9zc2GeXPrK1S
ity3eI/8cqScWoznY5851d7Mh4X6Pi2ZrV93Kig1oTjpu2/qaCFz/x3zSoF5pTj9Ftz6KHhscEpc
w2mav6DNhu+NyQvPnKIwj28WlNB8lnFaihTwzXYFddd6+G1D95bh1UGlWC15aAifrn/SIrZZaubT
2yBTnbZL7Vag1fEDpoHebTjcdqgZNJCXdjNPuIFI6gA9L4dOd1GFidBsKtIzdB0b70rwr9VjXWf/
8kms6KVa9Vxi1F8wGvSSbzXv6eV0AI3KaYHTGUx8th1wjvPoD1HnVZGhyJWkcKwaOq4EtDKVBVFt
qa8NHFMccC1+YnPEnE7zvT9m4z8lRS1kJKHiZGDW0aNH7LPsmTrGbLxukXX/83+yYfRq2K3QPgQP
7uz35GsTouVnHUWSgXfmgI3EalTCG1sLp8cpxk1H/kBkIE2MTCsvbl/zoy72yhAS3V4B/79QJ28k
wNc6okW35pIWYRRGFr5UyMmOcAjptISH/23hwXJTsxYvXOih6BXH0tUTd1TgpDUkaXqVA+TVVzhT
oiryWMegt/BnebUfge52wfo807UQuNssXnzbMTwZ/rf5a2TOUvR/ZrAXczK2BO2YVTjlf0kaYUgK
DExhDATz0IMHhO3H7mUyfFUcp89saxBe19ERhvniS2lMmCqqbp8w58tOUJflfSsKsaD2Efv3mgJD
Uh0QtxFzE7hS6XiCg0IntchNZg6ymNakJA9zb+5EXv5d1LG3C9YL9vXm2fjTk1E+utlz+HadU4bC
b07S/SLbA1G/Phs06clJHxjUaHwK+4VDFq/3Rjm82lfAjzYntTbFkgDCgmUMVNdaufHqCx/FAxOJ
ERy0PTsymqsl1YaownzigafREyoyrJcz+pcCFVlenWeqRCXvXBoN3DWQmSj8CL893eIvxJdjtyep
iR13GY1N2MH3mQG4RaEOvAeKPVvx015e14PlUWIylDSdD8mHNxjVNG8XZLd8y3SnyUqG2j6YYQxy
knAQ1R23/TtIY5zjHmypp5ikN/360H/yPPWUOwkopw40dhH7mn47XAGh9kk6iqoNTyKR48W/6nvY
kYyq6x4gvALb/rUrgx8+lovUg7/pS3AZb0NKQOQbhtgrw1Q5GYaT/IFbQK3KRedc4NaYqzeqEdqy
UEZw/bTZDBNQrhf1GCnZfEbl6y+6Bw+VZLxWetM4WpZKwtD+qpnjOQptzsNZqQsgzH/GdMUOR0DG
DFwnMPnTJUNurnx7dZZqWzL2vHpIPP3D12x388MPHPWhOYq2g3/RD/6lFD/8TjgaxiHni7iO2i18
e0RWEdSKPur/qoq72naYG4RXHEH1dANAp7n2BGxYTxRQuk5pkjNF/fgpJMlJC5hpf5CtvLjAOfMk
9CyCeTHRs0h3HIIWqGQylwjz1GL3R0KXkyv39YbwA0ClXL1nDG59afBUGYfWcC+5S6N4w9NOAh0z
LyKsJgzWK+pA1cNaIq+4BC0aqeIpafmGR/LxJpleKb/AcO1y+cjHbK7EEpopOUXVPBPHXRNRfAai
2eu7rt/Jyhmprg4fihit3IykfnFFD04cX79mPPISoQ1RV/mKTHwMId67pl5mIovw8ydd+6RT1qBy
KXb/kRVYyBMyNgf3WsxbLKGtuZaTx52KWzB05w2g01xP1XqpfzE0C0apN9T3bq1XE98fePYswY8y
PE3fUeXAJ8hmUdOLybXex9dvwSRBIC4oWFHQOHfwGeBQ735XTDOAycMxuWBH7pTMRdJhKmvyhbjv
sqc1eHtIIyqTY0/Ql4HnxEJk9sQeWHxrBZk7uh2iy5vXPgAb6Tu1R7UhCSlPqXF7ri+lkwoQ2IAf
5trV0DJyvkDRk20apA5HcDhrEVWseffZ+3qmvlwnepCaMOJRj2Yyh+HCjqnkjMsOzeeIjvB5M1+u
c8G/gWu9u8c8S1p+gil7SgRoK60Pa5SSpZHiRqRmxTVt3/NZUw2TCuYJDZzwujEnfcWT/AySMHHD
9e3fE5VB8VJ0P61JtUzU/Uwah+bSEcbGC40vq+XPBivjyl+UWDe90OjCv/yh8vSEgLduvM8iSNiL
MgVjDWxhTyU3fckfJJ7biq2ISiMJF/pVikTPOPkK7Z+R9w5Jx0nVBS+BojCSwvc8CieiXpgN/zbf
Did9blkuM4jjvirQQktX8OLFCRHE0ILKFpRr2k6Vfl55LPmFlZwNol0SxSw3nA6vPTegj1IybF6V
zKyLugV6d3starUZUNEh+p0fsA2G1esk2ocEqK20m06Km0s1REtxE9FIYMVlh19gsrZUJQafNYW3
ao4qdi+buAS7KbCKrZYO1AohU3oLXVPDXp5NbHgQZIMnaYipJqkbIUn5udMpmOK7bc/g++tdN+bd
MskrVEEWCza1aTJhj3U9Ulu53b4SsSC6eYkQKLr1dEDX9cZsAAtBSKp2QyQdfByzpdfb3tV2jULc
z+zLQGnbJexFibMNxCNHvWR9Jg9oIuZTYR8JG/roe1k6pHttAMDATJ5pGhQpH652kHF3ZEp0JOFw
LsCylVv8EkciLH/6DjMNF1X4/YCWCpOWr3BifZsmkz34ntnsjxXJVrd8Yl14EVnnbjv/ewI6nIia
bzg27/qT7K+M8dtN4B1/0XYBlFT7nYhpeZlVZHNYYd+QJXefFzIBbyhn0aR4YT5gnBFT1yLYCGLj
vNzfJ5GAKJl1XcVnq76US9T0o0LgeMsGe/0q1J0lK/TXN/uR53VXnOhKx2Cp0R4APmC2xOGOvvRz
cp+S6UJuKi+mt8/3hytNrKGgUIMcZCCtAgmvg4rQYHqn+GYOseSA2xbjmuTKDapkNP0JuMFnd+8u
w0FatXEwduK/ScDZ68zhk/IjRxq2RvC8llpvPhpbw7snG6rwGVxQwqjM2o3ekAK1HufGcqmJ1tGQ
Mwgt0zBXaDDA3SETeRriT6ACu2pxgnuOHdl/PBjMBV8jegkW59en0FXaiLyvuWbp4lf+iGrcwJFc
3OQsHtHgLavXSUrFl/tTvDwGuPKGVqOMsD0/8UR2E0dX7lSLqypaZJxGUD14cQLPUeRTCwz1cDSv
p6tRPJgeTAVKeDDBtqsVNI7gAmaYf6gyLGvVXWjBi6NYE3G2Iw6YLzBjnvx7X6RmVyvaCk/fXtxp
Wfvc+41FY2dA3BeFAHGijx/ZRdy3cz/K2qjjEryzB4E2vwKJ5h/3sWkcCHP3XB/AyQW9vW/l4/Bu
WTTkDY0hNE9W8C6POodI62RJqyLMnGuHogEYYrHHlEiczjJEuZhXoGL0WWgVyt1IpsaCH2tv7ES9
zdo6Cj7TkWrdee/GiWMZR0VFFPeKjqJ9bhdw+0HIekYvJOYyk+fga4xNjkahdAGP0kXPQT+5d/kY
lSDD0eSKFOTnay7vN1lZlsRYLmYtoU1JwruwWgIJJZWrbPdBjX8r+ASpSqDzswwgwxglXAY9b4hz
FzHMs24ydNKZFDkY7woYYjYTbxvDOoExYAPBo/fuih/pKOnKPdBhFosNCW60wt3Rx36R4Qjm+L0Z
RApCwg0JWOuIrzADNLE+sVBjbJszv+wergZHGBY+pktMm4Tcxj35MAoDMfG3siWbZ2ikVveV7cQw
Wdm66bm9B6LFd6SBMUrn7HiTnAVnKcJXszXbUUI0AOziCd8Pc3KosNpuRTT9Du9sV5Jf5VE+N6pF
rAdbhoZ+ZvIFfzLFD+OTA7mv4QoSwZMsEjT09Q/FW1RKoZ1Ul+mQB0V/RuP+eH1hfZTU6DNNn+D3
U0l6z2SbAM3nuKDq4wibqMzQOM/s3DVtmhv8oB1NB5cmxtxWj1wcCUrA1Q3r26eFIpwl5IRSXO3r
OErvOyhkyrIcbfsvnMkAtOciE+xmlJ14+FDtdyJOMHeIKwwb96eoSfUe2l/VIUX5BBx673UpjDRF
bZ2TJPAlcX0nzUdQ13lMOf5bymIi4GErpddLC0iJXkPdUV+ZtaZdzAXdwwrWIEDdihrvUgpdrt4a
O/JbRXw7M7iwmvc8xEkR6tmMa1RKns6yVflTjVjEJc5ZUSZSrUWWEKlvlms+sIXoHfxp8hE23ydB
3cb0KKtR5XpdZBDHWk7YLE8pncWAEzRF8irifysMu++HhgdoN9r6kaW14dY0iSM/FgZ14mTeRmJS
0t9qdHfiYKpm1ETHHfAMM0ZqFhCDmvWJOnAS9icFQvRSO2zPtoSO2u70P/GXZ1JrZ+JDkvTG2qr3
o3xdb8o0amul8QFLTMlMBMqQ2dEHlScyVeBFEWRWDGO14Q38mG5dVFkCLH/fE+6/56O/tgErpytH
Y7iHIXueKaqZPBUa5SRmej6E+hyh4KCJ4PzsDY6MTPiycpobUf0haBcLviUCSGmZAUe9InDbNm1M
Y57rYj52vQZebfXKB6lPkolHP6RW1D42wO+RwzG1g++pXLXR7UjOaFSieTHPapqBPjjnP6YJr6UJ
LZ8zFJxiWD+MqoFyj9fO0Gwpt+lenFU2hCwDn9p9VAFSBp0P3Pc0FpjVj88BAmNYPsxPcxshD5Ly
SQGEpG7oeqhIO/zCuN/yHI3yYngPM8lQyDwNPmduUwnJfTmeuax4WfmhhAXQ330LOS+iChd4U3XO
70j0wVT4/BYJP1hfSdQOsWFuYtCrzhTYnHhjkpyA1KQimsmJ9HKTiB/yfK7XVVZep0yxiDG6F9d8
M+RYKy/qMFyX8db3P4P3UlbNmeOSPpIgzf+pr+RVKWEcW5wKOpOafj7DKERqOXOGVRbOGjjJ/m1r
2kyEJhq8TJrgNxE7llDjrg3/D7ajcfAAt8koBoiITDa7nrR6O7tNNNpe2qJ8HSCufMBK9H1MbrZd
1g/pH/lsO7WX7mz38z+rRXVNP1XAJm1YGkSEREaZ86KIQWoin8ZjwENHJEdT8LxCHhu2PnHXeXXR
yZjIXHOBXFqCtXAYJquTvWErhODaLG29ZJEj/uBDoXqrzIY6b7+fjEglglKMO+dBc2qOLjiHzVpM
s/wK69hoX3gxA+K3ql4PmLhckYRm/zqehrmtDsSIG2is2J8XxXlna8AY7iemRu1DdmEusotlzJcK
vwVmvHtZwOUxjEFrUKl7mMmEt2yOEWIgRs6I7iWYAFkYxpv/HZI5yFyFfHRDU8DpWbITcIzjm5Yf
sqFTfJNdQmqdr4EWgUnyHXRqxSgM6buUdDxmX6sDMyPBD+oszJn27/F7pP+3+aDeF2hjvTyIeqnh
wFteBS5bpRx/n+HN5SYY0Zvi39Az2/AsuWT62PPvcc3CjtAvpMiTFFR7gSa/zv7Hgpcv8kih0kRC
eWeDAX7BWfrRll4RQGLurMAxMjPJnMy1tTgu2T/doenZMFe4Z7iYAqk+P6s0MX5no1IW2HbBypCb
kAGSdbE96+Xs2C4Sg8daOM/055IQYLijS4zwwkbfyPWAGrbCX7T5KXrIlzmnY4ORuxtWnFnabMkO
q+doZmIZJgwLJeT6lu+HmbdyCdEhGhBJ7eJlCk1WQ08Gz0pGh+TwEk8K27Rw6v6N+10ZWKtylio1
acfs+uDB33upYB9S0UJ5ETKVkc1xzSJYJnHIEQff+AjavVUWXM8g7hvIDpjFhP3sIWYA7vnOwk+6
iYmpjjF93OxQLRSR43Nk1y8E1ouUR+hV6Rr4eoF9x0knPzYr3pfo8u+NbTAmvmnhFXgAEsBd6R5Q
9mOG8jwJMGwXUNpGrYos5gO4LsefxMMx6J+yoHZ4MI0qRfa06At2xBVCCRFJbHCSnwCYnz9NEJwk
+uXsKJaapnA62D7U2wm+HI4Sf1skYJHSx6eizPEMb1pIeZIayF4N5e4zQu5TgHK7qrn3y3kcEa7U
eM6qjLICKSs1QM+vdH2bmLzs0lkjXiTE3nftpae2jxFfrB8z65IozqHi1sPWeQ+HkQW9YMGlAFBX
2t2kJny77SEIeREnmKORnleZF2bA6wpFimmdjg4DCJ+d3TEkSKiLBTYfRssQ8XMygcM8Pj5eAsWS
cX8rTglV6Ts0HDWCrUpZxl1t/911JtoYC60aytp/GaCAij1biUURPhQSoobOWlU/NmLoOYZQlSDv
NkcFhxo9WrLLNtmjTT+NgSuqDLtHEFqPNOykdLI8FOuf23AlVjQyOcZOiG7MAMRVQ0NS7U853oeV
8BBAyEndtMOfDufxi8BPyFtjLdAxwiY7B/iyejsJLjVLGCUHnr9Xn9XFhvXWb65LTn1zbgCd7liW
hrmi9F3VDOpBihlsxNHvcU50Ak9rrwrTfkt92ffsa1FAHINIzvorjSqghJGZvXui3wNMan1TjP60
+vEYzc4VQNd6Za+1JVdFz/u62iP1yzDV9VoMcxDAWHCeRUBDBugv+QEaikHqs0U6znhRFzRDTXtM
H4wMCNFECIbkGachLwHvZ+t8M9CIB6lkBBOpErD5bciMKw8z+nNWNa4cAZ/xiaqoPHibNq+omRer
Mc3G6E4VdXvR23XtqCQSbqbOho5gqIkxMX3gyGr9mimIGMx+rqgObC7VG3+hBACPFG4YOzWqT0iW
hCm5e4E2KNOjydVqXFuFPT9yP8qpaNY3FLujHTkIrBIC5LJWn36J4eci1IYX9nIfvcUVKL0cSRRX
2kZsdFcQgqe4OK9XplxuVlkQi0crfzWtRrFsmg8m0yCXbCspbMC4F/RgddU10XKEbIjSrZuZblIG
p+3bCYUzbckkPIvYlh/o7GZe4I0Ogd+Xx4BbeNfg9W32mHayQKznKzMuL/n+0+kSyCwojZGtsaBE
EFSBTiJhQ1EiRGVgPApPrszCqiqhf53T/Y/3GOxf3nEAwtWzPREbvNzuIN4W3ITLgLw9tPopSrFQ
vFE0X5WzaCftMwSJDj5v9d21eqK5sSOu4MsXN1Tz3eVTlzPFGGthvf0kz+pCA7mQw8yTwAOCFNKr
1qxVR45wX3LVyR1ONuhStCgVqpkRMps9KqhrC0+xlSbYjiUCx0npN47APDJasSBi/0oqZJR9qIHX
sErucR5tIwOQLlhibjFtetq4qKl6JVv4+z3ku4GzfQfR9But+dD1YMw/TGJp9jeR1ha/T753uGYj
N8+zMVh1oPB26ycWTfrkoK71dHYkXZ01oGeHrYOOuuav6EcKVzHtNVsDSz6m51RTGQv7kGGQWsLx
bRKoiNJ7ZMvXIkGpOhn/1kbcFwUAc1Odke4yEsB/LPZiUdcxFnBqJ3TejbhnE+4rKhOqfZzSdB5M
I/N1zkCPfeTes58tAOVjqyNYw8DsiqjCMZWTWw6L6FwBnCQDJ5ZnzWgQBDPfKRSj/3TgesHW95xI
C/H7js3/9cTBIwCbBPLnoQCqIcyLFbRL0j/8FrOf5or3YQA9h5NXMQTynlLZbKwRNd3sieIForYM
dzF9DYXHELYGqpXX25Z2H7rK4/5OOLElnmFQBqthDIyy6rpOvIBZgox0NGo0CxtjAW02bBVN76sr
fg8nDTHiQhtio4qiiCJ1L58+zeeS2KsKf9bLG9zmHfflvrrs+P0xKHX4SLXPjkUY2n2fqsVu+tUb
WN+GDtZRp0GHV7wHjp0tBwQe+5tlqQiRYiWrHapHM03n5q8a6h2ZuYn8tToa9TRIHeukMlJ5vNc1
jMzm642QYJ/6MPVZDRZ78VlGr0d8vmuyqFFSUcIro4R5yJoA2P6M1zHdaiou3z5RJND+Am8aeItW
MowNaS8s5cAidN/lbNLHhkYeNyF/QNC1GYw9DDOUmkzioCSlIPnR81M3Pl6vowbrd6z/z6OVgJSm
XGXYmYFhexsyYzSMMupKOjMvApXf+DiP6u44y+SY2iHS3bSc6VgMe0eWG/qt0K1XgWxazPyr5plD
3Tgs8mmiyymSGob0SeEilYww+kc74v4WIpu7b6EzQoiGMiI3VotWm43L+xwu/fkbPkXih27wGZb9
tizAAM+C+SfEA1P61niYQyUFT35jeCQMP3APpBfxoxssAABWPhvq6An7mgHXHKn683NPhqx11euh
ovoA1GM6xjBmZHY6XHKlDapAmEdxz0N1cZXuzJ16TiJ4h2sFrCT26ayIlop/ecwbI2Msh1PN+mV9
IUVw9oC+wy64m7YW3jCerRrzyqbe0eVBzHBxTZ0AkKyBf2oMIljQQ1FaM7rrr4bCBZJBMUV+cmZN
dZb5UdF2EZ/988XUEDxtJnHhXkYYYbdOMlI9OFwU/78fKYfpEP4eLlbb2GGd6Vs/T3wtfqAm4zH3
HhxL6ZU4ryZfZzJ5vZKBxY9BBkDP+bg+Tbs/pUjkRIxvDeO1YRfkg5vjKY748mF2oGrS5RK0qLSg
u35PpD33A7iwBlogwZnnIx1GPnZ54hOXabrSvbay1yUuCXFzTRiTr5RANmfePxJHdPljX77NWeZY
FPM41eGjwT/62o8XBeevZeiLBMQRphZhQcMKpMlvscDZiHc3MAAHl4EvlRE0RO9CPL+IjyqshYlc
w9/cfdpuNwiDFKBBYSwglAB+NFh2+efYboUbyXDCT+J6b/CQcED0dWGAh4FXQzKeBTOEsyfdi9Q2
MvNSq04d89ta+uAeUFuqFQ6cisQEWtdoLGzLMaDVcz+KXA4agRSZ82YgJ7mkmfOjK4VAcOn70yK0
8K3UwLkLTKhEzD5v9Yt9KTyCwkiBpIX1KmNgIpNfviJ1YPoVBmANIN5iBfv2D99L6Fn6M4Gu+f+I
ZB9oLnTsBVRM7EpmVjitDsRen/uIwT8hCE0AOikMiEIGLaRZEhT0ax5c47OdyOxofMr0yYFIB/F0
8PMxChy/ZjPfyzEnxyFbHPE1TvHHe8WYvs/VbUvQHW5KgB6Mc9NneBkdu0V8T9YkTthwgZkAb00y
WA1AZnpjQeT+Y4heXYIpT24O8abBtO1WrjMTgeQdgHMdBK8NeAH1lTWUoX3cUEiduf/+q/XCbmzZ
JDHNuQSkxjl8Gy74aGD6wV97dqQGBub3ftZx0YVvtn81JglAaFuIknvTTEXD7w64Wft6CrJTpIgZ
YzMwSpogngeKzXlAy1knw3mCBytLErtnnN8G7fk4pwhbcTy9py0TU2jxLf/74PGThrxn/67FB4T/
0aG2vRwBrBv/Q8O7d5mmbds5DAgTW3w3n5if1WLhKpfTjaMKtjpQjhT9OT0mlpw0xWkIJhTl71UA
dB3kLYEmalvB1ZeUGjyKybSWzhne6Kqbxz2ZDNUToVz6exo4K4iknzXHNvY3qXVj1u04xUN7CcLF
vm1ZBnoq4yrWgKqFNSRoP8qnVmhWOvt2FYtqydFYPezlKtgmCeyT3dAly8a5tUW/F1wAAtgLPebk
NxrWKN//C7Or8vdp1X/YDBrDX70spCsxl6+KV20oEwMjgbDgrXeF1hEjXHMmvqz23yJGN8zmiXs9
CbZB0hVIIF3kVuoGh4CSBNKs00Ey2faRBvbYJrVkIOxs5MaPeFPxSaoHU9+w7L1Y94CBD6UQGWnA
mzUyv7irhuBYPNuSTAn0M9NjEePZu/Ms5lEbxxESg134DZ3Q2kXwGEmsBKWwtf6VLjJED5gl/Vd/
GoNDPZ0ZSU8HNcLwBLgWxHXA5FrWqk6deNy87X02dJyB/7jdsc8KS3JoxYcfQkR8t4xPGx2Wv8RY
CwYp6NjLqDuSLTosoZqQy68bxXnVfOVUHFLarYJZo2ec4dGf8t9DQgieCsRouo0ywedj2qu0cs2L
PMrngD1tmbhKiXCviuC73DIQTOK54R9gCX6TixjxWXZRBBSwcNtHc3N4mmwkPEgIIYQhBxMOP7Sw
e2BTGYi9b4MCoINMDmDhMw7YXJ81RsP7ps+n0Pf+V7rfUjui8kzUWB1sA2pyEH6ovxV2YGq3IPy7
zv/5zGxAq+Lf/PaOx6RsCiAJie7PyMKjbsZzLacrLGSmD5xBPOeQY8oLxORclRQbLHr9+WNUCA19
lPlaem9mjQJo9L21KN6RYdSjl7RusvjcCLkvyeOFK/RfyuHtLRerHh/GpUHLtBd+kB2hNa5YZI0z
zCbdvQlR/JaQzF93vD/USzpUoP5l9CvjTBc4hQnq5ZLVFVRoXiOpTaYX56M3CizK3BPkY2Ze5fYL
klxd33EgsDtWu8PBETBt+nAlxPbiN+WaXeP+n71lY5rQgnceYpSQ8Z+U8naBdU8BO86llgwkWcM+
GAXOU2AJrC51wu+I3J8gHSa2ibzCBQe1WNZvnDAi7aSIJxNPPVo8zKrLAcFLgfWTe3Km3SyJNaHm
nCo52ZylKjvPaBzo2nKyGPgLuFE4e0uHgFk9q9rTY0JE1MTd6vSYK6+CkTbHNPZB4zfKXZzgtpXP
OlTXVf4csK4jHeDXtOoGRX17anEkvP34EwBGF7pUsp7qM3c22UNxUAVtlPuDr5d1ZUiMfd5v+R2V
ss5XiOzAu+IghgnYtzfShIMJLSdrVfdaPP++j3/MM38K5BdmWjk/Qo+Zt831KyUtCJNL1z6NuBrw
ZCCiG6rui22J1D9wxjQ8LSMRG5t3U8ReO7qRbJfTYmkxt7xscUSCuQz07S31xWkIcOCwExsrkA/q
HIPY72n/yRucmqGkJbDPRQXLA6Cv8YyMfuYwUGeGliu0RPkgC7cUUkj3IXUdhh65dkTKFoR+4wjR
NZUDlDGziTZr7L3gDpNdaY9eQCGfkxLiVG/C/OGhHEAEwbAwVlnVV6UP5Y0NRF64/2pjYJLEQRnb
qz/bJ46uIiGg1L3SdIYg/glLpAEZ2aAxz9tcHtdkesoZtAViPGyr0IekpuTYlT9FTnwygvoKT3pa
/Roh79JHT4ycpiyx/1qFlQd6viIeWX4kY7kLcFvWUohMz7Iq+qF4WV243Agg3DFy8keJcDdMbK0p
kDww8HUb2xX6payyduRmeUTJdkiLg7+WK9FZ4iwquhm0CCu3mXiAjfRkcfygPFaE7sY1fywtpoCl
O99tBMQZvjGHHQA/wZvQYeMTVkiQAOofysTmHivGswYyGN3fPuMNXq/YX3VB3kpmT1hzx8Zti72+
grMt2chwRlbFmpGn1UrV4qSFMD1NhSTuy9tGW8ttMylwaZP7kXwDsu6KouVBbf+VcGpqxzWRiJGe
8aq0G+RxLnGSlJU4ZzpwGWPszkZJHxp7S+ogui6k3EjezVpVkp5V/9DPAhIbZQexepfn2uOX1Q4Y
FrAAUkhGoAVpT73Nk+rt5LR5FVdAUuct4mH7n1uIBoijJ8UJEgaZc4ijzcRVQa+4HFOdJ9wItL9V
Q+z6PX28TBYNXPtuCgzntWbgDKRZcL7+uuvfpg+nrPrUy2jXzzaVqTh4+2p5QSkQnDQhjgxx2H31
fuVtQFbFLkKKRpnOA5RhPDIiHMeGlfVAkU3GKVAMXxZr0sLke6lrfdbI+zh697LAvn23Sv+jvEXw
SczOboo4SK5k1Yswri57/x52USIBX7o2sDNStaA/jKcbSLpg+CQdVyKz4LvaNqy1eAJWpZIS0CqA
ot4S7oBIXx78IHQFHxKEHYOHn3GitWuwKAnnI31JbNoETTQ4Wao4A1X5jDiz0lL2pZm8UwuoF111
tZ/WOEfE2xoIGA9y1dPFkyu1OEeyWG9QhDDIlfZM3W4DXZ8aZn1ZGCAsTYUUaC14L2KqyPP6Ef+Z
5X5kHp6kZhtaBevCu0LpivOtqgJco/3p5jDQOjax/FcYAnB25VwN/c4MOjTOauLPNNy1MoDYDRtR
oOiNeIYOt9joNmCgS4F7dqDIAPZhs5kyHglSyHlBXJcghP24r5WN6tdxu16JsrQaby57HVMsC6sR
04PP6cysQsvRbd5bvazY1qSroiPioinqQ1O0/OiO2pniAY8dfmH9kXjYcXHJSPP2+hNBPHfl18Wl
G2RBMjZ/jamPXbj7b6pVu/euAdDxVNZeYdwPuuXJs5YH+P0h86TUQS2dy7BG/BT9ZX1fE/nc37H1
wDO1DCvH57kbYb1gJRGd5f00Wkhj2+camzhl4qGfyRDKZj9KVDryiVfcpc1Ym7lyXQ2e2kCcsQLE
awEtORjaZRnRJWh7MoxM2h9DZgku9J9sbZ9Kd9LxJ4zu390asMGemA7/5PnglMVtzXzE7M4PGkTC
WbRQQudcRiCq3pkMmrqbYsdCBGvYYvQ4vXmAuuD44bgMNmgaVGrI5X5wcF+rxJrKIvQw5q4JRa2G
vqeokx+up2JfvAEyqZT46hP4ozhQlh5ljFhREyAz0ZY5eD0a8wXaMW4aS84Pr3lC3xEiD3AWEaxR
xSHeuP0BhX71NdCm6kgC2yEOWXAuZNJ5n/lDFf4F+b7TPPyj1A7cscwDeb8KxZlOZSc4pOe3qHGQ
4zUkg5nQlVOHeYPLAOQFxMppRVjQ7UdFu/9Mga9geDGYyZGvSfm4sYk6ud91ThI2A9KzZyyLaQny
ZR2ey6hUzp8H5gKtKh2CuFliJDC4cRHxpMeh44rcgGYbF6WOFMrZMu6am+tNZ0iBztHBAIj6SUlH
KhhSd4aJ6CumHJXc6MeKPh3d0R2zxXpRLjldsoJp/Mrx2yqNrMo385arBaLW1dEnFuouRwB7MGhA
73RyV9MJsnS2x2h5BVjITYTtStBRZY0uP3XX3cofiV73V7jamX2M7/i6T9LJQT/uiFZ+afLKO+o4
psIVRJhXWTANp1V9Je824CGGEk9kisMdP0lNluvvjozJfRB33ZFEDnH4sZF+NjtALqj+DhK6qkCn
nptucCgJnXKXzSTgORPr1Ij68y+vAvbNZIkf4h/21MzQlzL1N84VzsDGGL9TXlP+39QvxNq8vXvj
GUIVAl9ydiIaQXQ5j5sd1XFHYomAGAkw14WuTirHvv+tSQRhAk6UuXDw3n3MPLRa6vgU4T2Q5/DF
XGJ43flNduySp4MCZg7WSEuT2fmVsBiglKmFqA9cRfMDCHipMYBi0px+QSaIZv9UcSvfBPeBz7rA
RBs92SFEtWDUahCs+GrBDk99TxK+eoSHJoCX/Z5IDqhsh7TtNqAP+UjZY3WCv3/50+Bz5S4o3o5g
IpcLWAEVPxPYfp0osKGWQO0BTtbWZkmKU08McmJdqLs74+4M0m9oxhnIBkOUA4Bngxp1qcj1SWag
/2edPdbXoEZUVcFOJkEsOqIGSWMKk6dz9L35KlA2mVNwHTseZxasMWDFMNx9avsQzamjiU4rGHQO
cusK3zME9iuU7Goyir19Rxs+1CDpb0+jUk7u7EuSBbmGkneQivey4mNlx/QLLlQfdV+JtDDHY4EV
C1Flb6Og2GnZuTv1wGtYV6ToizAAYGcmHej48SNFySQI43wraJ6z6oLxI8LqxE/klfn8YGueo3lx
Zy3yk8yPE4Men8xxX4zr5y0+ACDVxYlQmNu+xvzCFmmMtvAA56nxJ2o3/jsQMOH+O3F2CXn+isWM
Sd33AxuGKuk9HdHdhWBbP6HkVL0qDLal9iEAOoP2D9waDTqJclQUhxhRh6CqhocHXYwfWAZfuJPl
cbnUQcCHvZix8Rbr66DJjJjJPMGz0sxKbJeMZZUBb5MO5cBXfVP9R/gscjzasLysnd4xt/L9ZmBJ
5Ih97FqnIncnL7CaAqGhYrMcYyN/m4uBq0ZEtpneCotkeoHOvx5NGu+sdetdsnceUb44UpIkj/ZM
SL6hQTsZLWastjEAQ351dgEFmOfeSXtqVZaoVf6I8XIztmdjGiA6jSxu3iiBnPXn34YM1t5XFWQ0
wrsG8v8SX5ieGhnAQ5gD+v+ZG1Oi1euCo5xSUbsZIqW8uTywTS9J4yQJsy6XJXxgWMI9DfJhQ8uX
W4bjzoHU1Mnh3L7W1SdSgZ7ngpu0M/iMMqxZY1zeK6l/pwda/zpF7V1BUJj+nT5zYRas8IFnmACK
ngnHOsRnJutZ3e3/U7rw0kUUzs0fLvIaJPxNc3D4HJVWho4pE29xESV83+HF6qeh7Y5SDZAJ3Nay
5a5AyVG0alY5xP9gtgs2ShFKImf4h1iNkJqierZ3MMeeK7cS/2k0gU6joyzL605Zt2vi4qCVl2mr
b6P0KWuhPSvW4kSEotkf64hGmyqTJ7NL8PNdxgvObfLc/Ue+U7MdHsbtCOJtzskr5/uVbUgYn0HQ
FtVEwspkc7hij6w3aEloRdISPAKLccYXhP3citnRQXqlGwd+EOJZtehU/LWdY2nNYqtEB0tDZJ23
/yaLQkP6e97FHxrUcpn+smcKJ2yeoE7iLy5amcMHQoYJ0tMXRcN4hiKfmkCGou2zBto7O0Wsuhju
5+e/dlwgNHKBhgDmNXpSHYivCAsyCmFv2WAuRu8vRSzorbct3uQAyl76eBtZpKZsx68vo6fqXDwr
af+p9HZo0e3/IVq+n3XyOoEK80aem+QCmt0dvMQE8RBd3O6A1i0pKpNoOIp9p5Ilv+yo0RnDX8Ve
KxZhSChHp9MSTbLSZQ/pLSBlu4ygrYORkGG5P+amwaGYzZE0Kscr2ClEjMt7bXRoudH0+AFKVNOX
2D6zRtCajTCQXP3gYnhp0ALVzC4IFuS4r+NjdZc3M0BYKO+NUycl1ZJiWqM5clBwfSJbkZnS0SfG
XHvuC4r1s1jKKhEnVRyJyTtNAtnv1EmLIFjBCzeh/zfF2kgvro2Bo2jBeFegEIL8WM2PngCnY5f9
2pr8C7PcF1T0THp6+jo0ZfB4xPpexmslzqC3jJU/mZiEZ95m9nnf3He01wnkXF1Ud39ZpAjd2Pts
+tqA6xa1zS3cKzwcTH+Z2d03ofl1bFiVOffr2EFFQBhGhliRIJndhxqo51BHaezHwRtzqRwfQ3Ep
BTCq6p//kEbK5GLDc6pNtO1x023BnFlLnChba5Hb6g5oE7NWVVzWNTcfQMvE9/42tRtXJesCIsra
BVjAJcH93LaveV7FsDmDQh+8WSD1IvwTdh0Tgla3j/0QOy1UWVWutXKJrLYlwdfb/mWyG4GCvwNy
dnBvVdfKpzy5ARWOs8EnxY1V4T4l2/VTrSMio/NS5vX2mDNy6nnIQnaQXVlC+kz2kEE1up9BK85H
lXnpv1CdxJYSEHTwXRNrGFJb8X8S2mdrotxKgkqVxQc/U7+4pwZYtjv6qTDDVS9TRaBcSYFsLERY
Gp5nz3drFWPFrYnwirDXcEyLI2YQfWy5fX0UburpRkZbxvfATl3KXKDOCUcsQz00f3a80FgHW35W
DkIBYdeuahLhdCWgK3wktg8cYSu4Ih7J0J1fYHxupITvVvpc3RkxakmBtZg2PT9BIxr7VaFFWDcV
TaqZkv0oOqzKHPpA5Nu1Bfkj9YZyCo9YNlVmkQCUysKTBhIvnDPh5DY++ZtSpnMqv29iFu/PWKn/
ipqvay43PXR0uVGOJ3AFkOO4qDLb8f4zHAmcIeki3aBKXiLne8V7s0XgoWBmlsU3FqBO+nPODDDD
sZzkHtuJ8Y+AG1oS57xouvPQzjvyqFeicaSNQqmLHHajfB1Vj2U43CanQ+HdqB6dIfa1xHpNEKw0
S3b4XCd3VFUaHau2khzdTNd/N/lrOr0+i0RrxJi0dk9BWm3f+beY8qife3aKASceH7n6pszJ8wHS
TSoW6QgakLelQnVROAi4gdaasiPJQpfOM1pK6YVNznasK9JNooALOXv7Tnfz4d5P7LrCK+j0naHh
I53bxzrNp8Yz32AlqcChQCjSx/MS8JewSXR6YcHcPcynSyOD7GvG5QpLvxIjQXox+o1uzBTfjWWm
DE/DTrnUEZj3/IW/F/XvzWN4/wX/XcwRPT4WYobBTtMhVuiYE0ekuqN+QNMF83OlszLTRPKW2fHh
AkG6EWGnVaIS7hvaAPGB9ePu5cxFg4ylQIB1AAyHtPQdxZnH1lcbIXPDYrl3N7OrswARCFNdbqWW
dcRwrx03+ytJLLOqQv7wlOC2P1Pzbkidh+2tZuhG5j/QOOrUsk3bQMubDo6e5fhuBZB9HqBZjiZE
jZJK03w8vpzh5kG3U9uIqYHiEtGS5b/QealrJkmXDhhf1tDB4BNfk9OaoJmbv/CgBo6d0Slx+l70
NTdnrjr1o4qFIDFXh5yETqKm1PfdMTm8kb+OoGLN7oKLybc7RSEXUV6dbtHwQLw9jgBjt+BNgMVC
oLl6gL34rLr+M1TeWBWMKcK4+FphoZ9Zq8rQ/DkklQ8JO5GmQa7mOehCCqaj6ecFh0jC3VqtRxWx
Zb5eoPi61UlTPZvwGdxTXQLs8xLzZ60lGn/51yBZiIXvY/Z35I/fh4JAgNfgIsmkDuofSOhbpcII
MZFr90T+z9K+o4rFZlKDqTyNfFxWAQoz4tdumCwbbIxVkTIfc3T0jUQ66MdH53i6ghCfxRbonTgx
EtG2P+VDLbFpWckPLdFKzwMX5i/VTIN0xlO/Kme+7W9NshzotnSnNH90VNL9TjeIPSH+naZ5Sc81
6gTiCqaaX7pEu6wCqBAVNEoV+BJCG5HD/Ym5mcN40p+lBo+fNIBazTMJgW5iG7TqtCp7zX8HzsFf
cGjbpKMfSRJtM4Gftzl09yuaQnQ7XgSOg30tz0bpgA0dfIO/IgiuEir8NFLX3ML8/OlKyoLBHfcB
GTS4gzfrduQQ5yK7TmMGTEeGRtCQ2zQiDenQ+fX+5dh6MDBcrWCTFWmkcNh3Kgekjhb5nWPs7CHg
es1pyeOwjxkjqIHSVgLSzQsMfD7Zli5NWMCEXBALsU4OHb8Fpf62y+lMPbKZgt9mKQPuhIJ5/W4K
L6e49TOa+rMrCg59uHLpBttS/7N/512xEsoKFRdryYdZIEyjHrUyVqMZ4cPifUm3dRmmlixclGgG
pRBKphBKw5ArTMsgDpK2TLdjAWM+Hf3l810fXCGjiqP4oSYLfz49un1NxdtHY3tWmrCWCjI37YJl
hSU6y6XbB9sX3iLEat4wiklJeiDSh5R6X4Fc16r0QEUAJWEZN4Oyx/oNDndzuOgIBmkuZd7EdSGv
S/lH+EDVt34oCB4/P6ZtX2Tggzh5XvDs52gXOxTySJPgPPl0WusDzuThtHvIoNCGPltQoSQjVpXe
hqV0xDX+FbN2nIkcC90QExWtSwne0lrdtbxjXVdrXQjDQ/amUmZjqc26ZDh2iSB3+S+pzvW2T/BI
4g4XlCkW2rdPXmSJ8lMuCL4DUdRniCztOLvmmlz1xtJFitfiSGngbgw7+DaGbawtOdmrS0v5GJXo
bE60DvNNAAoRkjONMyF/kaIhgr6PvIKChhvw+OMipNQYUFmU0mkjzeQironhiY/uiiZBFSy1uEhZ
VIhZGDENKj10Vbnkg55zl3c2rJQJbiE4qLnL/bcmE0wz+5e3Q9TagsRV4GXcN2fPVQP+DKVs+89+
CdkYyXEn376Z3/zPbhZ/DA0AWb5VsavNTWRHF7YkP6lt7UAgvkdnl0QiYS5zzVuY7z+iX/qvxjOw
7CjtQ9pfAOrdG3Hm2JY0YNcG3Y7PRR3OU+PuF1B81EUJ48uXzzLEn8sS5UPZPp1hXl0COejLZrQ1
kvpzyjF8wdg/hRA5A51yJPLAGsXUqmuePSLjC8c5Cesg4ASvvCCt3XQywjv429+n0/8DoNLHJoah
devsGrO+e8HXCitcoEMeUn1T0i2c/TyYkIENJQFtg0gyYjnm+wS4tXq7jEgP18hVxmHjVE4YWDf8
HFgdyiyk7YQWFGEjRe8/779kjLLIdG1ZxVvfvQ2dVli0JtgjKDsgdwr2Cy0qzfVmbVlqLN9iEdTf
OYuzKgeMeOJrl2LmDQ4dQ1BbTfcUfm3PtLC96obNeWGvsms6gqFqa7VWxkIaLjDcothq51LuZAzx
G7goOMuNo9IqW0QElUSJndMB2zWxq5pIk385x1cvBa488Zbu9UNmkHNW5cR/SZkXp0BKjMmYNdZH
YYRvtrY+yLRos8PJwifGfm4iXcLYLWZESSlrBibaP4ijtlBadM1WvQMyb1gtaU538dE7PTCSYPtE
GR0FBmz2XpWLnZD62y8mi4g4IgwylOxl0cDKYoZfiMm/HYiMGcQaC15+SfEW2wInU3q9kaWq3OiQ
eUedLgthPA7Hx7xbVoVLLQy+Pi0k4/3deKEYKitHswzOwhKWglKhS9O6wWXK74QMisxqrq4nWKJV
pxLe513EWRoC52YJAuhLhvX5ostMjug1TqN12CM2ip0t+7lMKe7PA/nDdojXq3IAjapUnooBRPGj
nIEh10kPLR6msALrRNxAqvnwrpxkWgPvvac1wtIWzoW/0jpEgl/S4LbYF0Bd/LRk2lRrnSQFvTQK
o2wA9/cEC7xlUvotYrme7i0e0l9ah0fvANU9O1eutbEDgvYLVM7OPSdlJPggPCcxWRv8VMJ62kNn
+yNCj8liriH2wRXsrkURYo8nMrdcV+d0gQDTLFNUzqHBwn4IZJGkN/2JwCrCmrIazLEj8MHvjeDK
Kl4IFUfwfmC20CT2gXbVjEUevOkIWzt9mGhs4Vbl5i+OZfLYd3JCJc+PC7z0ejo1iAPLe1XAupHW
pf8cgA3oAhzl5onrdwn3bzubn2t1E7QvfGVSX1H9sJeCxkCsw7SaqO0b/WCEbY22Wqe90UKmfLBK
WlKSHfuIkNOlkD3zhwgYR11/CWVo6Z2g9hH6AcaEU7HieHgx/zmCbOfzI1f8Zh8CtiviM0AjqU3o
3sdrXrPU8XjuSyF6eX+iSD/XRpbcM9mwG+EntrPZFqZbf01tnusqy9KEGBWm8T8VuIue+oOy1RO6
JCC4plBEgBRP9COk7mZ8+DZzjC4w5UkLYDFvHGp5OojNvYDE3ye1pKJBHJfsC0bVzr7ZpdW9VGTk
gY2uDLZ69JTi5IUoxGsSN3GMVTlVSguvwBqlAdZAHaPK1YUQNxzghOukuqaTu1Pz0Vq0LWiUkwE6
gZ2AzvZgZ0frbjAnrhxDf5dtruf2jvUQnD7az7if7jb76KejXzWm6h4PPG8hkoePn+hCyjW+gaCu
k23lp8J7w4t5gqfumdf0PajyBOyFA00ElenFOwiaT6Vx4thNtneuPpZJ+IICDLxZZ4RNBstZ1NHj
W2uGWPl+saN5rfBxcGzAclnxm6ukm7aZV7ik7DqEiZM0sP24zslyI4Rdz06KMhHb7ncrzxxLZG6Y
53SQK1DrwMBcDb37Nk/B+JPkpgFPz+2QELhJk96RCKHloiraZIKk37DdDJRE8HgDdkyHOIYvddSf
S1/FOic/lmtiS7RbH8/7uREfJ1xadLlD9qf4Zvm86kYpTPZUzSooeQOALYt7l4DfaNM+BKCbkpH+
uVvpYlP67KJ3d+lW+ZyUq4bDieYwbU0yEfduIVypPl36DRAp8l+o0t1WCezGoHpPD7lBjZ+EgyTo
Jt15rw60z3JWqMiRFMwUifhGUVxhfdIrGJJ2QbB2h3M+JtmEYDflkupyAmM3b7IpB2FU89Ilt+15
V5efGhgsvYDzCEb0ivZj2eRhzITTdizkajaZ/bj5t4XFX4cR+btUx3uo3pV1gEjCFqifAojF1tLU
YfN41jRPjwaCcyvEIHuage1Klk5OjS9QdaIa2Zuowx7cEn5SattNK4x2COIJ+wtv9ABUhiQ1WGfQ
+ctfyhZ7xuFe4ww0QTRAI/tkXWImI90dEMjZmHVXcSvStgdG/TlVqkDKTR3kHNBZr5fM3mBiaux3
xZ7ybUvMujvtD8BJ4TUduNER3c6cU1YCawEHuDVayttXbw563pkD+8o+aAcnjUPrJeDseUeS4lND
vM1DQ44jEzTGxC2DZvzyii6ym9AG6y0TpftXgWhR6qa3IWG70VDpVTZmcHfwR4Cz9p3tC/jK8O7K
3r8qh8I2seLVeSzBXhYSPkeGPY9kVuD9RdH5YiNvKsUURQl4WAshiuGG+7ECIMrtjaUhaqOnJ1nQ
I3QvVqkGZjJ4vITwHaKGvClSy6vDBxdT/W01eQNNvf70znmpQq1PRdjDnL0NfpfY9656ZAPNoOKm
IONDq3bqFJYgBLx6b1losTU4VON3djHdbditfFvtLdNIU58W7sZ3cRiLYgC2wjL0EKF8SCVD9CbU
0SpMZYEtRENXtMPfgNi0FeBOQzYEruvJhYjLUSdIxmco1zZUCq2yX+cv5IzMyjqx84bv3G2/E4Ix
DIVWLWvQxawc9MXAirXpeganYFLI01ln7dY+peW/eAaRyGczSiN6CfHYqKwIxEgKdI87XbWLpfYT
GcR6tHy7HYEO5SIoHsocQ+PehytRSg8GQiT2jK4gwvLedFZ7hdZtLKSDVlqImRkgC6jaCrxpEM0t
DJAIUDy4eg0zkY8P/mMhrrzvQBZbw4qHz5FtcvigzyFhc1YzbzqeM4lCNzKIoDlw/GvDLjn1/S6n
Ydf+++sqdZEiYP2RYQ6/ZjL+W2TmNslO+m2TdKwypeGY0kQB12bWfK85iUG3pMSxH/B6Pt50GS8b
6Ip6vJ6R7n1xqs/mfGkSrCMTgYiiSsaF1lLjEIDyQANSsUAMnRJRaUabV3hPq/nxK9HeenpcrLst
/PK6dys+M1mr8mm32f6lekkjX31ZCAdHKYbolShj4h7uwP7X1pFE20a6w5YCqJoXPrzWI7JtBYUm
UQDyFcbYTqvCHtjYmKJ1BqMws9dDVkjhAiKHjhOaZH4m5lsGzTIm4ETMEmfMAUYiATnzNIwfmaFQ
eKn5hohMRNJTTllwd6QJyslJ2cjV/oClXDI+NV9wmW8X7AzHtAAfI2k2We9dC9I4tx2fhQECJ4uP
Hk9TvYPQGjhh36FycnEJbrFORHEEHUfXtmLFIyQsmP6QuHg8I+GJgKRn9gFsQ9VswwspwmxEhoP7
dPKQIxX5A4Hb7bOx1QjC5N3HNCbFxiDwgEqsrJo6kFh2bxE61Prwi8QHpTw0siQMj/A1UGSUbOY7
yuJtyWk3FllGf34S13T7MTI7huYFj5VHFKHhYIkq3DunaUeayecXXW6CoEGpdZnLNFIykEgRFmZA
GSsejxReVlSaWO6zUaJdn4K9CGENEsG7lyOtaSgZsYdmp5H9AR89lk8+3RWqZiVR5i/SLpWaxJLN
C5W2vpaIjTeRHoHpJu5T1AB0qwyJ37ixpo+1ffVUu3KXayf1ioe+qVBHBLe0reStfd/VZhfZD50j
9RR01K3l47tgzq4b2q+Hh9X2Udd/iRbFHvvHG2zW6ZrF29LWPx7TPlTiiwghRtGtUisvnIMfwOy5
zdK6mvNBh/9JUMYBWugcNphQKD27KdlJArTgoK99IHiF6QKqH6F7BDuJyeZ2TTvWoEgabEMqm8QP
XgmRb+plVdgx6AoLWG5OJ8tiynOz6rU1cEU4Rrz6ttx4azswKaYYKtkgttHrrvvt/xqamAXMwO3I
lQexbggiljyYvi2e5AMz7puuBclCgqagvjGJmHqdQNZIQX/krg0HNBX2czQeql6eeQnoQYJo4xkg
aRfkoqaowiTY3Ui86CUUOTE3a3KBqiO2514M8AGPwW1HLxj8iIOOOxlrZdNcLiO9PlW8Sth5Hdx1
KNtUKah/P3fVTXLbJPG103TJyA85CPx0Q67WtQmeSQLyxYFbXNGHTZX3aHDpgWOCw7LOK+0hlwn5
32kRdJNZA4pIKh1UvZwjOuFlTPtSCmLMmjypS1iV1nusK40coSF9xsq8aymJos2Nez3C6Hp3yIEU
39Si3oCBurK86MEgxsu33Yf1G/iTL/K6iCnXYRgKSVRfbTWAGCM8H+VuL44j4kdyuhCwGraC+b+V
Mjb/tZWYEK8NI4cgg7TaLZt7KI4x+mYZnoIJ0V/rGh7GbZinzqRHRcEGepQHXx4WGN0fIQLWVlSa
CQOhCY8JrWMOL5rcu4oL3zVhJ0PfiLFMWyFcpUA7S4Nn6q8G3fpMPcns6mEOFSbqVXtAUhD5Yjjs
iQcxzFNzeDXyPPbj8q69sSvqPgSbRr5ESpbnq/UkSew3A0/HFCNRUzLCNz0gW3HE9BSZ2kp2UV8Q
A8m2zhkxhEYhiiyfu5SCLTr+2HkV9jaQDc/8Iz8Lyu7+H5hC4JONjB1HHW5Rg6tyL+jDFqUHg+fQ
r7lL9sApqKHiSIT4MvbT60jSVcBnEQ9UTt3YP8iWCKA2fAxsPt7PSoSAYLgea9sKgGx6nwNa7Fii
bzxvDtOJsu3T8msoriL18ZHR5LyKTymteporyquSgGScZPkUOZBkF5qwUEhUwvCu8S8OFl3OKt5q
m7XZwha3PuG9z8GNugTOrpv5zbPqkNJ/nj64lJLwUlQNLhTn4evgNRBM5M0++4wv438PkRP33LIC
kxYJC2+4SdGRvB2An5f7Is27HG9hI5oYn3yL2+DnmkvjrbR4J7YOarEt8XPGWcKPNWpbuIXDx1/r
zpwS4EWZYQ1XroLqJD7RlPSoPh6MpKhKgO2hlSzGdHaI/YgASOcOXASpTPpuhvQi2uaplBFPQQ1c
AzR55sCGGepFsPrAtE+QDDIwdt0i0AD/W0SjA4ZpfbirWeV7HXKeq3uxOIVwS0aCRvwb4sYFg4L5
aflIFJgQSDQUntvEGBryOLWAHsj0h8Rtk+6sOvRLtYkIpVwq59aDf8cixDqktFtvk1o5AGPnCvQl
k88rutZmjEDZtczuB+69H0fWDw9CdkW81qTFRIPQCEMCwq2fcyG5FPblEFoqHbJ+mmouT58tZeoj
4lfKTJBLACn9oZrHrOpuULUxTEEca3+1tX/8naZJYaXE9HFYyoFOxKNwK2ItPKGogAqShTXm2DPp
TkF05l4CzH/TtZ6/akWkQgfeyTH4AeS5TEjvOpMN6uG9PKLaalbc18Usxe4K4r4ujbG0dR+naUQA
MW53ZPbSM5qPP2pRLkLVVSIee5Vz1V/QtRNvK0/6S+UbVPrm+kN66HrrOlxM7U5TPK93nIARrC5c
oXldJp9zY/uALClz1zhTRyelVW3Iun1X7pxquVktgdEOqQf9XY7fND6UIXvNJOsi44XXy39cUaJ3
etjXdaErcb7TV3mn3HDBPYVOSEzqeLYSHmMKKqZKVVAtlUQetQZRI7RCH8gnjzQd3YZMoHiyprAv
zjh+7rGvmjK44Bf2x70DkYD5yzwAIxDvHKH47EGOflCo4WMv2BJz1VVg87igcwj8Qui5NvwzU0RK
sdxR1lnuxggAYVzlbuXFKNws6g15CaNxQnXkbft45fEz2Nkbt/FjdN+2JnCsJTg38/Wuw8+gxkPS
eFhvRXP5W0HDgXPR/i8yLZ4NHxjliBfZmT2dCS9LJDo/3k3ym762WoBzUBUWhUz0+Q91N8pddya5
1J60brsXeHwrDr6f6qOEPEYnsh568gaUjU8sCmMA76pbBPmoG6LAJxVc+zeOMXmBxkcCeUiVFudW
N2kzpEIJM6hkHSc1Qd+oasGxKnZRYHSe5ITuJV9EZMPHS+MDzWYKAWN9uSuex9o5RCzYSQbzj9TR
hleaC12KbLw9uQwDmpYObAUbjKc9+vJDh+ru9SFb54s9G4U0r5m5OFP1u9MHIgVjF2OXUP3HPzdW
JUZM1szc74u6/CFuLZb9Qpc9/W4uMClvRnn28g+NIkGR7nv3kTIa1fnfXxK1Sj6lKgFN2xleymWi
58Cj20FaS1Mxb1GFpMDtDczNI8S+kTwws6HcnFsgWdYvF07rOJzz5aQdOn8gdyM51UG+r1tAKLSz
40iOMoUOkZ/W0CGO7/GYXi/UlzR4RTAB41+PL80bhaObR5cEoG8lJaUSoT3KVp28SeeW0+6FVFjX
TTMerEDNl9a+w68GzUEZ9+ubNms+Z5ZBNCwBRck69B9v82qpubpTps85z3wYtfTfk7iKBF54YguY
1SOzuq2mGBOhAJYd47V8VtRq2rl2wv5IExLLk1tleXRFQH8QH7JcZbEVb/QllSvuwGq+c5VhPcM3
1B4EqpxY3FwC+yx+RUWHS4dQt6SY5g3+4jF4x/7a1yJJIYk2Z4ZloIHvyfxcrsruMiayVnyBeocm
IzFUXJbHE7wqFfUEi/09NLtp2iftyIMiIPvpwSIv3W73s6wtiBsdG7G2N9DHueW/2i7waOtIcnKp
yTzqqyLN1u+VPhPzvuYzDT9uX5qX9U74PYWb4m4DCC1bfMXIW4GFX9PnN3pl9LKXKYhMKianSarE
CyeIFkniE2Xy+3mG4Kw2AvZ+9rJcex1LQsP+V6QPgZgn/oYks516F8/2l3v6phITGJdj2yFoJtQv
gt2+k/o/4Y3SOmZYWCKt90kwq6c/5mZ/9orNxak9/CpsLe9Cr2qr1ev+uTwsQ3l/8gywyxFfDCIl
sjYSQ/fF1prc2b949SslktSRy/frL3hJyqaUG3YB0EPR5ayTYjkQ5GcN1BrfIlanISl0An3zHyde
n6C1AnxerlHiqV8IxFbrp5HZxoOy4Vz/vfkAfnBDs8zvS3StDASr4QpShtBZW2eFqCOp82iyQDtQ
xs/dmLrQpdkG9yWxXkez5S2hjYBW65y5OgwHwufeOAQANHIA0Wo5ASzEvRiZD1HEdEUgf9s9paNm
vjxVQZLvDSZTG+qS69au9hkoMvZc+tkN3Cr0QeMa4Atri9I6Zv3sYk8F5MZeXdR/dpD+RJ0Q3lRz
u8b7vV9aGu6NYElb3uLt6F6tOkek56KAf050+tCGdejn1fTF+4TWrCUwf0LZTFjpxG9bxyCElHSE
bqVlndzmb9MfdhV89u6VAVfJdtpV9/BSq7c5neAkgiaxyUG06jDe9cVmFi3axmm2AyasL9Htr9RK
VHcc3uS8KLolpROinb5GBA9aewInvA9qXWfmLE8Qfm5X85hZG7ny4OBKpI7hrW5qNpbVttY4jMkk
J8E1GGkcKiOu3fH/RkHwFFKjYCz5Wb5ItDkCFCHnX1IC5ACDJGplaX3ITLaJeSQiEqS1TpO03Hc2
BmMO5IMTP+ZYVOb3D+Wss01e51C+vSvUlfou18ZrYlAVfhn8bI4YGiLLz4mJLah1o7sORTb/IAeT
xj7DzB8AqLjRGDTwhuO0m48loXY/3pFgpdaKhNd2B1/Hy9VwJjbzS8OqU7yuRC0rPEBru0alreok
Yd7HHvk8bb4PzKh6B+oPQsB4zXFyx0NjgNvQjWuRdj66aWs3S0hQJISoUMA9W/VjBD/SknHOEM9J
+3+4TdmRAe46L6IRmpCzkgn2XJkBzKaz9ia2XlGmVUbwKnm5PE5GYpcqi7sdmETtk/Y5fHRTnZ9Z
SvNg1NzVrAodjlGL0SLAwnU5nqfgz3MAa6oiafSkgmcWn802RjXnDlBLF6e1A4PSsnnWCh+zDtbD
Z2dhs96VHz0HRA2tn3NnBt1ZZVlTlRBNImPhZm+5qrMhPcZXBb9C/1RIRPquAiQagDa9p80gybe3
Uu3PgXtOtBM1ymb6BQmKzu6OsdDr7z4yYElVkDm886bkeu21gc0FfmB/alN1fX/xU/bAprVeXaAS
YfNmaEvaS+AKXXY6PTsuUCktAbzgccc2aEabOvF1oqXPngxUy/+OZtFMVwbT8ODDySk9CGUVHRP0
kNv3lvpUXgKxA+DFzjQb6x7rPXoIU6o/oBM+nqTnbihysMUQ4OIohIAzX1dG5smBez8SIePQiJ6m
YgI5oUskkTV3lBILXx4FqtB593uPar5aSVnImCzgi/3ZGxHd+6Juvl9cwSv3o1J+W/HqTJB5c7IV
L1t/JY5EOXvg4kLQ/jDH2+L7wU0yg9Fdt4LXoPMlEDQQrlzU4Py4nLUbKQhnBLf7uKJAcpQH7peE
jnLhOcYWU8tFKuwXiEJT2c9Jc//MbsutCcnO4Xdygr25RZV3Rr1A66Sv+8twPcDfeL8ADjAWtqK4
dJUOjjNRUypE3BqcxYSH5BePNGiEiQzHLHfnLoFuvI9HvHCcuPJuF2aLipY80fiEdzAHmDelsJn1
BKi2JpUIF1K6kigvSK1qENEtg1xARBV0K5he3D7FRqwMsnlvfSF4Yd2Gc2mpQEqjsyMY1Q+XgzFh
zyheh9g7gCfYnRvc/DCnoc/JwbxRKFLOJvdY5LFw2OW5+xehysMp8eYesuvY8aRCy6W0zasVF4cZ
/jLaipSspnjQDJJbiQghZzDlDHwowIBNhP00b0oa+XH+fOLDhLw8UYbUWenzsOpZoofYd2Gimpn4
Q4GGih3EIFF86TNwIXywGAlWtG0uO96uDq7eF5hHszKVXEjSncj8x98s9ujnWnI9Af5r63vsUKNA
R5KfoxCpxM8gOwFZ8cQVHCJ1P+oFxNbv8r53AwE0OJhJRXxDWI8gpS9afg7leU6eOT3KBFii+aYR
HNQKGiS/LmKbz6+Lsv0x+Fq2Xybbo59QWi5QinHNGQXOxaBxvMu5IFfI++lSzyJ1KhCIPvI53fvJ
GzBYTSt0LGfNEaKIU6NgQGfNBeY3jwgfZHAPk6TFI8TrGwtDrZrSVJZZajpzhag2oTJtKR6/FzDI
nUzxwbEkeWD6/RU7jaBP4rugJzx4b/g3t11OLlT7kQYM7SOgB7ZfEnBQSNfZrf+Sr1N2IpoogPAm
PJ7S95Sz/Ard7i5CHPMEWmcsooBeorkOLTF2InHPbc9/C3KPCsmjji5jT6vZNtURC3i96Q+mKA+R
o5or67jo/YoZ/xeOxhlOtDnCRK9V0HoGuTce7c71x02tH28kxqNqzJ1hR+VD0d8YQpMI+xPL+hQN
8FWR4sYAuNphdm9R0d1YemGhIonO8HqxZJ+bwkMt2kfR3urSNGAWw87ZpnjeN/+fREx6smEBJGsn
asijMeL+9k9iFaMmYZYcUIUI3SJf6ZzkPfuNJ8fRgGNzXzYjjks8Ynj7KnWhlJHf/ZIhdAYd/qal
S4UL6kkCqo+YrZHMu+frw/xZHuAEMawZLQtNwoJyCBz3z9N8PyGpglixfZ4tr2AM1QdsgLSdexxl
PDhpyQER4uUWRY0ugpl2GoxYGNSNbFZIJi3SOiBvXfF4Fv6YBgy3r7D7/W5W2KAL1kd5vH7/YkCb
0wZruOp+2BtygFvV/BTbzUDSpfg6/DsjfC3eIqLLxsBnsp5GISa2Sj/yev6a6RQDLKQkA8L4deV0
s4YW461Y1dmQ9y/lFk3Tgtal0+YWT40HrVQDAU7xvWTVcva/14oWWSCCyjiLvStv6CtjAkGzfgSW
O/691beIn/ZekBbOuJw0JgNCs5RdGcVJJo7hk+fl21cwgdiGztNgFXVZWjqZUp/dZrmLp8KGU+xg
0fR/Effv4cPLYcd+rABQtc8ENJDHfV7fgPMfDBe/iKFm4SraphJOn14MoJWo6euOsJelXRlGpWZh
nnnzrVtpBywKeedKL5Mo0Or5bp6Dcp1USnuLka3nCtekfz268GgUM1ej2NFtRCSSIuyl4zmvgryH
WX2cwyJa8V9xzMa3h78hBszC5+6D3MRzZBwqF8NIyEMeqHHgeLf/L0Do1mqtsroyJlzxHfLM14OB
6rLngAY3lZVEb3StxpedPuTDVxS2WLaHIFPX3tfiOKQsePvqaZaVtTHovZxVYZ8fmJklXRb0vHo1
H4kMt/KmkqGxkn61RD6MMSIWa4oIyzFjeNfv7SlUrLvqAOd68hQF9IHkP0ZRiJObW6VaW0wo/i7n
nUc7LhCa9xqsZ6wR7wtXpnMUTC7bf05ImSyb69WJwCT1/knu+Nhg/EInBIeefJNAu5l3URc3NGDB
SvzpCivr5Zlvv2nylqPbaOt9GHuv+aA6ZB+KVwUgm9fVNxRwOzo5KIHwfzDAXxlrpeXrEaMFKYW2
ugqYqTutneZF9fuCDjLU9ehdX5Sn0FzrqVHuNjYfiErBbIyl+p6oRn9zgOhMDFFKPhjTo7O2TL83
p6vAYfQpi/2ZUNUE8BAERwO/dUMJb7br4w8XroO+pOhh2QPG3DUYuPctfytU0Xv6cKWtdvUd5umD
k1roz2IIv3OIQZnxkrR84UaoBG0Na5+WiyNjm4mCnIumOwcqibuq1wdLmlnV4VbjVpOHuje/YGdZ
sBSkekZ45T31cc3S2IV7M0qjm5FvnanK0yz9AOYB6JdXDlxQLmVNVx4rHFebSdLf3aTGbPkMRcTm
ctlMuZdaT3iKzxWGc8GpNUbHJbLBNFqJ8+wunyXdjhLnctzTUbbSZnEQGrbSX0LrPRnz6K1b/VlR
z5epM0Htz+ecnZHD6tOKw8OF2VnRbXhqkvwTufQSlbaDlMC5SLaQ4BSxqa2hy9Nvn9vIHyHAq5lK
FrOGMfWlw8an4NiNPAyV8HW+u3IwijnEzS6EtekGwJqp1B2JRVDBAbRwT3fbrgyTKTEycHz/OB3y
NfplvKIS/Aj2ERDvRrBsJNhEzOMCg/ldzAHewuJYU/XHrQhfpxeBgR0yAM5B+NMwt6vOkXptU+km
G00VsSg9mlpfnAZ5W3TwHFFerD3QLS4Xumbh7kyWKEvrzdd2yepBaFWxTJ0urhZa+ynrIVEOFxT2
497h4qf1oFIyKD7Zbyn7SKhIWfAjraPB9AOhLHyr2Jdt9Zx+iT/r8YvYVM+nEdxMVk4t6axgKKio
AeViqjFNAoiGH23OjdoiAv+XjkJwTvdeuBOK3EddchgSVhdxjDA8sqP80c1Ee8m7/VZJd4WqeH46
9etirsBywdHPrzo9M9ZyLKm9O6lDRgwq9+CmzFiiwP1HYkQoEnn46zJdGrlwh3lQqZZkB2mwHuxp
3jg4XhoOBKWoiDAl4jgGCxPUJujzGrUypa5J1cY4zGA/naptZjLp+f07vNU2qQip42jr2l62P3wL
AffJ4RQqsBbTyg7XmxAUC4nty76XdDAwgq1chQAomKdD/tEB7zVsNCdkofRLeCG5vmJte0gE9EM4
kq1ESD284RJJhpuQvRPwMeWwM2m+QTP7mpq7/JSBKIrQzO2/9ROfmwOtkNWYvrgsUYYvdLmwRlHd
GEFlDUoGOGd02OFjW1XlTSQMxpw/pL91NSe7jTk4ttMT9gsgIbISOUPjnSs98VjQqrx0ET06G9Za
sPtixJcODEDdY719d0oxxOgplF1NMsuiz9hO2onPoAMMKrU9Sg+PdOd9kL7QVvPZ3JR3BdXIHUMm
Z1Jf0nwqVcRZkiom/oXMOXubHirsVvMbav3RsExs4AqhpCqa9l3fMw6hBLq6J2j/Mw0QVNCOGaDq
5LLS9DSPMh95E0WlTQfYspNIYcg1j83YrrVLFEr3gty3+aLR9kIKk3ymWXFIOJabeyP098IuEnEA
XnW5XVSdcw/cF2/bjDzcrI2a6jnGOMiOsuGvNVY+M+q3k2x6hB29VL9VmSpJvHdUdxgnpPuagwZI
T/6fXV8f42L7roPK0GWcUF7aN47g+M9VVlf7lrDn1FYMLWsvI6DmF218CULtBiFOhl3OJ5gcRYCU
HuZUV6ELfzsVwZf6uBsTYaBXEHjErMbI9AGOZbWed1sFdbtUhhykbC+cdbqrJVgaFeFHOks2gaEd
xEivkuc0mtVXmRg0BZJG5xKQZvrT5bkss6/GQpHvPwcmOanFPHyoDH9sPgHUrclPC+kmVMb2MwIz
9dFM83dw6CBP2h3t3YSUXVdAv+vMkmFxkDXfClSG52W04P74no/FDCVEebfMJ3raOdlDlIHAs41q
0X+9QjVdMjlPs+Zu81QQ5q24w1Pg9sN2GGxEFt0ioQNeRv3BNAUDOM9nO04epQEAO3wj7zg1XtdF
6g9cOafBP4HXuUuM94h3A7+9LWUae1Q1pl1oH+pEaTnzYCGHTaz2ae7f/QeTE+GUjQsUxKDrMRos
yVzElUv13CL6n2PvaD7t+q7kdlHcjh995Z1InR+iiZ0pgwDZQMeUUUF7RE836dSvcHWo/TKNE46+
/1lenBoao2kXEpyYDN9Qv0471qxsNidwCr8Inda9GcEX9gJRrHlWwnPrB/uXLdSufy8ulX63CMFs
S31VI+aloeo17re42qbKev21kB+UPOlRJuc3OCD1WU8mgxuDtQQjYw2lfR59S7SjMgLRhouvDLaX
PoXcB+xwew2FigAUVNyZeTINWfj9iupZ5bUfPkhxXBK4bG2JH/mH8cmBmAbabneQ0JY6lG9+4OjU
DbDXX94cms2Qlm2IHbHNWOROIvCndiIZpTI6Hpnfa/CO4gj9nLemEAeaRmMqLIgNcKpfH8RBLDC8
1PFaKf6yEwbjqMuBhfw7btL6cHnaQP5CuPaXWOxHokK3Y6Lt66LZRFxtArselBQaS8Qey+9QfHr3
Ps37tNxxS862w+04fB/2KO8m8JStWcojULYKR2sFAJkidYEGh5HtdS+h9a26oqEQMvjhSQ0j5tf/
/5v3LrkmGoXuEW7QGpGFv+MUzaPKi086LVDMQUpDBc8qdktNwkOId+zG2fvBrEKaRsAVK+x07Z7X
FzUPrJemgrNhV0CiDCKGWxG/txN07CM+ReqEEpdgxbEPzbrZjPRRTHA75169YQAsm41ojOX38s14
29GmbNG79kLl6IOZ47xsv8Irb/cqsiXgqGtLNEkGZeM3T9+eZ5GvTm/Tu7eK1F5WCSQFXR065R3c
+LJVJdEslnfI5GEjZtgt0xzS+bRyMgZlFXI2EkbUrH3jZ5KzTSovJiKp7/dhSmd36mv4pPtEHUWJ
ylGxTohqcORRGQS1s7ytt5NDq5TyY7qeXC07WheoIPS9EHnWiRnBQGuJmX3eOk+QV8u2bc7KwtTs
g33wq1Kvqh4N+0VmCt+JuT1di0LCt/HPlVi0pyuV/f6Zbmvu+UPbanO/lhGI8UMgGEoOOvrbNDoK
2/F8caDjbwhZD9riQxtgbOHAKsNTwoiG/zRSUW5VMfuWf5S21HNlNkI7IDPB5OCnQCKJtfANoZUe
rwyC1n9g7m8oqDYvnt9V80rLEaJfYLSlwTIhjUPxeZhvfML6qW8o91peDK4CKDfFVOg+1c/oUWlF
aM4bZptok4rnYz3lB0J4tFT3LL1T8yUt9cmH6Dq8kgFvsO4+2nRLCam4MxiRc9SGSoUhqgUD13iW
l4bstDLuAFpVX/guo+wyeCAqcO62cUqQmlgeNyr5JNQOlSrvh3eQRqEpXi2eaPUkdtooyAkYpU/9
RQ22PrVTakHddU2s6IIzzQl85774RLgO3XwvEGYuF71YHyPjIttOZfd3iWsx+xNlfl3ikuCO6NcF
aV/UwB8o+UIyUEyBXwe4QUObESQRudhssgoD1MXvveGYQk8YAHPbd1ynEOessXRy+LXrg7MfO+Dc
TRmk696p/JYPF6Zmv1gYXc4RG9HmCRmdPmvcUinDL5s6bQmfGS5y4wnap32uOF1a5qcRSb5fQhS5
yIwXG/tIOk/lAqAoxywSxFZIPY1gDp/w3z77r/hAp1nV8SY7pWNoQfvljpwv4iN2jDQDvAeiBiMU
LBvfRvHFZQf0+aOn2yGxpkCs08WpwmAiysd5LQXmWTB9ILua8CAbeilbSZwpxrdWVFWZtHJxeYHa
/B8OiaVNM/BsDOvGsmtwO6FL8rJM3IvBJpI8tSToh9dWfwJ0/ucL9brGn8A/W21JMrJ7oHCh3tZs
vbumOwxIveNmgJ5956IzfocdKDDWuYHvn1SBtrhabQENrkQrKbsyChDj5LewbKQGOMyWEK+b8x3+
7fJUqjt5awjI86gAkmXgsFUROVowf55jLhuur77OaTec5Cs8pq0gjwQHlZnmlC+ESqdFeX16zAtO
p6DgaevDJJpFyyd59o+GXF6mpp8a5JWqdDOFcdG57j9ph2Wjp5uBg0FCuWZZpVCc83lTKHvZQj/6
+5ju+Y982+4P9bWKSROiujCFP3J2J2uuU1LDlSZdcZSNOzeLqW0rfP3t3H5qqY11f2GxurdS9dFd
W2xTesSs7ECh+m41nd8SDjf9FZDWzEy135+FiEIvhFzwQbHSTWsXtnQl6T2mf6TJvUiyc0f3kDuH
j4I+ttcVxcOvWFB3MDM8K52yQJBzDpVcUpDCOS4dibBS4uEU7yEguNXGV836gLPBwcOZAhGVa8AX
OmwJ6j9fdbynLaBW/UDaZopwCMV1+/CwnoohJedzS/6291u68JCEF9B6CB05NjQwb8y6bPLvtjxx
vfiUHOnfhtPsVPOW5nC3VyA95Uxu2P8kD3Hhq1dxB3rH6P3wYwA5gHXvEcFqQkgVMNF0qV7iApbc
0rxjeDZEOSKaQLnxJluhEDXRuleyLE/KtPADh04AxzEZwH4fugr6ErdLshPPTHhOVR4fg1wOGy2/
WeBtAKz+YHMj6Q2/UO0MLY/0nw6IH/xpojClm9xNdlshJ6QWivBs0lzmonvkPmve5a0vJDRJ/+Ek
QPA0CSHa6CovaYwpg8Mqo2RB7Hq3Rik573484JO2oya5a/mNhaH4VoMOseKXbHJIVcrwNaQhDBgC
0/9/zlSlfPBvceoLU6BVFe4pmZTDLDexZc0QZLyquex5NCDFbVi7SPf9GcXc70Go/pctRZ5YBAqs
KQSuN5nXTXeggjtE+FxFCBuNf18LhFeKzRgs8VPKMSgGffqzXzAB0DepdWLjDL/ob2sfjJ14Vs6i
JwzexkMF9xcOfhfVy0H5pMkOK5s+23JGsFI0badiQJ/9ldy2rEIEJi3h9Jn/+ORs5Fdf5TcUUyyF
D/M9eq0WDcwBAMsPW7Q/PV0GE/8Ig/pyF3VFsY4EP0VCj/XJiJXhDAmOzUYr/H6YhAbk5VPs3F3q
waLlHpTb6f4M41UxiZ4D8kAeW+ZMzAWNYNFg5YWRMxGZ5KhnlqxKpbg0I4Ec0YqRJyKf81+9ExgI
CqZDIKwv/YBwPA8/oEzrekO4421DHZEhxxi476+x/LnPNR2xG22ufEhz8EzyrxY96gBmtCUF5gGT
hgm2evg8NxGgDUKkPXGoB2zOrGffJTptUeOWeQwHz4MQlraS/8S8FcDFOhIvvCsd6Zn8B5vx/VLW
oQ94MsldyCOmGvAJ0+hIxc1w+DBiYsRrw/Aij+LHVNPV60jbaghqUPD4HfXnMhvP/66tZhymaBUj
K0daqhJR7jA3RVcuSw/9EjldWqI/jNwQsKfHvoN9ww++cpSOj0XLYY1GtldP3n6LnKcAR/V/P34Q
4EWKwPAqKpOhVHX5vgEofScpgAkBkBGhkcg8H/9fzuEXee1jS4Drui4CjwcQrVBAcHbhdjjawqOZ
vgsL2YWde5DbZFs8JvEhojXJJZFUDhUSmQ/ykw5c22jSB8DmNGSKb5LuZh8Yq6VSHo3BC5kk29I9
MZzHfdoPS9TBhzcF9zu626C1Hz+GrYfgj2JK8QuYLq58iwuM08cIvg417+nLbRHb21mbsC685B5m
8z+2/T6eGMZKqKUo9uzv2uLRu35wWmILq46ixLcLXkQzSAvKwPwBbYxWhCBtzBntueMbTSU0OVDI
sQZZ9U03tGFcviD/NhduBUbWTXfjlAS2nEczSZfnay4fCJlP64Sg1o+D/CBiagy31qukAJPmdgSP
srcuzw8gbulct83KN/2Fe5EXXgkkrv+H68Hm+/19B1GqvQu8PLcVvL4nz+kUT0K7Ai0pEpLZE+3o
k+m+vR8qzMfQBxa0vs1bWv1RS/Z9xjeLVsaXIY5GNmNmG/b0LGunViW5q3me6n9lpTHiaSf2EWJg
IbUfdplcVfmCBWm1/LbkpokM5GIDIB5LykKZuoHSo9njhpUQw+ukR5Y/FLoqxkPbNSGsEnltXQhF
kS0xu0wP14b2X7VdjWqTtgE2NWkaMUV9MKdOy44zD0/LJP5VSlkEPrWRqP0ajEFlfOd/In7MQ5oI
7y387Gw2qmxLRKa5zLTqQAXjEcqnOv/TF5lDCAOLI3QfXiQcZJ/drjwfNDnzBkyvLBiQdD6qlmBD
PEsH1+8J3g0A0kXam7u3hLrr9ktWZ7iBASeDpM2AOGJ+845zsT0VabjtHxeCyNWAhxkJwsKy5Ysz
EhTJVKsBpvcmc9BFUYXCu9X9BZ+fn0Z4kiamBUDR/+BRE9JG8TVEA1hEbBOzaaS3dekdQ5y4//iO
mdbvwyNMnLoRnzizt6kh8FNFUSvBpYBiaQooKFfm00y95h9zkgBzF+CBNj4RaXx1QsfniwDcWHqu
XvwsGILNF6QbJCYGu+mKiT8SWgg9wNCvzbTmcQv4pi1RbGrDQM/b1cE8wntk43aUxX2VSFxcrEpQ
yRS/lCN08LOXLI1jDxwpW0afTupojXBjYQwfgJcxNM9LX86qrW/Krzs4TSuWUz3D93IMgk80DjjP
TrmUJ7rUrdfrmaFARIcr1XFjsVfXGE1i5atzWSAIa4zG685ZLMsAmueH9XY8oG6MR0Q97OVWpbmf
ZGRKGKfthCnyOBuG72/v3dDF1Cgf0zb61uQKznkasCJWV26jWqH+bIkQNNOhbY3HI90uqAnieOwv
2ialTcD5s/ObDGGIXP1+boWy/DUV8zaJdMLEtzfqitSLggXBVPUSy1okPD7LAX4eRB31alnQdjvK
daVIDtk2uoZIhh0lgrmIqjFKYkvus4mrUO1w5zLvCXEujsh64nby3EmcwAm2KCPzixgLeVZm+xBM
HRdGaICeh5t+AxnCr04rU+NAI75O0MNdpxKmfzloiLk33c3kRDeVRWNAnd7WCslmrJwzV6iHmNrE
x+AevQ1YZJ8JggNTliOvQMfMjUOCZu3UX1XvFgZPC9lIBJD/U082YozKof+wOuKtUmmrqvHJkO2t
/rbYOLYRhsTmEd7Jhx7O33VhmnEV2VgEzDMk/ff33IFPj4oQMt/8Cv2sKRBJF/IXj/eVfvo5tKDo
308CYZBukxWJW4tjfSBz2KGCtr9Nvgwc61i91EfZRY/b2iIlD8w1q3NhYv1n2vVdq9yOARsZaThB
cJfrKV14v+6hrjumKNB2lEra/WT4q93WBUNReWylZJ88SKXOqls9DIWEhilFzlffeGXJHuIJg5rq
ENvCS+kmSVrA+oSXIl9CyQMGd6cNvHEGz+tJR05x81Yz5Rq+9yJJguUMUoJyhUOztK/Ky+XjZTyQ
fi8zeVsBkhjctX4/G2spsdvUblmM+B5D9xqBa+XiHo/h5UApWs6ZcyOG0/8+DTWGGTx8m6xpXhHQ
cztmkdHMHEDgYsfj/DMY+RaJWWWwQ/kltpRIA8YSinKVh2ZKx6rPwGRUIcaDIfAYdcj3umQW2rik
2gC/gRvToQbZcYHJ81ygfpf/ZcxvxfaNxw8JrcG6v598xpuANHgFJMDdDZm+wEgHci9Y8mWjjo12
9gc1DkJZjc8tKkWRsWbCVLbZlkdA9Qu8IN50JspsJKMhbvAy7TwhRY4GqfY1yX7vQAtfLzqdqgoi
JGccKMpNjPHJKyzWXQWqALYzdOe+NkwQKDrytqM9mZmD3cNoYxwv/1RJ/E5IGessJqwEdILpD2vX
03fXmfU/PAoM8tY43HGVY9KM8kxxx1Hj5z1LB4tROdqDurIMJznsg/s6yRSHHP/TsEIr/W3IEBSj
o5QR6G8c6rYIyn0vJwzhX1S/pzykzTv/HJNKimo13C0LPl/fc2njR8edBvsKic1cNAmgKrZJM4Iq
7XkEjFBetyeVTTdyJ7EUPSkD3GXqh11Dnwnj5lhlu4+VJT9E4wlFEOlYniQbRwhz/8LSKJhhdRRh
x2KWIWMH9E20lSa5Yjm4mh3HLvazLQQfVANKCazZS6hgvF51upwIHDD3QFtYuIV6QDkz5ohJsE9A
6PttdcFEWAais+iuT4WsAo80jSg/9htY6kMwrtp2xjADXIdW+oqSpRDpBp7D8zbqHCuV+HH+1Zrc
Xoe4vFJpzAVzHSja2NDoZhEZ5tZnmoi4lZ/2I9qDTlHPAApgJz/l4sF9pt5941Cm+w2pRpzeNIjX
hstC47dzEAe0yzo9Lh9QR8olTllDz6GgADcaTFySCVb+bNrMZafGsRRy/e42coxuvkTrWb3g5oU8
+wDPZ9QdyUQcFvuDWrZrA8sUW9gV/iDVnU45OHExPtCeda4jAqi6EUfgz9HIykvAFSqeauQfSZlx
4CgPD8aUEPu3KS3LOFfgPmee9wF9nXNy+TSU9kC/qp5Wm5zQSZOxeA4FlVBNFWlhiNxmfyLRLnE7
56R04cob6bvvH1OsezdFHnHQSaTSq/RncAdWDMPqtieNjd8TQOQTK2F500FzKjvQpVrFrtGt4zdU
NtEJIlW98BztLzE/r+XlBJTaMWU+Nmdwd7eQEzsecCkf95zeRuDcNP26EUyrhwM3Fz9Iv9Jg9y8S
+C+2nRShlJDvwcqCCPeTEJIdg8a4UZnsE5KpQ/GronqjH4wmO6xFIJfSW/yLK+wCvbrv7a2QrW2e
1RwgVZrIlVCOK9OPl22moKuFAtTXuzFLuBeis4BFhKrRqE9eVKE6MbDq53dsVz+AipLWatsipSVo
Q/rl/B0/R0igoC3lVYJ5mucsW6of1p+fJc3YC+tS1KeqBSxSVF5huRmCvi8kZoYbeL5zWivu4gxD
Ia0XDW4V7kA9eZVZvbuJznMP8UwxKiULt8aEoXxrL3++Gqi3tM1N1aYYNjtTn3eojnp+0I3GCrJG
6SW6w/oOh/uVUjp4lOIxyAZixp/8VF8pGIfBNa/WBwJ/2Lu0uuiLD05No8sNBkPwtG7w3PnXGR1H
VYIeymY6u6g5rAzpDpejPQd5QWry/CpBOr/Ev6rfSqc9uwgXfmoWBHcWxKAa3uAQyzO5jAPlVG4A
j1l830jFY7BHTreYJ1yJGFGHI0NUC/k/8hciln0BrW6xq9XNzj3bgTUGUrmL2T4W7X45QgD+A0Zr
CKz2/2wq/Fq0tB/L0dFiU5r0HecNG/Qt5rxuxC4YXMacoP9S7kY/ke9GsELEjlkINZIQs0dlZl8E
WDezKTueHH5KsIwXDEh1YcPh8n5mWXbK3Ka7Qvs5AKglapy+AzDVg9V/4nXGeNZNN9UwYJiRV8cO
+yXNZqEQ1XbL3fkkXLAzbzp7f0KmPL/DJvNCd8Wu8ht/b1sldbBK+KAsaRzYJcO5085kquaPQeO4
A5xTaHpjwNTgDPRz+G3tzdHurwN56X5rBguOMvVmZeFB0QAswB2Gf/ZpBDkFF244Od4OMYv8abUQ
uUaZuJ4KePn7L4bSGb8mdwYx6RHnPe7PnHynG0aQ5TZqFwu8Enls4KRmbyUDqZJh815Z+fb6whvc
Snf5vGkKbjmRCNDOfZ8t68n/NnfY0iZ+MWabuxHaWoxI2j0Ae1C3lAkjlPNSgyWPczlzGdGYxMHD
FrEVI3nBUbBndv+OdAL9IEJVrXyB9IGeXoK7/+057NH9dB3cEimGNxfMHsa/4yPdXpAGvOKj3AEd
v2aYTHYz1a5vpYTdAiV41AIa/JLfTBZd3NrA4iyt0ZvzzlylO/4pdvhgS1zFmaag2Wg4vL33Co39
xkkto7FcaBXbquTrR+jJkCn2QTL6hvzfdBrrkl2GOUvexX/mlPLu5T1xj6lUePn10apNHcjWhK+B
DyjvtuwJhN+MgaJkkWRedzFRRj+eI0qmKEMDnQb3I/UtNCo1FwfQmTMC3xkFYkZGcR5FletoG1uR
z2SxNh9B+OJiidaBtxMvp52lnwbmdspZRbwboxHUcsEKds9L9ntb7YlEBHzBexNULjLbUtC+NC54
gW6PqXtv8XPClLr+7Jm+xyA9zcV7qt3Lme0+sR+TlV7GxTenLg3BCJpwXR20uJJtK0Zpgkti2SzC
UBZVAbmZkdbmWy3H/sU4Fg2UopZw+WzHIk+SOUwP9ywQF0+3AIm/Qt3ba/ebC2lfPqmZr6dTYUZ0
lAi/IJHYwzejWmOKf9cw4wYWKF22ZdIJcB1OTuQabl18Rv50foPK8AyKA1Sj0S2HJmGnW5Ibz9M+
+ybvgnAMdJ62wfkrEdSGMgzXfPuzlIBzuIWzArcrr5QrJe+tuzjschArZEYS6gHI16BO53idVssv
+YtfkjLbK4T7xWrK/Z7Oq6EijJ36X4fFra6xNrpPSA/ddNrl8Tw1lHAuGBlY80dMikf4QHzGTK10
NjgVnOnzEWZGmSAVrRswMXwmwNTGwqKPgNZ15gRDPEG1ztDPXcAl3yblkS1lywMKxlv5JNrzhfZ2
gD1976QEqcov4OH6ec4D1JrsvVZZsif7YqIZbL/l9eznzn4qfT9pu41QqVN/WY8SPxD0XbnmpsS0
ObqoRjNGz0I7GlwH/oXmTKNXI9gHsbmIIRWYRGYKt/nL4SL9QQocRXTLc+gmq8F51Uib7km/nmxx
kCDde71eIHqfPNd5w9XKy5eWPp279D6j767L33VqqtXeQACIb9/BVZIz25iENmYjrR/fFPm8q8wt
FpxdkP4IZjukYqd6kf3EpXOGuHwOzfa+lHad1yWsR40aqsJ1XJcEo8G5M/+FCw6ZkEAkym+Q7K6Z
PuJCoe5KCuoo4DVBJti0D2/4KktxD5Mdz1K+EyKSjLpjQiG2AE/WKTj+Z8J7CYpx0oYsNKuMK/NP
jwDy5DpS5CJ4Bt4W+mSo6gZQTRq62woZS5HkFCcGjAw0e0eFjKlCHW6NEAAMbL9IwrFRYZCxKqsw
Vlb4zf2sp9BE+nlRujsYx73QBda96uOvGOSblEzm6ReE30yy3gA0u0q1bEoujUZ50woiPdP2Ai7h
MjFEj/sKgcZXQW0PRIK3GMgbm2t9Cq08g7VWDbmAxU8hw/wA5kI0yWeq6JhL1fD6TDdVcOJZEeXU
DBxoEENuuMdjYcJ2bg438X6qlf2wQ7Kfr368IiuN1vQ+taWPk7MU3aVr3ElZpmRjYedRLiM7gQ/c
UNs7S40zGsWUz6qat/GRJHSZnvKxrMhL4+F+2Ex6cVAn+6XRdThGF4agYXgIFT4Q1u8vicu16T3H
CAIjdA0vNvbdKvDs9RPmQPKubgB5lfobW5xzILmpyy6tyXosaL64Z1213/fYCSa/BZ+Hm4Ph3g87
bVWdhXBiGykSJ/FIbU8AfwdtqToV8khs62kyvVxAQLk1F0i17jup0DZtTCCofKRdA39mwIwPJFhL
fMzP7uUYWfE9+VrCdAyhq1Ogllwl9gnk8gvURVVj2DIFYMc83HyHbG6ncT8MKMzyF/y98Bvi1PiL
WcYirX4AS3boxUwnkK8VoC3ik/Ns7GNiiDhQx+nb/T8R+9wa+ia24dg7nuy8JyshhmyLmc0H1J6d
TZBxpEKRtkvermS9qIo1ex0zVfYPad/iwzLahcwNyRh7fOkB7w6g8HapjwfNSbkxhjQO3NDTMFxW
b7uuC3Nzq9jriaRFPniDvLqYQhgsAST6jB1maMVZQbEai/ORV7AWESGyc5/czrlz+0fxvrUBydxK
hoMkHMwJ9gkEoBkQrPty0ahsKiAQFOoCiNvFN65u6HnNeL+SgCUqYzENWq6ZYg1Z1+o/msQtumct
9eoLPbk1/vgC4OXkTVua8zR7SO+cZQL575DW9Yqm7rhE18Ct8zA2AkdwMQtAxmUkyK0XCK2Gz+1n
vM6KFS60ryVZuQGqk5kSg2JNv+//8uH4CWRQvT3sHYxzQ9kR67nWn00pl/T1FGV8/7OCIkWEKiG+
audEPjvWjiIy0D5Pr6QNUyGPPRDaLg/wp/eli8ceiHZOX0SLIGKqw4DbukIcny/Sj3oXIyRFjfYV
kbd6ee6oPR9yIAZYgC/mQ1RixB+xehos2CL4iM4Nos28OcKJTePrZMiNlMKfPysoW+3pSPLs82GO
sLTyHUIfCZkJQuZwOlK/cfWou3/DGWCkv5bcF96F+ZuBp77SgO3lreUyErew7UGj3AUuKm9G1uGk
j782OsxLyZCCURAXgaRaoZdQo9mIjILn/Oe2+nRZUXSuT+8ojlFM8kb0jnozFZeOdk5jKkzpa6Sd
QG0Xf3m1W3Is1eQbxNpHWQ89FuL0TFHTM0WiDgzguhYGChHf2KLEuBTCul3atKhraccCy1g3/1aF
QZRIU9z0inuFvuCvpb+jwEuQQtGrk8MK+TS+cQ8ob16dJBivYPni7dLNzez1REOn8V3Ya5Itlxoz
xm/1PY/0vlqDceyWkhiQK24n1qCUDISlhkh4w9LJ4RIoCt4VrFOOJ+Brh+q+d3lKRtWD75o+24k8
iYPKhbSv8WuVO6IDxiQA6uI24X1xvqsgm7o1QiZdndX/FzeD8D/HvWO1uvhC7va+UHEhiQ+gKLoc
5lbqL8xZO6T2j+lnadmzZ1yjL0uU7+4/LgE3Le/LnI5PXxiQdKahvbIORLcsjD4Rf8iRyBVLIlLn
+rzHo6ciTH8BY2ptlCuWXsn+wgio1bvaJkaLRba7z86fE1b8QEQfcgcIE0NPwCyf5J2lVRbWolwK
cnp7PBBbmC9Mp5DjqknlfMXDi4A24+saPM/C+Qq8Ob2OeV99ieqx/XP5MV/S0vMpBPpVnRK6DS+c
r80+KWgqbQUERE5hVluZ/TGJhsKDoPxuGn0/46SxjCQRVg5GJzJWO7CHhW70N0u8OxKstRprdA7I
sYymbWbHMAfA2lB8DugfvbU5O014SuObmL1LrWLR+18CHlh5aLV10lUjgmBFUGYRilhUKQD88fJf
INNrwqaKU+fWfVhV1mrNyN3CfEgPrkN3Zu2SpUqKeSjMt6s1Kt8Qyc1UXUclvAPGpYVTok3W/lwv
/+0s9Mhu9f+3+o9BSCRRWVhTO3ykMk0CQQQ6iiJqPmbJtW4IZAwkf0Y1QanB0Q2jlp4yAcw+3ab0
+R4ApwEc9Ih1FH78ZdrSPVXIAx6iSMLb17NUsKGWBvDcSJIeQto55raULvtaIc8SwiqNfmq0gD37
L6Y4jmKbPDpCfIZzPbjLHkUl2Ulk85m8r+aNcdlRC4XizPmWhG3z5FNxSwGZC8SbWGuFuaAvro6X
Payev+U5+MairWjPIfKmUD/WKFjkZp/3/p558uPsTelBJml54pmPf8P6NazSX6RTqmjHDeDar1Zp
bkpRFCuRR73/oJUu8rUqNtjMndVoiCdvqydJh4lihCxSzd39nmgVyL4hTb1sKxFAfTAN7vB/DOfg
6yRVI254ZxM1dQbYZyViAz2eJHg+55ier1hOpWapz03vZ7OTz+lH+GsBB7sOr41azx28GpLPg43q
nJ6+zb2gJtMVrbCsC2RcCRnbn24JqIOTYagXx0AVqY8y1sl5F8smiu9Sk4Q0V3/DCy4cdVgFEsZk
otUmfLIWqB49pYRZszdLWKDdvDH21CKnUkd7LpWynDLaYY9CvIxkkE97KPeC1pJdWOKy7+g+l3m1
TedeGQKpr/soCshkQ4oN0K8Drj3ft0jJLebDlwtThIsWGbD6pR1vq9oRnphDcoJo/CRuLrwvqxaT
cRYPvEcV8nYkunbewHon00gVR9cLUe5w45O00tGcYR6/O8vqhe4CLvCQt2TBrQxPuzKXZOQ14G0H
1ePCpKUt//2iJmWZVVscojr/P9R6oXrYaLII/2rFTcZ3MjEuYQShu1/Xy7tyQuZEC23AaKTCQYlK
7J2QsrXLHYjrzC5mDSzRTB7CaU/lnzEyOHpKqEfGPrahbdDBZlXGAdUqHYXHjD8xZALKYNfXHv0s
z8osMU0G+uZqN36CEJ2RPhgoKHVbE5x6E6jMvHzWX7o3u+j09fmobG7ObFFIBQjngvyqjZeuoSVP
ga5J5XUtGyolLnRax7zFBfOE9cdg9QSGQNIboCxbNkX5gVMEi14IZPuEC0dM5sSuoNcQPJHkoQCj
zxnLMV0XBBIDJkZ9PUAFyYWq0fGwTHDrpn2XefpF4ZYLoRYhhh5F2HSXdB6ibjUFA8Fv4n2gUK+e
45YqHGlq1HtTBIfieibkEi4npzJgvz28a+sPgcFxSv+QP7FXTV8EDlBt0H0UgodBCJhG592pbXfy
UfJgpp20hageeZScjBRChYGTuDBdVob+qRtVip2YMhMFo3/SKP7lw1PO4Lm636FJ/f0FhZhL58hl
Miwp8iH2WXppIitIsOQVw9Bs7LxeINbLMWuwjdezhFgvlnTiJ0+CE1WISjSjJmu2Z0zyF6XIcI+E
Aq5g0DYeAXz74VNufwGo/I9UzPqf9CKMQODAbslCYo/8zgo3pGC8EM4LO5iOy3ZytYK0XFdEutLp
DWlBExtf8+NV/WrfZcBbpbANMXU7TKPPGyBYSMyvmX+U0mGusra5Tm4eKge+jrMBqLioqExBSs4J
Yv+RjwO8w2iuuvrC5daIt2G6+YQl/6PBYcuBcN8L5k8X6tZnWUuY+K1DMFsB1RomHYnR6mzvl7tT
Uesj5wt91Fuweu8G/ALWOaJTyjcOV06hRaj4meQAM+1aw3UTcLO0Rl018IoWId1BHznTjUDylX8a
xG3ki1C9vg0+yLU/Zi2+0HgXvCzosK4C1FnNT4gUWxWIJ/1ivoej12SK/AgATiXtZCM24jnp09TN
cxheD6ckturnn+Tqftvq6ae9SITcBv+r6wCouCjbVYnRS/Qejt1Ld8dHYpgA+ksa3Ho8wBeA/h25
hWhjMxE69bsXhp3GGp/fIWImkE3xMaX3J131rIP3985+vhcXEHEAxHS7efzT9Zt8r+JcP4tFDEb2
H/k5dxYp/KIKf3ErZDsQ0oyZgkQnkOBZIVci4V9Inh2+vt/vkMSxVRsbf2t+JvMPQ9O21/R6l0d/
N/QJrusUSLErb0+hb9qdL5awlDvuPzyodTB9Iix+ualu/icGcTXkSp5WerxNt3EFEBckebYh5+Q0
Tbd4/BHMmAwvvluaSnJpwsDjdnSvBRkke3Ig5PBrE4Ot+5hWy6cTbLAfAzJdpaBISZhW5sFHz0OS
HwmDT6DYmilYScYV1tcbybsB3MXDCx/5muBY1FAcD1F3DajZ1rYgvtKPE/qdZWTPv5YXsdZRsYL9
u+evlJK9MomixdkqZWLbigU129+zxWH4LCVkbAcr8KQNd5D5gxwxIBdXTnYkkgtanCgTI6daOfH+
17W+pltXAJyLI7lksfmHVLkPm8uJXzLfDubh6kPNtrOsLBH1f15921Mg/e8ijlsx+qOgiW2Vdm6Y
Cn+a/Wmae2A/vDw4yHdltCv0UfOGDQxLQvZlOgQmRzkGyrhgHVBhrg7x5mqXp5vjUYKRZaJcQ6r6
3DPCDslqC1ShRuO/txuiX7eGbacKhJvmGxrx87L+4vB8Lad9AzxePewTN4w8YCGdLlYHtEuEFTWg
KTiqtKysapEuYy6EY70uS8nqoYKYjFMyOXgYEY4G5e2k48jeYXt5MQKuIuM7dYG9pAUbsHZKrg45
UYVr0tSsBBcBRElCetFU6KDAG2ENLeBgCWsUmUOrng43Rxaue1CvmtI5xkX/8fvqUFsN3I54uG0J
zMiZp+PgCJl//62kiWcMldMGH8DmdZCXyy6w8s9oIhzDai+wFyB1Xs0TkTdBPlJEO/CjwBG72FwS
Kc7JdTb7x0m6LSKUdYcw8V4D0PGgdRMkUXGcdpMU1EiD85LGzzq7pYB553DtCSjLfYv+P0ySXAQj
JO646J31jRUYqZ2HAj78F/gNqYeX5aVH+noBMa/mflJRx5I/BcyiePtrf7qNC5p2zy2sfVfycSJ8
u3Wdwhald/l5Jr2YsQ566GS/+zdP16Gb5ivnQUkqcWE6XaWr/KLZHq/RmcZmBEgkk4PN/oYpgNWU
9gNpvgPASUSCargJsc/RZ2Hl8TU3NBJ3H1z00VlA7q9fPHcqsNoGMSj95qpoyDGkGl0xbikpT3Zq
j6QHZmWxPlnYtfdGjTz1Rk1GwBudgqy0qN7l3f2GdxqC0T3QucxBrErnXOYF/2pItWvRk21EzxQH
509Y9yfDSZ+kZchiZ8DxE0xP5NSIa348zAzFIE9Xp/qe9RmAQw56Tvvp9ozwFjndYiSORncBLX03
IUcT+j0nc5h/xyP43lbfTnqPzJkSGU2vzAtaS2AmM51QHbh2tYOfgPQtfVxaaKGf4Oi/gMXKmmTN
89vcgxqsZFLn33G1mvKRldLDo2O8wDZGMbZ/Nj3vSHqIsV4NO4RHDb1BKJS+klv+6CJToQRcFh8f
eV5lU/xlTgYrxLfvVeI57nuZQqEMr+4ow7QR7KpBC6+eqinkPVrh/xvYNxjG27LA9KbsLSGVuVsd
1Fq6KTIyNst61H5gyoRJ/CR1uhKh5gTPDK+FC19v6p8oBuwNVoCZEd+wIeiCD5EO+2cdNyaGAcwy
HSyghmgNPUbrTFghNOLpN1z4U5aGiIpodJpgNpKONJh1WvCQ64djs7UzsKOkejwWfU4pUEuXUgqS
2+q/iVOgRDvi1SX3fh3+GjCOGFt26uGjbNcsN06ve6MiDnGsudZj83+123hq4tWbhzFiUv0IrHug
PyFxI+tVL7HgT5j2X4YJ0PiVq4T8LE2VmUoF35QGK+Qx5A4A6XBQIEAGrXlpv/xJ5OzQ+tcsKr0v
rLKnuVCHDjjKqTTmUTSDlvoyrCwPELXGyLrLr6G/GslIlokSBodQjz2buYvU+3hsMjdsB3CYy1z3
kOxSyltYohGSuSTWFV1nAubXXt4J63zVH0g4ZBf58tirr3O4iQ84muWiUcc91oqYWFasdZfxn0Nr
sKyyKadX8Ik4DvoOvKTJVUr5fObsw2z5fL3+ztCwH3hrXRyoM01s2m/YYCQS62MLoKv3ddWkYajl
JLcn1tNALMHz6Wjv4Io25taX3T0r1aLHvt1L0/vV4LflXZp0XnK24aLF5lKViH1duG3PZvXIGCZ5
8lt6eKKy1IUMWkPFv2OE2H8UbwRc+qJ8YpyHiu4KcxI5vL/hE9SsMjzNlDYNBU6Filiz8eSxw+8x
gWcptyeOEylMAE6m49DWoyeKmz2+3st8hiNgv2t2m/WyxFP8PEiBcr23+46xAje+PDZ5w4u45M6b
B75d2zSWvHvZmuE9MwWleRm3/jrAlAcmZrch6xo/Y4yIb5P4MMq41HoNGtHQJ9b2AqVQqI0dvaY6
PFH3QyxooLsmqcrZQN/ngmXEJYHK/sYqgzwsbSchK2jbRR6cqs+8dmrp/JmyDIyWLdrnKvs1ntYD
DHsMwZ1pSaTH/V45ligzWW9YO5ZgCj4SR43CQPp9AQVKQxk5OxN1xwb69/rDCzuTr6591bzwJh0H
O5X1GegR1PxJa0MYioRv9dwoga0tJwvAOkXIGkMxpS92/hI1XmNk+9ISZTk6HrnwKYCqa2OwM+6x
HymYMV673OF41nESEWP/KfXmk24b4hvaBXCk9pKozF9fxg8k66L6XAPxy59WQQ7ox+ErP2/PqHcZ
9SJFTEWUSwGpKVP+4MSSSkfc459Mp6efxyaz/Fr39669enn3OVIpQbAt4plIeJZnC7zVqXo9T/LU
DQ7D2ovvhjcxDmOCMAEUzP7kQ2HLsySHpFJIs+cImW4OfO4lzpFyBkD3WmZleFcjE9STHCD/L+dU
7Zfo99fJkPhOQKsZAP1xlRQGwcBM/+rcb+E0TsySQg5lXsieLXwOylUh46PDCpGEuR1LjLtA/ncl
TKyP2laHnsPmM+V7D18XG8sKOl/X5EPcIcVKO9dW1s/rxxIpfY9s2izl/PgoatLDrYt/slZatKct
oI37D+iD18yZ2N2Yy/tPUq47F1x8eCIvj/JYZY6mQoM+fCXI7/TQxyHzo51HgHrmzC+pZmmThp8g
TmXiARbEBQjlfusJojjwduSpBUmlY8yfCoyllS/IEg3yKYx2bkcL+gX691ZxupmtQiqKmsM2yuSX
8oYgFBOOkLI4zIt1srk/PokbaeTAqNV//LOwMh9rOBkgxwbwA7XHo6HhOibTMW4z6tw9m5XrAWsA
RElXKVLDdM1Wqu0iFKImURVxkBsO/PCKZOhoeJ+HlV9sa1TviKqk+l4N9RV4BTWsKNRTQUMIk/tZ
UOlDBz6nGBi2IAITGXXtTblkHvUDKvj+eSRYqb6yQiK3op/oFB65efZPBRQVJeo+anLxgdoFJp7l
sLFFJeViI7NRdzS3YZtkDVeRcKSY0vb8OTNqtEjWMbqM6xQM/Lp3CwnGvadgfHExbjL7YUqnSliF
9FJYqGT3PuAZ45GvZw35eVT+JgPGdhxwJ3Klev61jef5vr3tft8CSBU/bJOQNdDVLAcFNNq73v0M
10pFbcHwT0NuaCYfzhrMRHg+h/Gm3CLmjMW3Ri9T7glqYdbAyfPvCumdxuCY6EfScbUiz+Tqw4xG
+WfZ5T9sjyCcT4jRfYhZ0QCzFI+p2+rxljYtlgxLNxwNWZ4tb9nDhHZmYfQR34HkToIbCnQSolQB
5bMiRekUtMO+SwmKOS51Nce8RYy5hcJa8gux7cPyn91We+pEQhRcllEVSZrrtOLpeIHzk3qaLUJP
weWhW1TssKb8+NRkRnmyiYdjG+QF9giKieE90F55okzPzprIZqZeCRg4LbuZt8NBFltd7T2hB0Vy
YnTTIoso7m2J2j+rzSb2RybNs0v6QROP/5WTElsLLu95hLr1Jy39tovh42G6xIw2SQxKCB7zI5BD
a0XMhQYZKPAEDvG9Zx4aw5AQbLrdkfVPa6OR4xP3ZyC4R2ReD4Jarw7f6gMJ9KpgnVmk5kr4aXOa
eytn4VCiwUwAZwtTH8eVd3P1ttMIRdb/eWlXERbJMA/40Uyn5Mm5AxYOuAGWiw3O+NduOSPRxi3c
59eQCfPpK5Aw2rYQPyOoDgulrVdmV+fWKGocpyemIihczisbH0Jf8KYMhcFhTURWvOz6Uvd8WYpm
C2SFtS8FSThRDJdNcnrdBgNCoKb8BzKJ7if97dKqinm1x+AMsNcLEUHeZgXqfh5gjpX0E+MFsoe4
1fhte/YViSchMBg3+FaAtxqRAyJHgjjvwCtcriVUhjGlqM/9TnGJuz9kSfjtzpdS6vdHX0stvCaP
J1UK6VSfwW4bDhrsuW31PEm/licNhwGjMQkQzukdufRsIX5G0fDZtQhAR5t1XuhfQAppvawU/PCG
13NptORVfV3GopQu3VnpEgAlxSLZ43Stp5/Nr/29TIEiA9Um9FESwuYUlo8k+uMWSrJId3nIA9wD
wr2fJPyeI5HgyefDgGCZHi97ahrn9k9e4fDe6KME5huT1OR2sqTQLgsqDS+gX/1Hvuy094QVb/L+
hvojrC/kNgTOMn6YRZQ4Qy//rf9yBgr24Pa3/tA/uYHstr4cyqsq3+INwvBKskNZswHsZ+IMrbYJ
I7/53XMgU6SM6y4JjlbD5SWssRCGPKAUnUwEfmLopDCYbNRjRI7nakrZF+cN11HM4qdgZK704WqF
0ZlOhTe87g4AsaNzvkNSQPF9yMyfTfmRlGTZ27fs4vF76Zrsxbelfa0yJPHqNyw5JY0UY23dUe74
X684zo7JDnQr21zNyKJUOzJTCRIQmqTe9s1mFVXZgXY7lGv2VlGhIg7napeLlGeblRaYXyI26trf
hGg17riBke3s4W4PLUcM8D5kzMKBfFqheK+Tes/XTacBvDGJOGoAzqLHGmhvAS23QYnehXjtpFgh
16mRa595VN7b6d0kbQ0+2itvogw3Kbx8Zx8ebV0LC09SHFkVc9843xj+9njVuNUZCtYA+8Ry7QQM
E7f8j9Sl0cea0R8EAVYs7TTPNUiKuflhNNFVYD4pb0QKnFEnCHyP4TtYcQgHB5Ulxnfrc/4A9W9Z
XsCtO1Vw1T+rIlw5hMueTZvsGXq1vnw99TndU+CIomKQwRwnUudPKWPpjwq4Wsux1377biQunyHb
BC9jzHta4jCiWE8yH9LYYy2MurDRQY+t6o/H+dTXQbcq1ZW9tTC/Rr2pwz801UvE4s0vHXLkmk5+
eGbgz3g3jpdszGwqzt2SmhAILZm9PbHF+ld3Ycj0X/dtOTfSqsYgQr/hcZPqh7L6BBkuSYMhSI6Y
EOCOWFLcLNCjWMAlYrdLBEi268mN9g83s1tFimH1H1jBf+PC3SdXH9wcgV3mY//1hqnA2T7Ofb3S
3bvtHgRvQ/Z5iL5NTSuQSLqnMna6OevZ0Har2mgPn9rd6wx4sZ1JlsUXYo/r5soy6kOrcp6eZoWd
bsWEKP+5OreIRZgAD0EBLdRqcBojMsav5Z4wd87LCubIloXNZaNwzR5r7cDNkiQjNZw/xeso6puw
glPRrfbjDlpL2MC3Cm53JLHbxKSHNwJICCCuRdxcusy45Z2DUX0YIzBxyoIl8sl1e1aGHXg2nMVO
Zf/bO6vTSix/JLa88rfAhU1xyYceAFn/ekfVUlPVR57//GXMHxErP1gwKei03BOkBPDGmuFGU+SL
Sft9prPNf4FxwMLh8ySnB09yQI4bCFkN+S8F58BB1rfpVb3zzcsPCyZejNfvDy/a0y0hn4WUa9vm
azFglGmGMMk6wxvSXSzMdY7sWYmvr9f0lN2pWUHORHXnAcLr8ftNuy0ALLbUCxYK7ujP/g06AtfB
N7FrfLudFW6GvVrA/tNpXzFimlEa77wdEC2hYS7yaa0HpFOkjKk84HNQrVl/bMkoyhJPzJLfJi/Z
v6wy22g9G7ZClhNTLwjAzKIvvovEvlKjeyNCHMX9WFsO6TGOIEJKkF8GugHKS6dblYaOVLMk49tV
yTfXRL01Le4jEb9rU/BMXIOpHGKtF42BsdY7KSkfomtMjNtz8L8nwMeDPd46On4e6vxMQkOFgtpj
J4UHMoEEbfxNdfUVKuG1UpB6BLomGY63oPCIUbJzTJ3lW/gzvI41D2VkI5GRH06rOeGLPby7cVXU
5q+vNhZlT9gaem89doZXEJcpxIq/+hpStdZJG0gJvEmiQnsomz6RzP5qF+NGFi0CiUU9OXJaqJCl
VwaCHZFLqd85Fq1BSBBIadRqy3KwoC+j7eRViKydvEyEOA643oRFuPb5vOPSTGbGP3t5LTU4X1sz
SJlyJiM+U2vE3TlIOvQZ2q8jjrWNDdOcmnOQ2VRYqAm5ebak3Odv0ClbEqeebiCDyQR9VCvdwCrn
P1x2OQi/dyLfQjoc1tdp9Ticc86cNC+CxzfZL/z298gNSornKPQoh/RGvznVxlj4+EauwnB+y2KA
n9r+tiTkD+2+1HGf9nhNzfb6fmM5/pRljQSgJHw20E/zbT8mor/bF7MIL0ubz93xCEpTc1AIhImy
afnk1bcBaJP6HP0qoOxEt3y0eSMtu8FNdo4Ub2gbALvTZrvIKzmVD/7fK7R2+Cmjm9qGfLcp1n/6
s3hxF+uzq4ysk3EpFKbTitRzf0Hsm+BqORy0MZQ39kaOh93PXVn3HUxXY2kS76DvL2JZLvNa8Csw
5t/xTRRYCikiaZ8EwB63lnYGrpMj+j070gupSzKTPylHRojPtCKSkP6K7klED14zSFqFFHNRh8JL
VkSUPc10z9jUH8sT9aoshckfHxGpeft0gyanPpn97g2VvDEB0a26/TcCGc6QWYTLBfW9eA+dFwRA
ZZcyekANfAeVRDOu22yyMHygl10D+TEp9YUsjz2aoq4xdoQKCC8Z00gMr1CH53Kuktew5KuppRPk
Z8NVz1G1Dsg9Z6zlPsBHNY7z3T1XVTutNFUSbA2En0KmzNthOyAifAUUv89qN8zShzZ96IHwGAkx
fFhurroU8e28D+FVroNxRp03AJj8hu/9ceIVg2HECipN/Dhts+HBBqjbfMpnWtHynJF05R4/rE4S
2Q5z310TdQIqJeyDoUsc5pPGW1/8lKxnmEhuI16HCmze50+KQxXmKs9i+lRiCRGbBbqCkDjeXpo8
W2BLYbx/7SVKBylmZT2D3pgShTEPvkuw9s8rVrXJ4nfA86MU4VsgPRJYXGjSN0kup4AwhcSoUcAK
mr6E3tu7Pu4S21VVG1GPwLFjzaIku9QU4DFpzl1tXBRzVVjMlCx+0/fsOWTWw2rsGOegoouiFT4U
VZVmwfvYUe35ju/JFx/nb6W8+GHIcHWj5MLHBHJowc8tRs+gAXFyxW58UGNziIHB4V7ScpjV0KVX
YPFZ1Omos/YPCEM8+36nyXNi8kJA9KGjWPCU2DIE3k87uIWmefV1O1pa9YlC4o5u+JUvHqakPQD4
LDMINHpMUofAdX8hCardNxyT5gcH7dtxLvr9evQAfsrlYgemVTk+AN+GRKAZgyU5Q9w/Ku26bl3Q
5sZkWrgyLqGPJrQB7GcJLHwJZK1VStB3eoLZqW6m9Bf1fFcw8kjH7NylcN/GEV2h8OMCisOOyUMk
2KX0mAcC7qzLDngnqQquDqUkyYMyiUCzwGECpOvOwHyfyqnLxefdCXtWnE3dtbpJqdMq5P+ZVFrq
aQs/Gq6gH77fbOz4qtQpihsU50p0ODiI4gq4Vu4hV1VPC5no5sUvfklXwFzYnSdSHHaM33CcOaZd
advzhIfYm+POpnWUz1xWlUVqlZPkcic5k77YJb/aI6BwGftqkay3hMSS07qf3jIIGKBntX8r8kma
92+nFFNn6rxzqKR+WDLwQKTBvZYLV5IBtLeDqYeEQXlCHbApPNSJlz66lx+6zDquc3lNBnMHj2As
ERohQmQkrllxUxG9PaAvvI4hXx2GqYZFZq7HqRw4GMAHaJ/XHofIBzqg6pBc0zaRVMpUmCIe0lyq
ImlbN0QmUsxoy2uFEMJHvb1iQyHjUMb3Wty6vbHcAL3Wu5r3SfVXagti93/gcA3D/aPqneYJd4uc
KB7iwAcoSUJY7GWsGCjOsFriQCIjB8FlUYBrp25zfm+XCRKt5veqIQkYmohD26elTv3ywPTvxqJl
IAOU9q3TyAuGAQ8ZyCDua5wq01oR/yOC9E/6lVqP3P2uXU4BVnA/YtFnUZkkIGb+SlvdQfzezXtT
xNsOMmJaXpMjZShAtrLnJP0e+ifNaDWcDvpmnF/ItaZdgbyAjVPvU4U8vRdyYTHvozWs0jKw1L1g
5P6asO58pw17yZyGN4SLmnCGXAUu21+7p1ydgNrZ2h3b9I52HvXFyGqLbTs9EtEyylMGB9OYRhbq
8/R+nF35+wBWfHzF58QL2MrdesT/wSqUEBFR1nJMBnKn3UjNVmTiOW8ekJqd3x2XfR3TZQUXwVEU
3skGez5cvPMPxtFUfElWMZQhpGgPcJk2ZHBff7gqfYrEUkmneZwet5gOJYN4gvZ8baTPNQTdBcFN
6iuiEH7+Gb7wytNeCzsWbKAwEkgqmN/QufqQoZ0JTbcQ+aaDikpDwIdvL1aCWzE0EAKqnHa+g1me
95N7JG9MN3GJVkxk7JyeklrbyOGgCaO0FlUVelIi9BTcTQHDNiIB8YojP2UzPHzE5YCUuWXKCpLU
TsJBnmYY9kR33+vdbBoZDinIhMJ+JRnNeoQojTP493ngQUCgfaoojf6Nvdv5zppUY525c/KBcaPh
J/UYlN4qoWvjCrEk/fEQU3WtJv1dN8iIZ8kSlAjd8CKxhVPoHpRCFxVjWFtmeaJ42dESlSnsr0oP
wc3ZxVtO4vpXbJoQSXmaFomVpWeOtr7fboqINHTz1BUbELa4EDd8tedZflx5C36jXdhu2QRgVLmS
DF0Ew2/n7dFvlfNRdYbad60BV3NS23i+yscXmtGo0ZrX2+7notjn7qZg02V4NbA4B0mw8Lo7KFeV
0NNhainuoa7gkMXddgtzqA/4y1LPP3sL8BaZuWrsyDtfMMMDWYm+rUimX+c1/sqzuo6URdxmNQM9
kNr6IYOo3+6xI9r4Ga8vhdh2rXLPLyBoKZqqe8qcvpDUzyj3TWfiiKrV3kN9msSwSpCvMQ68vL/o
qE/JA57kTTH7q0cW4SFjlqo4suLbBaPd5mGoOuPiCd2/+iydaX1jBOJ1jLJPca9VAsZQ2rHrQJaD
x7PjwEqfMEXg1ftM14xoKMIourSCLcDtA7Gb3Sr3lSFJMtpF7opvYXGhs7OC+kyq5btnmiuFN3g4
evuok/jD00oJE9nJg/DqRh+m1tJnIt4x38WBvnsHM6RvAcIkO6tKBqze1HPlUNJH9fQY3aOR+dCF
eb4e+Iyn/nY8AmVDXyC5whuRWo0WI0XRQ9exqiCo30TGk15na+vqRyLiLic3GFM4hLOVWsxGdNLi
SiChAuqHiyoV66f3a+v6oN/Ojz7Fp5t4fSprIJKITaThM2JPQLfaHiKN545p5O0ybmxNWt8mkZG1
/mQBrzyMal+RZtCP4dLmo8JjtEWvSkWomW3R6t1pt6vAJJaZmbQyrkdjAbHu0tQh/UHe6mosFMDo
d4dEaIln/AVNFqofzlPbgLKeLDsz2CTt0NDRtbqiqiKoOIuDhwuwvSV7cIP8r6Tlgd5wcWmfrc3y
b4QNuELbPrWK3N/M0e8AQ7xBiLr9F4U+gYgsi6VnyCS9d0l1Ofc3r4oIkHbfaywQqeniA/0QJnNc
Yf8Wlv5XKL0rMHd4eNVdIJzWMieQjWBM+fndLMvuhCEMgiMRBWKVbyPkfcE6iSnMaAgj0AikwW+n
oHd1oTMGu05pKrecsZRQ2INTJCj2NEAYq8ovmkIGT0YXlRpIJxH9jrgBzAILoNLxuMgJ1pnVKLjK
Vm3q7Bo080HrddjKQQrlYFE8+8vkv++KegVAgKe1ennq8T6Q6lMriZFm8PZZMt4sAxPOhAGumpM5
TRq710qEBhguhpDWehPP6Ki41qmQ3pzwtQm9CH3M3Zn5bKwX7lppG/frcJfRbRQkdG5VWZyq6+J7
Syh3Pe7LS0uOod7LL5mZx726q+QYOZgg6qv41EXdGx0HQ1mEbnCnXquPhZ6VduC1Sq8kWswFmm3V
1F+qgsOAFo/YNFyHU+EB/5DGELZMpQFUGK6PKIp/6LqJD2CdxDlL2u01RzBtpO7PHgwVV/2vhGlI
nDYSBtdQWHzxdhvSybF1TzGS9qBf/9cDERf7W9vBK3OpbyUqHvLd8omtco2PbMAS9ECehF4so0m7
+oW9VtLFwn93uyO9AAkh1ppShlYwhYVxwcMg7ysABpMKbqBr2M2vojgPcyjjazmOf8uKm8Qi54Vy
0q+roOhhg0wUGkHeJ/BoDmQT4ThO1IBCOBWEa1gFCj5hOBj1iXGZy81U4Nec/8HYExw9Vv+CsCSP
SWx+JVs6n2nDwII1jsiJDGMSg0Pqo6ZIxm0yaLJQogG9mY/xQEsmOMJshK+S0DYKe9c+FK8rKzxv
ivt18m5H+7E8oInq7iIBTXzYKpHu9XH0/jpHdmzReraVJluGMKicqWF/RLj+ml6WK7M+fZyC2U59
kht6Vp2QODEbpgShYmgoJxalyF316oCOUXM7kw0a4UyFtszwWzJWWwUPa30W4riBHFjoC+JR0y3I
Th60zoxmuV7Wt8k4odZFqfM8AomiWCunOuphB9OmgbSLxCLWdQbGd2ZexFhsHfCgkZ1dCu+wsSoI
5Tn7IrKolUPNAIgPn6XAqo8qtE5b6EYysHK3JE59zE8XPZowqIYoPfYeo7Y2kDC+pIbTm1wpCiOO
hSGcWWbLCmME/Kz8xJ8fmrbxtiwi8BR1oTz/nczmUTCSIaRDQSZFQDGdqIsrydnHa51lY4m/c49X
lqeTlUxJGzLcJ0V9KwyJI1hr72uWT17xDOLLwb/RKMBKOZdSlC32bvhoPVMg/qAVenZBWP64y7MR
gJIwwTAjQudUv7c3zSiblWpXLubhPSdgi59dp1Frx3fSxDhflak0Xn91RGypjFExcKXr1NhwdXTZ
jsJmoSV2fglblxYws7V9amO6fFBGg4YKUeW2CBlbXHs4CDRBmVVohu7V7Jzc9UUVPyAu3BdHgncJ
6XeS4ZTmWW1hScF9nMglx6VLr9NRdERlDuR8R+f0QmWti/7vfirNf7oHwqNdFkzGa2vEuvfCD9wc
2dECxatNZyPGe756SIugF/Jaugp1tRRg/OZAwUuNOrI72oGOKvVIWUvYXUTFNd7N9bDvvNn+kEOX
YbQbf/xt2Ynkg9vuO4p+6OBuSSecSkaSaIlX2sLlJ0lAU4rE/Gno0Hy8XTo0HcM8s7vhoZmE+KFi
whm9hDbdnTE0km1C0qb617qEHtNKsa2nGfJpDmkx1dbOiUSMvAX0GWx+6DV3zNOqJCIukCbKVB/z
w/s+Rb8hVyUqwabuuH633JURChipPdsFv02t2MLEJY4wFODy+97p1U6ws6wZhUnWzBFDLRDI+Td0
pkcsS+eVbSKuqUlSkVGzc8ti5+qiUMreW++3uRnqjtL4rJDTVr1fBI0a7RqAZ+2Ha0m4tAOS7vME
v9AeOhioG3J2g8aw4ofnC8SgPxw/tRWVeSKlYqgU41FKHfGHywa0PnQUb5BgtmRu7Thm2KWRrP8w
CbsOpzBgbdfSHj4WtAlY8JyS+2mfHKt8m6MuqI4nooO9bTvFs2j+FZRZpwMfZ9m8o7u4QgV1tiuq
WRHGYRMpkftPuczRfVy+1i3CfAnQwP2PBvWnWebaQYkBFF6D0HqrLzZKrJrvU8forViA1GIOccy8
nyCNBbs9Kzqg6ex8Voq6SnpmjZH/YuHxR6k/qq818VHZnNrmtgysaEum6Q/ZkGeGUHZFXkAtsL+r
MshGRdLSXERNNqkPpsP7x1fE2aawbjxah0lAjfZw5pvD1cabTlBwQ0Ex3BvpGMsM22HZP12IZ0zK
sVZ43JPgQnRmBn4R3EE2rINVc9g41BylEdQl2CPkyCYT+Qbr6EZWJ9ftJi/2gvc61HgNSOWO9S6F
tslfirE9rBTjTuvOdF7I4lYkBLqID+12xHsJm2evmwCn+HMz9LElMdJNem78bx+HYffWmn8cIDZu
PBFkes+1DyH+VVl8NJ2YsuLJuGkVopdO7k7efM5vUv/WRYmf7fLo79JffF1MCAZVCRG6IfnPEvY8
MQHZo2FgCt2+fK5C3zr3wlmd71wcUKaPg1UQG6Cq2YLqloOoCBJgYf1p+BGfFpMRS01Uy+Pmazy/
cfmKOYHsVEorn/SEyr27m81Om6EtkYn4hqRYuB94GAEF12d1Y96oU3djYmTsMHys8D9tsC6jZZ30
9SHk6T5SDps3eI4migga1vfdi30pMxqRYHL8DIEzCKZ93ZYQCIalTPJnFj64OYRaEVlPYeLguXUP
jw+FXfGED1GC/tqtUpyKyH9us8Lsdga44N10CNMuv0BSGva1jelX/ut15X9i7aJSWddw3uPOXZi2
1NhQrzqEa/HP6vbUhlTKLsBnh/D82p8A+O1P47l5CQX5NIxNZ/2TaUnKZ30WNz9cOT+75T/pOcBX
+UGRVyO6M4XCQYiLYGPenkITNYgzSolTWMxktqPa4lgknQ15OYK3KAGRZObLZSKGGuPnVGSNtYVv
gU0VAaAujv9YIaz/QPhVzu4RvC+sSKBMysS3wlrPBpl0ccPPrVCDmF924oTBq/tQaIrV25nCwq1P
2ThhiTtRDv88sS+ovVYYdmHpgUyrc0LG0otvkWn0hD4ZMFkY+7D/OSflaP8/3np/PuRN+Nihaa7C
JcbWIFMW3C7jpiTBFGtxufCARK/tqajaS66Ct+nUCXtCd0aXpQdoZt5hVrZF8y2MuiPa2NW3fQW8
ayYjYbur+7F43KW5Bu8GKYuXelJV1+RCcvzdWXXhgR5O9+mNA4hHvZC0UgJEdKr0Wu6yoQDTdzLi
C8a7PplyeyB2s7rJfsWxRdZw84PGstyHw6DhCKnuGRUhWa8ro5UTaZo0e5UJ79zYrvf19U4bc2uk
g9XD0FBi6u0gynibN+RJoQWk5Ykc4s6HWfgfHLY25q8qdo7WeRIgm2PnwT1jwfktUFFalm3tVYVy
8jArak60SJkGQXeE2nUq8js1aH4go1eqBzA/MEb+V7s3MfxBIK4MshEsljHy1C0brSs/b1Q8ZqVK
7044ayETxVwwnGvr4C3I3c7lWjCLHZHxYt6jZItg/iUX/fXlbGYN6QeUknlnmssFps399SRNQ9ha
2jjNeTrFywmwofqkhAMGC3zgV5jA3nP9qTXyZADhIriF+ba5nzKRA/AJ63fw/GwCYN1LjLm8LDS+
D0TkUarOfg/DY5FGNrtwRF6usfefo4WYsO7vwuHi03AOsa+Y8bvdiXDgHuR8QvscWYVIJ1JzcvvL
vxb1CEzjbKGZksbdBj94oQhz1+USuBsj2zV4M1FdxFLm6IxAL/n9vEUvbCSuMWGsMuRBjHocjgxL
xP/Pr4fTYUtFBLbrvsNwV1n/BaIEFpcpUmldVAA44SJPQwTdJWDdn6vKoF6puf/Le8QDGczL/rJ6
KOPSqf/Zgn8CmANWxDZ7E7TZXW34cvmnM91dtg+mcPfbULUD4VEd85KHbMB8Nm9SlzjO2xpZqVpz
3G2XMyhBGJZBuvBSr1X04pAcDpUHAEro38ogAabKH6EHBauieuGG9QbxPu0A8mLZSKAFnHKgXlv2
+lxWgEBirEQUh/t4v8C/jZBXy7lMaUlW98kVXwiR++czRYC+vdyFya3ZQlAEmRLwo2609SEhEpI+
DBfNL4xA8SCrK6VgYiVGWUm6VtoWiB5Z3mzTJcIKvhEUlJADvhQDT/GiHV0mdqrwiYRpJRJemk23
VBT4DbLoh2OxiVHR3qMx8/cmZyEs9aMCt1ctfJn3rGyhRa9aFIt9Vo1Za2r9iklMJCPRz/rzP+sz
tVBn4ketCdJYZbZU46XGofkj2hxPUCJzrh8MiIPyZ1y1y1A0sdeCcpcS8NW2pRn6gi2KeTFVNpn5
rYzjt1kRZXoS5TK6sdIKpWCMd6a7ELtYHO6VTVS631oyVFAsDd80zsEG9JuWKQk1dHXXtLCwwHv8
+A+3M6HTHDtMeBGTwC8Jb0ZmwRgabgVgQiD4D9uuDP2brI2dIttcBvGYC/mJ7GcRGkNyZm3V9rIE
uGJHi/7l56vvj+cXPi7uxuKMZyFyPG3RsvzMqQqsth0uNuDezerdiIBrFWQX+hSFEU5pg/5dCVxt
mt5gzSL/QfopQZ3sEgRnYR9wqYsyika1Aya++8YjULczuCh+o3xWaf75D2ZR0G7NdfkUksfyo1Ei
d0B0O/DQ0a555T1TeVsVTcaHCdOvUg8i4xc6Imi3NYbD82IWC5geAAi3k2xX5qzhUNtGbQm5oMgc
URGlE50/ZooL4eekrzTkcOobftSr7QgM+WKfyhjj2Mc6yTIzPr6n/5o/IMF51oGlKBGBH2/yXmgy
B3CpDxjoYnj0Vrp6f2/uaoPdL+PVnnrmOU9GVL2AartjFRW9DPB6ochzrWdgA/Nqx0KbPD6ug3BK
W98fFotWstTIgxfxqP7kfu0c8ClVpVOnn3s/qlg6aPV3soA5kUxu/XGz0UQCzoAmJPmBweA1uAQQ
0+oxmBE3WZqY/iUqM2pMtBT88fT0oCzLD5g7qRWeiUqoFV/uRrg5eB+DyyJahT31V/R02uMcd4du
UrA3JcpYHOAqMZKh346DgWajBxBZupNc7SX7G8oYNaGBT4RxVcUs9q9c58A/84NaEJvJk4moVc7q
tToLT+Ig2LWw8w7rOqgyeM7ku896I/LIDFyDK97gHOBH8904KTa8BtLGk4Y/U0/UBEkm9brm++Et
UkR1hXPzRYFAw/qhiCuMW2KhaJYfGBL97pF9eiJVaaRz/YNZwxk6YN6TlJIzJR4NN5a+gjV2orvB
nhf2oqwIVSlHv5S7Ej0deYM5OW11wfmxEeJmB7FkkdJveosN+vHUnYKf+EOLZGHoLmtb8SU/HKSB
iNTTBUQ4rl9JpER9mwi578EeKarvX9n+JrXrXOGzyjxvdHiurE/VpDiXuKu3pvEf86Eg3+Jbm+Mo
UGzvqRafv6n+tBqK/7GwPzkXlOHhc1BRCCH1XDdJqCIMa5HwT8mNkIf3u2HodstdkJ1F/NHgaday
03IVPpfjC0rFYZ2sacu4TZoT8aUDy9fCIp/Q/pxZHKzooHfqsi1huDR7JZTYGhlFU/9b7p96WMDc
1WF3P1JtNiUVCJSOVtiCmsl16l5peYCDcplrGeaexIrpsiZqEA9nAKVsx0FrPwvZJ+jiUxyNwrrX
MzY5JcsFIyXIM/i68iLortv1baLmLB1R15f+Ge/D8gz3l73lnog/u54CgrHu5avCKdCU7e+GEpnK
1g7M+s03A46HWYLS/o22m3U1Zcqsg6DqdTFNFByJeeG+KwyybOaCwlq0Fh4TNwMHeeHClUb3ubDG
xJ4hOt1uK+0INN3C9OLW8apK9UjFHty9sWT7077zw1zTzhRPdw3I8IXkShunPPxFy3v+3hBZ+Y0r
4MCCQ9oEHbf6S/Ea7esiRCYJX72X5PhyCHZM8naKBXQa1bEaRn34a4cxoTztlPoycbV01MAjc6zy
JsJ1nmsvZJ1AgeS8QZZIAsyFCsqvhE6a1ArUjMNmayTp2hg/vbQrCretImPn1QTWyHvJkIyDG0dR
Q4ISJFBTBI8/PsxM+dX46WiLnl9rXeYAE4rmepnbSK8YUznm85wVngDAumYMM5p1b7te9vSyWN+p
jKDc9/TU2qJ1DgPyoC3EnoZHamhLMMIMMvtAepmK05mcV/6Q/m5zXzHNdefZ0NESiYpsFvehV6nf
6E7kL4K9cJzKouWfxKq8cLffLVvisAVt5XbCxdRLoRssKxyZaCAhNcKeSo8W5rP2OTsZsBv2RPdj
P4GuRDm3qsBxjsz/IRhT/FWFVkZ4tZvJA79nfwpewsBCqOKh3XY2nRnkfMX89TA0hy2jqTq9GMeH
nNFCgwrrnx04XS6x9npF9jR1VkFzrgx+Pbn7U7TtsSyyqRviWLO7YhZWwtkCQlHn7FHOanw8rcrf
nqnOvF1TyYHLapIQj6ou6hd6cP9wI5/KJS91Rrn2iU9HeuI46pqG0a0aj8TiFIT5o3FdBfYhV3j1
kBluO59CfANuiSf+2cMSArooESKdTEprfLjBuFbjpxQJ0pgc8wqJ9d9GVi1hCuNRMXt4mLAFt3eA
vV7XIUFYYae7DJ0LfFNI4ycN/OkSG/XEG/HqcWdhAIBO14RoGWdpiKjA/Itkfr4Rif66/vKsTfHd
/aZE93tpTs4r0sld1/XLNBPfaur9TyXdr62Rhe1cEhPgNv0ZBYXO7mBgkqhdpiXGEeBB9/lkMD/c
A1azxqwrVRc1a4AtE6UmhHo1HAJ7orwm/OKEKZuLBh1XppBvAEo80Bgs5lYQpcNJ9b7dL1HBcZUu
Z7diEx8S7ebrA6MQQMwjEQbzZKKT5WiU4aIVERfllRcWhiJfhwtYcdIXFVeg6l8Y/WsVKpYQEFWS
sXPAV1t8nc2j0oNZGQ9f8VNN8TBIozlA+IFRAt2ESOl6xuvZeLguHoSwWqkFSiIG5PUmXADG+yql
RY7SwtSQCWydPAvwR9e4kgfbfNjWmUV+0SRdxbSrWNgmzx0D2nohugZWYGtqk+C7YcAbAi2uzv0+
3cytFpqyAHUJ9i8kpHza6LWOMY8rkX4A0oZ+uvTWrO314s8TJW8OLoByM398sEEOivveYr6UyLyH
N20Xg0MbbWFYFualmhWbUGk5UGM4OneRUfF8XYQvKA4H0LzRQnCTaHqn/GrQYIsyjyFr8xYvsz84
bDNYJZJNiw5Me6hHI0bC1R2A/Qa14sPoJXL+c9orCLrD0rpiUznwy2bYi/8QIIca/+DHnMq1G5g4
+w6wqUv4Wqf6w71IOYz4bXgSyBrRG8nsp+APuXXGbM/FSOEs4v3EDwtwVSBuVSAYgUGnKQIEXiY4
tFnw9Mjzkl8CHUPNT1RxJZO60Yj2wSdxrOWGNBIPlvBOcqBe7/Va5qmD7KQLY9lO+wp/NXl99DG4
Upl8vrA01+KomC52AhtsaGuLj1QltqvyHzR9/vgzv3ALb7SIoB8JbRluDzwRsiQ4DdfPf9jn/yux
LU1NyxHTmgb8P9Gylh2zwiRInkfOupZK2LrRYnqQrp8Bxtr7dSd4dREwVOWTDj3Rh3wjR7dhJPPd
RZzgdgL1niCgpL77Iyhoil+UXQdLPcbkrBbhjFJAKjSMprE2QjhG0vertxClz6Ah51BiVPQ7aWgo
Wgq+gALdCkhYg46ooB7QpjUxKbs/EtuSKhhFB63gUDirFFoeU8IOvrZsddAtEGcQxfvOK67VRTWf
kxMthxdNpoQVocdyqFeD0D3i/kszjYPU4HIsPi4Zqld/PszJWn/y5wHJCzdTozwWr/vyB4WlVkk2
EChGP8XDQkGBfjW9WLh4obU4vVZPbG2z3nzMRN9dtUrK3J6bKcYQ7DU+KcNSo6BuQ9PsS3d2VZrj
G3xho1R/OHWe7vg8DGO7tIxGuRD3Jh2dEi7/wi6r1A/RNJQjTQLpD8TgUlJ3FpT/23a09EhUjx/f
UxilzgzlJ4Gib7WZ1hjipLf6FqZJTO+dUTmyTi/YaZi+uRLfQ3KWECR4NQOnHiJ7/k5Eowny57AF
AUTy+LTy1XZVqeb/bbqI/hXUzd1UhqVmx5HUcZnQU3tn+EfJU+9b9QlXL4pC3uPgNXTzXrhnqV+T
8qqYrcwb2C/sX3EdmvviCsonT4cKebLAepKbw9oA+8kEVr2m2gThXLbiRf7G+2iatI4L2Dn/n3mQ
4YeSf6ARaL2O5u0z1U0kShzmCWPVl4WOwpdUWgS66AZBTmktC+78kB5GpqJrC5sH5OfoSQOQDZBv
Ed3Yp5H34T81DLUIPOZ8f7HqWwwtZRYaF9VmlBaBgVJFcsbQN5KeZjhQZlv7E+cOrJ7TD85/95gg
LGZfMDNh7cbttPZ8DUotYdWDSnNGQVoboQwbVB5sDlj9JO0DNzzbQFo1eCeFq/xg5J/qPRxgA3ZG
Ga0KA/NhZ/gv4saoqovyx7WDweCoBSJecrP4J5q/bPx3ptVF/CpOtyGyXwEJrHYMdxezYiDhKmnm
h+vaWCNTIerMp6j8gwKRFkr5dN8hIKCWR3oOKtCzlfwJjbvsllA0mYBdPqFPDPe5v57IP3/AuTvP
ZVDt26580+oQ4oxrKi8w+IoyDoXcpV2NSQc2sp5Jkhdn6UkxA2hTOPAtLoKxyiL9UwcKetGCGaTS
n8eiF5kRICkUY1YlrfrqR4XU0zHUll1xd+7i65N2KolztHbQwwb4kQL3MyCLzq/CluXvt4i9y21E
CqkSOsH4FTfoPmOZLYJmSS7R5s3BbcWf4DYzUicbzGmdxF3iGhV2aOjCvnP0unXCePewKlky2g8v
3VIrZc27gp6YqW8c45+944g5MPp8ZVQraHYPmMWtHEqi7JkvYT8R9zHoDVehAWlwXfz3vM7PrywX
yZ9uzY8ufV0Z/TCNonpmojM2W6PQu1mA1CpWTkfV5Qa3Yw2WnTdAEudkQ52txu8szeMpS0qi1pJv
lSoHDD+o7OZ+329uOgwIVqs4HpuGXS1ul55Yt3byDp30rbKsnweuB8l+RrVwMsV8CWmJnmgJlT2d
6i6qbYm/5tGV0EbZLGV6w6bp4+ErDPZ6B0G+1lCDYvEjCN3haBVmp02mW7nYjjVwEwve6p6OjWRD
aZckmL0XSENPhv8nLM9YzdE7dLxR3NBZ2QqZMFQgaXc2NxMEsg3bp8dTo67aRZ160l2he8mVhEVo
Vqsq9370SyEJBlC1k0yDrgROG/g40NJWN6Z0/Kpa1yAdjH9D+Vsc3FmaC+pABjKAgX3nZ7jEp35s
MgL5vML7pcWXaa3WAVzcZm7vcL/Wn/sN3k3QLULtMFPbv2u73eUggS3icjmTZBLzPb/hl1S4xU79
McdcvUMUwwb2zfyczWymkN9zd0vfIQg3P/7bn6bvAwpEmVxhBgZ+Ei9YOq3lWPbVtX/YIhavqdi/
64BaB1uFHQGpbJI84AA10Y5KzxQQgITASD8RZslgNdPZSAayJT6mx9Q61tJKVQCSlEsraDWftBhZ
xyNG9D4Z/b7l/hPkAoDs1Ri4zVlgWmexgd62Oh2SzPPSUxSa/Nt8badlCD0RLPtJuESfwA8Xq+xa
bGcrwTNVLw+MarDlpsB5mkRd9w3agmrXpLu93W9IV6vM+1toYe9DmSt/q8McJgCnVHbAxKxxZhvD
XPVnUVoCVIgfWEG40Oj+xtLjxHKichjiy2wcmjCHHvHsq3XM//+ZpFQwueievx1vQpFcPKyu4xUp
0+Gk9oExwbRmRPVNITM8aciY2cRcxtxsMxUCapfBwuNMe56R7J4nOaED1INgLutzRu0Yc/ZVo7tl
XjW/pURW67OBH6NKkbe07TU7+t8lS7Er6MRIoUqf3+PHCrkFBdX28ZSi3kNheUIZfDnO2bGyMIKx
2OvlXwF3Jr6MYaCWFj2pEiqDVY98YTA/MbIeYxZqYEHo3SEjGzfghXhkwim8MNU3cQSKUHQ7R3nz
KI3q7FEfJGZeYXDMMB5/5ScVM+I6DMEzNkBSmMzxPLIQiXr+GWIBt/m9jLQRCs4PKuJPDew4Bk7T
D37UUrFONm9IHk6HTyQL7/8FES66wq2AiLO4pzhdg5FWeWAOLH5ibg6hFPSi2tt9eWqiZdsVltJi
GigqkMXwHpr6BkZmROguEFbE6eFmVvWJu5VQ5n15sXOTQubhx9lzfaY6N4kU7nKODdoPqhtaVXXt
/Vel4UeHN9FugL+bbFcv0oOeTNBCod6EkUWIY1ZtVTis18475dQ8fVw0sEvarL3b5hdPCffPc2v9
rJCsNJYUl8qoEUAI+JhYO/RC3Od8btQ+RMm5l/1shnxsm1YeFTzwrSw2BNNnPAaW5BLoqyYzH1uD
1pFRKxJDz0lgf4EBBfkMqJGgJlr99c4ahOYjzwLZdUO6n+kGjKG7kftNDRX3icPRChrnCO8CgI7K
OtnYQIWfzNVbG/TcTpDqcBMCTblJt/seXMKrol69CUPld59JA/JEbcTdrfydNED1kouEM4yXap6e
jg82h/SQrXi7fSpovaQSgFf7NYJZNcUjGKIP3Z2KCA1Yiop/1NW9uCcCGXiBViSLwzygClqs/wDW
07msdIFkNshHmcEKkyYo/6RIxAtl94l9VXAeKy91ALIU7dPCGC8LArGbTuRpEwfclAkPtwQgH/gS
eY/QocBHazuQszwHHA1T2glShN+6Tpk388NhjwnPxpwRC0In5IcKG82UIqq4SfANruVCWFiymc2M
hVRHfOvWfXHaeQhuebXPL8jPBswL3IYv9d6R8reSzx7h3MaAXZpkvb+hp1nMwI+MaLizRRxuKh0x
+HNact7N3qSu7zpP3UQU/Xm30OVo9qQd4a5tJO+VawhuGGV5QOSiVQoPHCNoy49GKn5x7RvbC3jV
wo9bVLJ29Lf5a8Njv7iGe7TyUpdzMju+DGCkZKNo9kiNB2Bi8Hb6H5h6P3p0Gp5eFe6KjwoBd61i
aHP2hAlGqkUDwOti3GDr0EMidUH+RFDRsEE1fSY2flhJCAQoxn1EfptSfAXXp+YIZIwVqgkp4vrH
++2KY5t9aWUKmx+VADwu1m2I+I8ifMJpLhFYhzEGBtJmD4/pjtUKjox+0YBrWmU3khTcQuG3Px6Z
ta8THOpc3fG8DST+MR07RYyriLHlgM4zReWfJWpDQVUTilf6CERrG3Kea0Qxt7EPwOTmz7qxhiTB
wQSj7LOgykauJqImOoQWGNriZ6cLsMlVeZ7LUsA8H2CFYLC88Fync/91B2K8E7UM1SJHDBBnFpL2
XX+pZrNLkrNjhxuyc2WKiHokv+6TMJ4Rsa71LZXybp1iiz0tODyzSJxMloMC5jTxwZ2p/IMDA8el
7IWyee42yBr7deA4GJW6dHhJoYmm/tKo3skYhMs/y3xONt6ZhIal5BozansVGlf19By1jArIZoWS
cv6Ycl+JmKXSQ1oBC2s8TU25MQRQM7q1CsfuFUAl0BWYvwNR0lfky3pWLn0vdQAj5Nyej7bz7eFw
HF8da9fi2MP/Xo7XpmFTduMEE7OMzwRKCnRd9vGFv6IQO2Lg3eLfeLX/KQ5lAJRoJN8/kkVyvXq8
3wYtWp22EafyNt+Ca2IWPxKvfLgDeaSBvoJuKxW32c9T07n9juAbzUJn6MyEG6gnga8TvpfJthni
W2qdvYiuezzBR4dppp1iju4Tv1IokXTABY4d4NJlg2tNt7E8cYoHLNa99ZjS9bIwAsj+qpa/HrJX
25SA4Sbjjla8MJNkFJuG+dlNqbWdme1I7RCMlog9o17GRb33G/LAhNmB86IUNtn3Z20cGni4f8pb
++689OwKXFeMAQyORPuFOo74W+VXbunCLOspHVLd15OngXdYXCMWORt0ukMNQ06sFtUm1Yw2Oe5R
2rCZyIRq1qFjaFK4m2YHZgmpLMhBPUriYLvNwDAHItAqbO2E57yU3lbjZ4LGc4TPpV1KgQWXlgkF
MRUS1c5PVVDxxImcEf395ahhDB4E88ZA+ekjg8RihLHudY3GG7SEVEbhDsvlDlMdlQzrGtiDgIl9
YBhY9OgKFMroFMBtdBPxSEL/Vselyo3bxOA4NN2pD8VMRUZTooAVJiq0arz0gTrtuUcqcSpJto2/
+z8Q+xAmpzaJ49P+QJ9fkqeRRP/UoYsfGe2nBw4igJOn81yBxWGhpZC7HTb8YHw19RrcAjutEumF
zUX2vbxqNIVdQWNDqZAM/A/PZwe4DbvselRprwqSiYNT99jJfSF3C9xAvirg8r3mkNmS1lPQBw7w
6gXSjx4md6gFXxkxFGHyasjPceUAomuXbTDJfyqsglqRDIMXoaPvfo4w8i4o11CAuQmFxMaPJ2vH
EkwSWfrkFuM7iJtZRYTfhdGHXp2kGaQA3uA/bOl4SXl3W0ZLiiuW4JwyIxM5yiehoQ/GRUDlYZmY
rLAgyZ3sdNXJT3wkEXfsl9mpbrltIEHcygsB0vX+T/LPz4zD4AOjiL76GFamCJwQcvTdbUp83NhW
HRttaB4WNNvIhH2Bwh6r3j/CFSdf514JzhFbYCiv9SeT6oHgwg0ubAogvXzXrW5H2eQCXQHTGlAH
wOKVKQCOPJ587P7e2P8ZwR+DykhhgH/k31Pz+rx0/6Rnn62ZbKZgOQbs1FGQtDmZr2m+hAxrhBW7
iPJCfZhlqilvtzn5jBRzytZQ9uJOCjhh3kv7YayfNvF9sUZ2HiY1xRvo1IcaWXid2OMep3mvnSFi
SQltzeWcEqLeDZImj8C/hecdvqG2iaBkMPj/MGbWc1AiqMuIH3aMd77d+NiCkX3UGuSLxI39UO57
gd66ieN3+DXLfAEDSni4aytvTwM9q6DNT9o0GIJ8UZDBD6wyz2GdxCiQDIybe9VX9RJQyUgtY6On
0yG9A0qUwCaTb5UTXMYQVA2LQRPDIyyYp76I7bpV6qQw2BBtm2B/UzB/M5PJNVC+8DryaddL69Vq
RSI5Ph/I44AlvsLeWRtsbh5ZtErwjeSRshWD7/PLe/j2Zy6wfmOtvDKWud+JuOK234HpfjEMMvTE
DmAm+TpzDRvwz9b5ThKHpossTd9k1yq73Cfal+RcXVy/JvhwWPj2w9ujFlDv1Y6ytssd2RHCL8Gu
bwnq/Zh8ofKmAjldhK7tLF5OQXWVxVzvmmItgZQ9/hHTLDkjrWWVPRE3DmVIIUBpCd3PXkBulEVX
IWGSLr5Vbgx4gidf/VYOg0vHicw9X5E1StP+MI48q/Ho0ur20N812m6u19CmsaVspVYOlue02C0b
yIKynOPXQD+I+H/Eh/uzJeJvf5wDXB+MLV8wmK0+RDvNJLYx+pFZMBV+wP0I3t3tBG69WJjGp0CX
nlRfSVuCjfAcQUpsvf/cUBTPZFPQ8GamtGRpDPq2UewFQzqygJTUdNNbCXS3yi+NzclJb/nEPSXx
+GUVVwGFswUwYWu42fLIYttkWFUiYth+gDRK6f2ShmsKaFVlLgu9e7a2o3KdULSJ8dlKPRIkjpG8
HfMBPmO+p6mr4kc2ndwTIaybjx3TC8Uxm/meg9UokTrAXPi3YOUnBkuml5q95CIypDvhUvSf3Rpo
ReDfNZBOR8AfMvLgULOjDIo8M913ZdmAlA2dxjOcwmFlahs7i/4rGEPpszTH7TQePI7cHLm9Vxzy
KiZIsrkrBOu9BTCcM4/M0zSEQkqNa19DfgoBGBKVknt1fzzD1jlUxJHbfVwwqPPi8GSmXdPwNEXt
KcPGCvozSlC+VKb7wOmo484i+XADcy8GfYRlyaz1xfwsIzPin3WG2WHDz7piQERQytrg5KQohpEc
LJJcPFxbwq2zybojFJ4EfJsPdrfep0SmwTbCQHn7ZQNHDP23sGbzjc+lvnkosPLHfrnR5tPDPgha
mP9ssIOgcAz2EKe3jt1elBTqCiWJKgCPsz0CUgGZ6YW8TneEGViNUO/1r2lXuc8uxiu/nHWQXwne
8Z3V98QcVJgRPVwRM6tS/QY5AFc9UMjfAH3tyLtzrs9CA+YlcmvpiE37el1IRvLPnYITVJVbIQ25
tTcYwPqpjJ1bilPdDscHs1PqW9ztTe59MZ8v4/Ctnz7TsglJrIqOs1e+1danS4RSQbjpaeSw+FsV
TGbOrxi0Xiq+bGljw+qQZZLUV6VBkMTd/skwgA8u3qoZSVb1EmEXs+R5yKjLtCGmOe5Auf2wiYdd
bZJMTSf1IajIuC+025zF0BAxXbfS5RrvLSPia4PoQFvX3EqtEcSzsgZZpNU5dcKcNCiGGLDlA84L
jfZr//nSOk9m4+SWVKIxongl4r3NXH4YFacqduw7EODSJS9I5n3ff7GwAebj4lEqOiDabgEFF1eu
y8be8CYfnCWrGDHTjetOFcvwxJK/4jbPUj9W5nNk6XNwbcirgBnhS6ZOcH8QYK4pQ9hRjvGWo4b9
dzbkjrScY6ihgbbbbVFaQ9rdmP5l/FwynDCFDIedkXAnLr4pE8DU1nLUl3j90CKerkJq4QXHdTLt
5dQ4eKUwikYZsCGypkPwqNzA0nsrzmCui/sB9YYLD78Bo2XeZNZRV0tbuevY5m8kwzv5S3YHnh+i
i26K2PyiBRY4/WfpkE4hUBT37ppb76pXh7uiwlTXpw4XtCAyTSuy3OsVgZEmFH7LYe+UNY4w3txc
DOowp6tNIem1CzQ/GqDZhewhWxSjj6JIcKrqoO7MoufHJqWCqqYlqBZmCWcEOihfYqrOSYi73cTJ
FgTX/dGllh6bd9oDoTX9fOxG91TPziDrrh5e7xC4q4vQeGEFj/WwfL3NjWC1IXoV05UJ68BlXz6s
MklFwTb5SYAKH+eLyDIX2pHgt4nxXHsdtffyqgWFuXYwgMlq5aDIH9RcCUzbgwiGc7tsoWu91DE8
rSQM4dNs8r3M7AoDdzcGB8WFtBOvbjJVYCYJM6p5KoXvLwx8yoiODGlqA1m50g+Ow2Wlw117JVcZ
eUfYSj1GUeHmzNcTk2WlhtJsX3webwXjHN1QMYSSnZUIpgH4j0q9QTwqBnuenryoozHNNBrlF+GZ
NXQiKX+TVGbisTAepySjtdKAgFIy4TodX/kgxWMhwWdTmfeoRVKG42XFqqiNzcb4kN0mbkYj+mJQ
OuMq9Il3L8Z4aw+g3VkPl7VOs3vZg3x9ZNjkV+/7fFChcr1kx0M35mkC1wastH/S1GdkPLei/rSf
+b7wf9oJbkXWJJgxSDyzQaj+0s3LthYl63TanH1ecGnlwjBqhG6dDelHriwBBvFD1lcEnJiFZnlt
8ApiqBadCPXBrmwN/rIYPpYWfZ+sTMRwxudiFON+nfoVILEDFkk6VP6LixqMk15t8faC9o0hH3Bp
K+7CFE2Kd/CeDmX/5rq9X+WVHwtEl6p5uv1IviUviF3D8n8rzDHsy7y4ZltkIpQ8rWSDsdiYfmN+
RwIgAhhaZAzgtZjn9I57bNuM14Lz2YCGtDt9M+8qq9ybtFOqMVxkOaoWS9XRwrysBBWf+XRliVH2
iLImj5ccqEz2RVPECrDN1kaur92I0KekhhRnZqM9I0aQNbgY0N0q/tbGKAWMBePclSk5YYb6RB3m
QHTmoszvzUPSmPXzb9hgUH8aM0AkeWGdiOhemjnQnSnK+LR/Fbsp4QBrq8od2Fs2Yw4qGcfV2nn6
H3/4EbalqPNb4PQsKrI+i0F/W/W9L01x6JqhLnzMZer3XeKofaBlhSPh4/rdCuLtzpBy+pQ30J6F
in8eRSopWcsQ26WTN8jDANrucAmH9L+cX9ZexdNPY86SqrHSb3llWKkcOEh0E4pmh+nfZS7JZGFc
A+b2rzuhlzdxExQy99T7nP1A6Glsv1xJGjaG8hna1/P4JVBVLvUhVB3n4i9ox7Fk/7xPN/uMyiNK
T5uFVUAFP7DZ2j/EE59Y9z/aL9CqoI/BT9xLNzUt2iQ63PcKuw9+4mjL5qR80dcdAFBYZBH+UT2+
ksLhHD7z+i8ceA1ENnN0zh640c4/P/IiLYO4RoV68JcLc8z1ehhA7F4ZA+WovRxEuXeJQytvOVE0
zzTj08Qhzn6ScywobGT3SLsY9AC2q5a7zpM2x7IjMVFD6IGYDMiZftVnxVRU8BrFyhVCdLJDCFoH
xKsSALTPPa6yjF8SRDhKz3yizkORMfcp2WF+GdGYNqsUGWHvj1IH13r2lZIXTWCASAzHUHJbo1ZS
eFG1RzErWSXyao5tiSxQ0P7aE57kwsv1YMJafbarjOrcGkyZQlP7wEeNrpKTiOs7tE72e50snoxl
4GzRlpIFlfkOybvC6JzQqDENe/sTa4OjOtEg7C6hPyIAmzVQ/bRnmLZkA89XIfALAnoCH9Vn6tap
xCB+iVjK1v8dkh2JOw94GtGagEDL6fsyWV5I4Izee2jvnkyplEpotY5LSMjIAw5IDc69O+Vy+Kaj
mlr6/LHbpd9GFzxwYwFehHBRMPgit9rnhJHt+U+6kGKBoWhYzOxO4htLdMMY1t6LK7OgtOrdkDvb
zWXhwF9hLTE421rpT10qm4xBMnA/gBvhtwJ5pWIC2Yqg5GAGAP44Q4bnnNaKJ8nXMYD0Hl0X2PuB
m3Ewn3pbXiU1Vfo4adCgRsFlG9hDSQrFmBjURyMwVQ41oHA/AREY577TKYEngZJ/yI4y/8T8jg79
/pNKcsGNUQ5I+SWM2kBhh3qKp8NDVMgGHnaTAmcQWHi+wunOsGwqFxuz2CfrQPRZZFrekx8QwC61
V+dVTYXiAC+v0b+rhwG6zXKKYFe60wnlqwaYW7VWgVTOjp8ThS4bAVZitMrft6e4qSZUORbDdtHa
LBrsHw/ue25RXmyORtOiuNgd6FFBseNJBx5f4jOZa9NUj+UCyULUjehQoTFTJQKys2CJv6KswYii
ComDwWM+J8HKd5zGt4mdjv/oJmWOL+0Lp22l2Dshwh1/yMXqcPd3aasec0M4TVGDkUppVJt6B42V
ZZvCIUixRIQWBt5Uf3Woht1TvylKUTveutZYJgOeG9UogQxIflYrdXEhpTPZ7nbpCIAwDcN8HlTd
4HY+bsmh3/jmg57NNSBT+l2sUMAW2KYnULn6kiuT/JFxl3VNjObHeJTk9XoR7CdTmDaX0viKQy2O
6IQGLVjaGUQxri6qaNu5SPmbKGf3n7xbZy7LnRYD6eX5S9HkRNNnKLAywc1+ImCA1mHmbblY/UqB
PgrNYV9ZVeRSxyOybsAk0Vvdx/YYPKJ+BIdR3hRp4/hWHRYMEog6rLB66N3JFuntCYvduauVgF/F
udlVU2DYD3g8HbKEFN02mUOowmap3nJbayucrQVmwXhWNFCuYnHNuH9JHE3hARxYS1IO5L+TNzeJ
PEknSj+apUBeBx7aFAcen8gfhuCHreKlcmDdpk1e8mTfYBr4tQDK33CUy/jCTg07/LxAsja02x5R
ZKtEgahpdiUZNT3AsXKjkPpM3C/UXrrEIc9kecln4im0cS+E3rB0990bL1ai+FxlnBGD4bcWXzf8
vs+ZETRAp0w5aMN6KLD0Ez9GV2OaZjOWRXjmhvQN4m7o2zP4gV/jIIz/XluLfobIlqcbG5TtV7st
TF9EvMuOOGzHFm9/L7RXPA/7oUBYksxoyBXsRUFhm2pVwnncV/HG0nuqEC0YD7XDaGopI7DI8TQB
jd0iuUsSRS7swIY4VKCRsi75/t9XydOodU6OrVaOxXYRk5cXaOaYUw2DhkJBuIiQKH3FvNY3w/Qt
2j/VTJLvA+5QMx+bbZP2NQcGjRaVwmyMb5KqAouEkSCW33GvmWEczGnvSLrkMNsZr7zfuN94EBiQ
1DV6Mlr/J7dixG8LQ3PT5wIdVa84wj+aduwzpwBXRcInJODc06XMPm1KrK79zmgOINKQRW07ZSG8
gIKUJRcyTfmuqUVfw8NVpwei1yhSfmZVWJfs2A+5vckKoo5ZlixVTxtqSjMLMvLATWFiPsvUXjtr
Nus+Dc+rdTjbqbg+hI0RVpY0giUtCz/rk5SEhS+FQEbsnLgZddf1hYJyTpJrnZ6bbitBdUfdosW8
flezgLFJsIqIFKmgaSnEROFyY1rLTBHJYxLMfDyGj0vMUJ4/O0KrUJzfh2Uc4pOaa+igAGULowHu
WRGf2lWwQJlncXTts5XdVvgFQuxDwwH+JrPyI+Hul9xYyN/DpPw3fe4K8dGR25aJlKLEEE33GBCs
QLjO73OS7glXbuB5JBlY13KAyR7pYLaA/FD0B0Ct3E59Zu278FjqU3r9A1iA+VNfrHA7xXENJyed
wjzEvhx7zyAL+Ao4IN2S7ERPrHpwU7zQbwPm8z+nNakVpEFefqbEgx5h4nkV2eZUCsEXwLqfUUUJ
+2gJ6c/Q5yqDIRjzlPS5yNnNK+zB9zJ9W9FErlAYZkel/oD1fjtxdXyNd5qJMuEptBv+QmGEG1Fs
5ZnnFoKvUqtVDc/h7nn36ASB4VOxVvr9a4QkaI+8c/O1tcC6rHNpR6fuRn0NTNkry+I2r2Wd0rIc
Ew9FYHbfwcOy4ELb+WXE3xcxkhzb1jNgpTJc8f/SrPfAk7RbCLfRPg2buXgbHiE9/uUbjnZiazxM
tlvkGlF4dwmZ4JEhry7DG0NPUR5ai2lmi0aRIpaQMzxK+7oNOocC6Kh2N9kfm7Q/4wLQRakXQrTH
PF9AWHr6t0pPphRXaO2n9qoxtUQZZMzawhFxJv5KPWRR/62v5tBhtSFDicfA7aFtQl9oiWkW1Y6f
6LObFuy9VzuWO8wvoKxRZ/MJ49UUokdKaGgOaZZPj1G+pQSQrSayA4BHcNp0QkrslfgFiviBkX5M
qa444MlX9qgSrR/QAbselGyTO+ZEbcZTMAMnWb3lmMOqUqw/kJyNIxTfx4ZT7NpnD+mtAlwsj1hc
vIzUaZgujO9M6Ohv2+tJ0Th8K2bCS1UCQcUxxrjs0NntgiRjhlzcnzDINHfwgQWT5MroqwdnsPaZ
dkErX7Z3KzdpCCXY7yowMHzHZLr2rHm0vkkEEBBuUqqFh8rizyyaP6zEoKx54uwngt/Y6aH88JsH
qnck2KHA4Vcsmvk/CBK8SiJ55vrngsTVWWDhHYXF/wCVsfzUthyO808OUbHVydeApCxP+aGLw1J6
oZ3cGqUX93/5j1y+2IOzohQiIU9qL3+Z1/hUva2i8ECkKIONmYf53viHfSOOVBbAOgR0JGZkkClK
OfvMPtfiAqVKuszaS5mRK1K4n0crnkyXZkkO+C0Sd+/oKjPfTx7ajK2b9Hx2La08KcdJp+Rnhi5v
4RsmiXqkplu9t+w/J2YKohXskeIpjGPGOanEvVrH/WjDtMdGAODeSCyD9SxBbNkZNv2K9Ao0GYYI
VXRQ3Hdhdz/sG8XG44aQYuLzGA8mxesCeQ1D4vRT1Ohybx5Z4FBcYBofFnHWtzgHaLwks7oIWGR5
xyW61sHyY7qMlO0zpHdhk4S5Yra4U1EcaQPY3oX8cVpSty7aymRGZEmNRfq+QRo3mesI8Q8Aek6E
OYNwh948j0fgwNxOTIzRkYS1Vpx78PSJqxkO6lCMuXB73ZzXiiAhBVXr9Gnv1WqS4bOEQNSRQgg4
QpQpI21IQXSBtkNmk6NhRTyIZZDRM8DqpJ1e1JCLIbWO20xwcfBfT8JSkO0LpLyIMfyMpukj4LsX
yX5EpGMRsNBu7mJ9oG/T+3j0cvoxA753QBjenTiXV4lXpwm37Di0/3/rHpdX2vXL9InrQgavs/YO
CqZdS9EBNfaeuDjU1JzjsF0GYoOMLY5+a1W6KNRA8cMXg+l07dUShm+e9ywQZkN9J72cZY3H0RcH
Xt8PtDUNI00aGtHbvgczSADL/DATJlb4FwRr2V+2p62/JotYcd9IYCN/ZLAHVxudEFk2O2pndowr
76JigNgWk3EOsczhGGnjhu5GtGxRR0tRfDKIkdApf7fZvQRSvb2V2MyX1X10L8eBgdoUVgrNnMeD
O7pk3T1zbljIGm1Hr5x45sH4HzZBXqanwNzsJcfq4y7ub+nHpQONLkAs/bn6IxMK6KiwJlXSzWaA
7DjCL7a59WhF0y4s71zgiGJSMLmMJUiQIAY5pnPSrin01yUxFnAb0K9SG+IQMepXaW9mgLO7cT0R
xKk1iInMnMdlk9ck8QbzPOeoWYtH+bKS12z7RewYqoOGUHR0CHBmhKMO9SsWIlp6Y9RnkdNC+VCF
r9oDpsUA0ItZjq5V3qpNxt7zeA9wCwUwNDZJw/iSqJXzdUFjasN02+65R3nPlXO0kotDmgq9fv2I
CNzRh6txhq4GbsaRzedTdb1Z4xY3UZ1lGjmWaqHOE9BrbJ0LTeUyIWBDvjoD0RySG3xVmh4YanRN
CZkfSZerJB23HcDCKOcaapidEAj9P0WF5s/BlKJf8ZzATVK+pdPIWnPGcKncK10yxYIbsXaqTr0S
p12BZqLcVzPmYylakgYEv3REOQaeAXYGY1oLgIJFAcNFu7lFLKluDpvvq0AT9HdB2Y1cv2yURELB
YAwM70+MaKTCo4/CpYH2qt9CdW0rnp2S3YigpQB+7ro4PKr9PrfU8BpVPh/hqcJpZugPON0IIPGA
EWj0l6sUlYDY79zpaoE7sLdH7+9A1kXnN2OEamkwhGbNTV4wRLD/1bA+RFmkqE1q15Tz0Nbx4PZ3
OZCoAOmQnzwW7Jurp7kQpFnVDLnGQ8246YxcJ1xAvQK3hYFWXrZExFwrzZXRPfvt2J2HWkvOGtF/
XxK7qGiWE8/josxDLiS3aGTzd014jAIN75VBEDlSdAxs4T8MgZ65xuYe4Cc1tAw4sVGbjXn7t1Pw
x0gJnGbrKBD8aYwlPehFd5rRyPqOsMCe4kzORhWmiO6oP7pB+Ejfo+HxcUtEqkeVibe3sD1ZvNcV
QzObtVR8+3WOaO9CxYrrcs8Uc7WW4kSwEHxXnwekK6B0YrVtHymvwkVt95F0yEkrv2RYmQ4HUlo6
iux/BHMtipZK6j0G5PGHa0iqCnqgZfCtf2tqmmbukM2cErVoWpL0mXO9aOfRWxf242Gyi/e/PzRx
NrKPTkzXaIr472X2u6ZDMOWt7WKxP+0SiUldQbaxvuivhlR/7smCgqXAicdieHJgk9vxLXQ0Mpmg
6RFKgVWXnvjqpwjV87mpVUeJe1TyxvFbVAaA/ycEXU3jgMhfz2KO8qwjrsmQdNtu7kDce8ultRki
tEVErP9k781hB4s6A5OUgZKEn9vuI5bACTpURAj0G9wM9wgVSpGFEIIawzKlRQdd/9VQU+Vxu96U
G06RCJQgewXOSprYjw73Ub00Zz0YX2oMCesmWark4A5yejZSGEsPcH9R+vwpz8YWMXB102jkjTkZ
TjAj6PV2GfEYc6dBVdCLW+u1kJaqrwzInDmdeY82JMza/lQCRALE84gq2yAL2GpPcDmQA5fYuKnA
2ZgOPGR7SKu2wY8MAMYjRE3MRQ1FGom1f2+4b98nYh+ur4cgZ+E+LwWUkFOFDag0BO5DeVFxOf+0
4iovqZfj518hHHuTjVe6SqaWlzN6CVUWBLfT6CbVcXWJ2XbFOwy7CxeHVF4xvD1/vw/uoSnhWcO2
qbLl/l2Kxo1WDcaOHD/Zoz6qVdmD7hcx5W37Xvz4lzB7gosl3n8wuIHrofB1E0haehdkFTW+sejq
fAzSTr0f0FDnU7F/nl1qQm6lK/K1mpFVxy1Emx2SwxjGn0weD3L14L19haYmvn23V9ijfG1zmYuD
LCZGJWEZPNBq5DbLNoPpp49Xi7sISqhXBtuGvcD063DADQ3L2DvL1VUi7LCeYk/d2ssxydWt610w
HGwHYednt8/m8dkCdqrx9IyjBKwnAl0w7lebAhBH4U7uqz5kg6tSyupQvInPHczbDH3bfZb9jxnA
dmWkPG5l8K/nftO49j5p2PMSOfkvFmrNe19rryNc/iUDC7wSqtvkVchnc5LoHq/vS7jTjrnJXCL+
0jG6mwCC/h4dkR1FqxpqHSxFkj1v4pKJXO1b4/gGJsk6VbCLJirUKp8QDQdBQnVLir7/Ty/+qc+O
FX0zkWAExf0hDxCkYzoBbEv68Y7GCImQDbs63MhciD42oxuZL6dDzMrvH1EgGg9rd99h6DFXy99F
6OtD/x1H7K4utoBcwlGMu74UBmrK2Vui8tQPmp0saQQO1MiRRvfxHpYpgPljxPIiw9uLJEzPh4JK
MN49CfNQrcDWJVcjdUhryHYSqf06AIchBso5bcr2GS730cFv3wYtC0AordDQJZFuDhkoOaTP6a7y
XRsG+3sVgqOLEPuY1huAsg4JOIHcai+AyxX2GfA9q7E35FVFU9hd8tmh0ZF2vlXk0xdk52eiuH65
pRqQGuZz7LXtzUZSBwXodkB0n+tMCkMum39nrnaDwDTRVV6gU1tdWuwjeV+2U8RIjD9GRe9P5QCL
8ZmXSI+cQ41bqw8116hSgAmhxCYimA0qrYt4nsAD1ykoqbeWicen+ZNi0Ki1QVOnKiA8nzB8gqAb
+hblm4vvfAsPpLlC+yJEA3yhfnHPiCPVMzuA0B7M8pAHLgwNQ4gPrIQ/yJDV0kkC65PEJomTpSwv
w9PfTAVR5P3lAkAVa9ZIxeJmniuAx2Ubd2SVz+3TQMc30y3YxMGh3NenXKR1/qmcyOZgDRPD//WG
OjwIaw0aLNIkdH4hNslV2D+WffMxixpciR1T7Pwa01hBS0tT2qUur2s7p13ErI2FlNs9XKVMlVV6
4PkXWUWQiHmfwUp16rNr6L8Y95di7hd4TyNIFJDfoie+/jeXJlXsYmeQvIrtHTfg10/rq2ZzWc2/
8Ks/P3E36xJmi+5SXbDtDhskB2wFhyV569FRL545J/OQGt4wF2ZS5BvjFY76yqLRnsS552MNusf4
egkdD3MtB9O5hOMZPaMAp1tIyEkI/SgVG4UEKTNevdLYryEKDkaNDVjfBoMS3+KCTk1Na8vRH81i
/rM4YpJf0GVBc6Wq+Xwst+AIyX+IPAZXAx2V2Rmog6Fe+KQqrAXcQHuP6Ut7Y2miZJmdADlZXyCK
/XH52nBiCsKWaWDDTAAiukHrgPWUTnCUMe9mYdDgy8wAFKrXgDdnCFrNo1vrFAF+P941J/ndjK/p
Dhi9ZRpkqC2Whzf9bigmyyEtpsTw/xENNI+34sUYvUGyBJjaGu8kg8Za9CBjEic/KFHl0VW473u0
ADlnCLJ9MdXyNCqWF2Pab4c1pDFFltob0Z3up1IIW8ODcBbtdlfF9+ozhIg3x3Uhy2S3xqXHyH9z
T0yFl/MBM2K1W/btDw9o25w2WsuOAk28rlXl2uvXiSFOB2JCiTnxFlFZIh1/nXeIu/bLmcoymLVE
ztWdN4MhOYJV09E2YhDvtRTBrRPY1f7LfHyS0U1TpY7Z7YrNVfl8NRkUJERxx92zLpTLRn8n/dUb
Ln2Gg0t6QNNqpdDC9akUyPaLzAZIuI2umunzsDrL2X9iZwsc5JWnWQe5PZx5RVrZVv5EJc9FfOkH
CgjiK//Oen3Dzgi3wH2QDm2iEwbrICuyGYBPC8YxXy3x6tukUhWhvkMOgHpmM6n6CM6A0pg2CahF
RBNNu+dXf3Ih29hjj7NHwdMVb+h6Jn1dX24ANIsOOVe8vFBhftoowv52eckhURMpEv6U/38aLx1s
vbEkTVSGVradq10QNcrtE7ZRUibDvrBIjl4qynZFAd/jfbAA8qBItPhYzumS0IAOM7q8JaEJH8KE
OdoBz7XQZL3DyUKEdVVPE/uywIEloIpBMFFJMG/50XJlb8iKHeNU5/pPLvD66IxAW+nUouyXjkNW
UIegijKQ50Tx7Ee3oX9mn6Bf9P7BniZRRcm0lMIeVpUSUxuHgXof4mz2tFXWYh0ZXYp9W1pP9IcW
qHSFjX8VAF37OsoYH9EF4QFhoNwayxbBXC5D2SJNsFAthd6TqUQjDMbnnXoyG6zQkpT98O3PEl7n
VqoA/VCu33i0sLWrW2JjHPNy6ORBlfHMvtKEGwNW+7/E55bNZBGDC0yqqyY9WLS9/bxj32ztA7jr
tE/xIn13qs98APmmRer6jyGwb/j15MthFA5IZEBxuKTPHrCY2yQpBqx1Ouw1d31GInxmAia7uWed
P7KlShFbXenWfuFEzCYGX6njSJbPyf06wdFvruhIjxlZhECRe7OOoCxEiROIdPbszb+FPmKbSrdX
6T9whpPKgVQdbTRCWatYtFcrC0FUKpW0z8wzcNKD3ifdM8QIgCtyFvWqCtkURjuWuYcgtfsxAMvU
rrifPAHmYgMwLkIZStk45JRBEl4JmTZyZGa8u5BqBGCz9jwomrHRKM3f0MxMPHT5egktoJr41uBO
8p3wKdno6kRs4+pLIJ+uXUmaKDmVj6wAQ1VCQFyaiE9VN2PG3Dxsqkv5vICj2NXQ7sAKhCss6utf
DQeBMf055wiOVk1tN+0Q3OurawVd55GDdJwZt4itAXgMTWV7nZG+o1Fl2BrsrKIsxtoc9zouBTr7
ofvqlmmlt/yqR2RXGvYM6P1c2MeC8ZE9+BVdVBnKD/tOWejXt3KAw4ItInW98g8OSVe1dz0HB2Ax
FJbZRjh2DkdBpQmYz9bBzB8TvJsrFgzise4vNSbcIvorYfA2JNJjpIwYaUgIRREFhIqU6z4UKzCe
Lfj9HrRC3KKR/tQ8UjzkM0a7/N20ISvhhkOXYogcw9jBSOPK3OQoGwhwM2cer/gtEJmaHgRGQJWU
6MHc/FsgmkWaIWnKymrMs4njdUtFhf2SAohLRZsaxljSrbtvng6MRReCgbsWkHMsPMiMWFI0KUgl
NWVxBtlmzxsiEIDgKXHA8hpXyMLWiuh6WodolHRZ3TWvtJEJguAhDLBFXsE5LIdwByDxU3HLSXIB
CfklsZd9egJRE+f8dx97wcxq70uUWu2mpk33I9k9cJXEmHeaLy1YBLwNetlJCuy783QYPHy9b75G
7XpLwfyONWNbfv/Kzn1mLbBPilzmUpRwM9hpfO1n90cPpyL8IQ2hsXfJ06KsmHhINJCY3K55A+gd
k5oEmjmh3uoiXvCLtMIrQWT5/i4pZiVT2iEWgJThZ4tc+xMrHbeQygaokjJBn+dZnYasdgCtNqnO
1N3VXijIV3p0Amtm5nfaHW+fIcMqp+kYjzDAJXLd/+Si1+nwP5HI9kgJ1W2Z2ntngU6A3eMF39tq
v9UjXuTHjooC1JgnRHVef5a0evAkqtuAmW/Zfd1aTHiSMW5LIfUmc32g2nN5se0BGHYlAMb2Skf2
G9+DVh81Lcb2GYT0f6wCYeDK6rIGwhYO7P2toSTAwvpioZQ6lC0vXWbVTAnOugVSOcyVUoK/ZXNR
bIzTTUf1UeYqdGxeKW4SXH6++wLc/3Yh7UPU46dv/rmw9uiiT9npxbEmzK62t6MiFWgJhu80wh4Q
Wmonn0KW03dh96a2A+2j+/CKTM8lyhFyOonWpUH4XNSCsHziRP5fyaV6Kn2xgFyb7goafd2PC2fZ
7KpEXPi81wUk9VhssB5DPuCHdI8LtID2zBKcBaGaiy5U0lsgyCaJSAsMAbj1UNj5i304mUd5c0Ub
TxpnNekBbUDbmY4vcHUZ8srnwisFFcvXG87eKS374X6UggVXOdDkKHCurN/L9Vj73GoSOL9KP7pI
3BV/MB3cDrcVXfs22e6BvJURVySnu6G5ETXYvaLqYie5qcvJ85sI6W6hUwlRmC0vHrv4wrrgFIit
ZK9x8zBJzpR7fqIOJfw1Lu32T83xGo3Zo+ZBQHzmH5a6w5NrnoUDju7C2whoYi/tYZGRa9hkieLv
zmeX2dXvswv2HXfBu1Ou8+KzD0jWaniV8wv8qInR0GF73tVDrGmRvJ0AwUp8nFgR94Dr2AUEHdgk
gySVl+X/SsawJd7++7/btH+OSh2Z8iXoKZ1wBPZhTNRugtVqhyP8+uWaJzUVGo++AlXaCLVlvQcJ
OmYMDMC7jVVmbwUqyyFUgQHRUsMB0mq14AwfXB/p1RKcVajz2KaBx6/1NLY2/WNwnS2Pfb3AXYEd
Z61Qu7Tl2EsN/cRtpNGZP6+QMhQXJuitwgck7adLcndycCX+fTqyRj7j+Lijug2kOVtcnnjY1eVy
CpsB1nHFNq3DEGFg8xKcXql9NX3HHqFr3e4Lx3XKZiUstWq1n0a07nwhcNvehAYCQ/VbO+2liF9S
N7J/Jkhr+4otXrU2gPDjOp4jabH47KL2WNERY+mzTPXTp2CLWxuAkIuX188ciMxXEuKPVIwSH549
gGIy7zRLwqbFjWyxFO8k0hRUuj4XvpsDDhl5Y722dCb7XSZLi3S+3zWZ2T1LIB4L1QdYT1/0YQTP
rs5pEqsZXVO2jjwGWSHVzjivw03L5M36oE5y3TOLtLotU8vMMaAqDis7SQx3EnDCcqiwrvBTSHpL
8zM+9bja+wm5exDf8jtyqzIkjw3nDiwyvHeKToxNEvCex3EMGdEHoAfeezmLMMkRQpuu9CxqCwMx
6l4fLn2LiDNz6n06SmpXkbthPYAE5tjS3otQCEk6/9gvK3XUaRqRQOX07esGDI9HIsMBYNE7zBC/
SCCR2tnBHRuBAX4ekAA2DFSpr5VeO+bT1GXLZItkP79rdFHiSK7AUH88qvoRFXvr63Aje0aiHoem
VSQ+dpkIFaKt9/NR79pnbS1xjbLQVJpYEBUmkWuqykCfnSbctkT8bd1TvftizdUeS/vIczNOjrF1
bhHWC4iBYBcp6VR2AZPtFQVXY8CN6+tjkWOUHO2ooZl1TlK2sEHp5Tro4yaW9fOAUMJqNST8GjpR
Job41H0d0vOgitN1xcdzT3RxXCv/o1xdyCW7uiW0ZOyDvgnmD7XyeDuA1ztf2lau4lG3NcJrSEfI
1aI4maRzE3aOd5LCFg/NxlPtgziwjU0a+xFN59eG5hRt01DXUP2g+4ncbYRcgbjOD3oNvs817F+g
bcEoEJHHjQb5ypHulN1ZL4/04RMY1Jlt5sDnkBOzmwSCa2UkJD1Levb60Mn8KUNujeUj+wX/n5e5
cG2gHktUZGWEzG4EJJPq/UZJtIzDh0lJLtOU+0fMZh3TsdCBSIUPte3AILWjBR3CRGlRgs4PZhlc
KS7tIaPiLB/MMLRWVrs/oH/30bxCUXufFL9CmfXia6kx19wRkgwKg7/4nErXKmv0uVZwnDHMm35H
DFEJFTFGRuTOGgsjL6mjnpIIBn13wDKLwkD05QVRQJDrzDVtGd5QinRrygd0JqcxeoOjTosV7gr6
gJSMTJIDVyKz4Ph8qha8dE/RIJEFIsHYEPg1USQBoLzur+u+I873r20i4huiSh4msDhO7KEocEga
ES3oL2+1tklzfSf9AZd7YJ1A9LRT+Bdw661/kJIO4ZDupvayqVzYG8xe8/l8NxFerte4//cqd4UC
q1LTTvFR+ea3XGSG8+SQxO4woOTVA3Ypf1O8uQjhw3RnlTykm46tCISZDmDsI8hiBzkiISoxV2gJ
+LjU4GWn5hupFsqJSJ2kPmrTwq9CkHYFXrzMat6m7l5B9IzB7kZYX78H4O9++8LWlScUDoF9lWI2
jtaJ5L3svc9QbQ7m4tTVBefIU61LSxwq8AfFJeyeQ5atgoDd7z631Whk0ASObE/VM8vd0TdRs4v8
bXY+rwLQ0NgD/ys1ghJnE4gVLdJAo56844hhzBTni898qHt70r3S7TsND8iCrvOUks4e7dOfmvwt
Hvhm3xNwVBsqNKfgvbY2iNwEKRsFVj/bCQ/RGtgKfd53atgaWXuYoI5xASLKdravGpCBq/ylnusV
5ODROmhTxqULGyWMjBlPnA6KzWdIykoP9Iy4KNnoAgUmHWYSObR0ktnd3sXrnCR1Z0yznBvan8ir
i3asjp6hqlxyz17acLWEn7dqHcmoME4cD9wO2VFxb+q84CUxBei+2BIDpiqsyeb3NiKM25UiCjua
V7fKTgEJh/F2OGJdsNxs1f4juIwl4MtHUxsSnDLaz8XP9IboZ3mwSyuI1icY5Ac3XJevZVSQlBQY
S4WN+EKHv/1XYLz4kxQAVk/9PZy4jW/vi3PTwlLJq9sXXN7iCiw5QYY3OnpNQH/+yleZh97q1bS9
6yl1At3fdKby0aD3JaKF43bpoNc7RyyxVS7yYM9AxqbX8z/OEWgXtRicvkYZh23BUhrOEsjjahJu
EZktXvE8FRoTXlTrSj9VsjnkLThgkimZvIfQqbh8v33Fs9YneuFNBGeccvCemnvlizJbGB9bYc+P
R7OpE7EmA1FdgsCIR2PcY+pVeP5d7/KeRv2fo7ZBxy+Kgj7dTMBxVj4j+ffdNucymFSwmIDyjzqY
ME3CFQXvHtfIhaxPYKjRtWoQucW/GMq/EqoVMPuCBzL2hzTkEzZRh8XHcL0VkaL4zjmZeeO8m9iP
IlsbMlv3JVJseAy+F4hrvMPy7nc3rF1cnigLzrh5PWrlSM1kIFhTIIelRWK0U/I48xbTQ61JhmWi
e/KwWEhl7Cu64FZLaJp5LJ8OFNFQDiu+O4hsYY26ztnyglqDSr70NYGnFrAH0zvSK8pEAN2i0fDZ
qHjhUqz/05h91ZkZyQlFoFG2EzJyb6PWbr+o7EaZnv7qWp22OxAFbzobPgllJZ4TVGs/frR7OZDG
Mjel9Cu2VGR3kq6CsprawYsYbDn5pr3O3sW4aERunkC/Av5ujLrbMcxFM2fR1ClymOuS9tXUt3vC
PJLUtodpF/VSnNXQpP06xdmNs0x35f0RjbDGv293asDbE5KbIfRA7UD5ugHxCtFm09NxS9uxgb3w
EZLmuD5K18YCnmAIqFLVb+2rK/vdyHTmGb5DAiRymAHzoe20HidEvQ+hYn8SvjSoyg7u0FgFkUnK
Ev4Q/BWolDKR8o5zRj5Qs4k7VY1wb4SHTh4Vbbdti4QPdKtBNHMEwhMow64TL/7CB/eBjUpg0MPb
Cr7ZlJql6vLtelcejHAygRP61u5YJ14QXXjB1vo/fRRt/balRc0sMoQ7tmmxB4QEzPsIBn+wc3E0
DWxhrMlosQ1aTp8QudnkROCCxSadyHuqbqUvAsGTqokdKtUmVaEfRx/rBS+/CXx5lTuLDDHlmJ1g
2loiMnkxuNKmv3uJo7e0lBwJCggli+S4R8Z0GN/45pquE0RB2cdstwr6hQBBF51cRALCoZ8kMyso
OtHup0N6dmf8JrE/SE7aZRud6tGZhLyL9mk5Ttgs4nCyiYej1O7eB+eLWmu3muszTtIBtvrf165q
aG3Lg8zxvEO87M90/JKSo5n9bPocWijO8PlDr+lRbNLRNvsyg9od31eBINxrk9ez1mWw4Ib/re79
NU7qQ20C4U/ygAATVIBnl/eFDw3Ld+sjahjb9NEBAQM3+fx90KaLcBcjMe4VQicgkUH9rgfC/buc
QT6XmG7IpCvel/3A1nT1I1w8RHX4otTO2RN3j0Ecjn8lsnCLfsGwpc4VSbK7Ts83OK+ped9LP7CY
kSo/hjzBo5mwN6dKwnnE6P4G6rVVZwAE+gKRaPTvAVLN+aFpWCd7gzFvVrw+bD5hegeobLrOrFlP
ZmgWMT8i5bINMO7653ROD/j673tTRSU3bN5bvZF5oWBwdDX29KvKxOwL9I0VjTM3WtfjuSC7nsUf
Ush8KSnYtvDD2zTHj9qw4ycYsWlz5GUkAp2VhCK/UqHQdF+F47FW8AO2SUQCcZ9JcVouEufGT+XK
JLp6I4TiVzkHmd6A4ZiarWQEN9VY2EF1c+UYhHqzxucd6H8Xl3LEn31LrhcxP4EH0W5EDr+yDth9
jkrVVcfcivVyrTLouXbq2MuFIal3yCbfEfSxxKBzUha/LaEb19S4Z1p8BMDX7hL7qswRHyCnsKnc
bMpWvSwQBItYSPdSAMn6mzahXhS6+i4qLe4WubWQFsXnVfN4yGMu7nuOP2vKicNgBRWaos2I3mb/
XkwaDqytNJNvcYvMGn099qAhOZ8RBigrwKBouaLC6m0Xa4EwS1IK+GJHReo9hnniryZObmGb7Gtl
ZfKkN7yINVocnaPS3a7vrJTthCVDF+qhkggBfeTOGEZOcOSEcJd18OqK1U1HhqcW/BGLM0IU4iYS
EuP192srVldF1c2pcA+fPpCjcMHMuhQ37JaGgpUBGYcrdIJtE03gZAgrQGHsPXMysZ17VlFuvfJb
HrhBMliE0qijrNDDKsGdWbrgYYVs2vjoHIcgOkezzS0Ng2laK51ckIGyf+KfJqxoK2iFRazu/AYk
m1eaZ73oDbysVSfvHvVa1Gk6J0AxmCUk7qy0mgyOI5izztjQNZFr5Z1/LQBJMZvBC/4m7CuKWLLb
HAeZq9Qw0GXt95uogwK/9yaaDc1qsprvwVwKDdKkchmqCW5fyb8Z1shuJEGiPhjrPjs8dSKHxFK3
6BpHgkz7MNb9MW4uxj6ln2jb637kQbr+qRSrdXFDWWZTElnuK6YpZUV8VyoOVZIX+RcbLpo09cvL
me5LEybwsIEYisoZaZGp2jscUUpJ5zIgO26i86dwLr2PUNUW3poeHL/QQxDj3j89hUiEQNZ4ZnRW
4fEB7RLafGUbjifJCrBibvTtIJfKncymyW03MHWeHGtwMIrIDH/UJ2KN/gO1LP6Hmg8nU+zWk/1o
1KMib5CaxHfy19dCV+GtuMzbbA1KExjETbXlXaB84TeoPjaTBxcvbbhWPcI/TGT37rUX9+HPZLXO
H4R89O42uv84VVAAgWeEBanN7KKs1CImf6lj936Rr3uHReZbiiGNKXHLFT70ixuoCRJlBpUt4q7y
gBFp7uY+lnAO3cc+rdqTOWA7Hd0rABC3g0HsIv2/Bdxkwuc0I6Uv1uV0fue8LxTwDtB/HGZFoEpI
oOrzqpicSPuRCVgwN9CD3ryqbzF/GbCjoODCJIfJ+h7c7KosiPAp1e1bnEOryuvRcuy5vIE0KGCd
Ntfu1IyBrIFTHDXT3uWuGcXt93mklIB1HNj3/2O6g+hwbjUMWpGVWpAK5LG8Dc7d9n9A3jKBL+cK
aWPzNwqrit6ZdmLlanWs2dZUO/eDVlixITWZKzYTajYtbWO3gUtlEEoBfuTwpmBzAhv18m5lsnUs
PnyhvE+tBs4ndP5g3jLwL4l9jdgk9a9fiLJhRl+xe/dOR+zlvZGf8YwkuAG/x3sL3BteIXjZ6vjl
TgvfhL2LVyfJ4nkwE/+M9r3I6MNJ51/s//FAW1/pA/CQW/sZjddJBVKcPeh4TBk46rNozfoHuO3F
qiiYiRNknD3x3XfNh3cTItz2oZis+2jmP03evGZvHpJY0yz+LJ4GJevINNcfWDK5yUOKGcDTh0Dj
yuSJqS+WW6Rn/0M6s7B6CgXQc7k9CbKZqpNJAYkHLeM5ZUUK760Eu3xBknODMH8AxFraviU+/TW+
cTPYAC9MgLoskJ09X7lEoKE6YpN+saNJjDdW9tIjVYlVmUr06m5LL1WD5ifJ3Y15X7hxbN3+uakl
4HD5e76T83nRaykrg5VRoa/ASfNJcx+R0flHVmsOsIYjMInU8Ph3lyUxdZXPofoJfZH5Tpzrvpti
HBxxEqEyHJ32e56zll3MS4yyrgX1NMto65KWPRLR7X4+ENYX7f+A+T1rB+M9D5AHDiGbDK0B/Iwr
I/1+N48j2yUzGL8Ad7hZfmf1wEBz1cgzAuX5q/LNLM762VSdY354VPLtBRPLjizOiczmLVneSikH
LhE44SSmdBTMWF+KwEsf/WvSaJ6jrwYgtL/cGk/a+QLX9/vz0rdlZmrGiMUBzIY6H3yY1C1z8qrI
xe0Uso9OlgUAAndYBrD8p+ypUYbxUDyDcGOAr4WyC0+twdB4AW6PI7+vFhZewPhPUnNJmOWlatjL
PVoyIz7kEvKqa1LV7zwgo0nHZnFTeEU5qeyR8c1wJzqBFxuKQ9JwfDx1biofX03SE9/sWD8JZlTU
PXj4eRKNh4i3RF0Ue/8rwGsz6/P/ZWG2VaEtPtpuJH8dVVYREI/dlB4Ci/ZY6P5uLADZw3EtySIj
4zB0kuSNtGSZzr3cHOvrzrBVRcQ/9VQxHdhluoNuQ+kwRzmpsCckahKFFFudnCN/xp9P34RNZXsM
JiCmJuEv5zxiR4N+/b8vMjY2XTht5TL4a19WP6oyJ1ykoYzHZDuTRLWttVNiTTX4kb0wb73bKOZ2
8HNoln6YPXbgHSq+pdLNfOOdU+ynAR1079fm/TeKbr+YOLKpFAG/g0B2G5HhPhyuQXbxi/fePgo7
LnxFxAuwUqpPYp+J0X92yA2yXg7vEHv8HuepcJBg64/7wr0ahGX+7YhLbvyApIDPSrwjMhKelcOz
tFdkMbCNTHiOMp2ThVcDkWdtHiORXTtSEwa7FQ8pdVLz3cYX4yBkV+IdAZpskiJSF9jiP8mjV/bG
LSa/AK2X9YiGofXFsAQmOT5HYIP80NMY/NANJgGx54BuaoIHV957Z/sb6LK0sKUDRqvEgoyTeJp0
PLmyZhCaR7rhvfv9r2hat9vPtcSZ8IAI0hFxMGjJvnDeuyIFY2F7fxAt3VpQ3wmdmlHonkB1QLMC
2IcRVQtlJtY/rYo4EmerWrB0fhv/95HIoSEQuKvS9q2QWXxy2D3Kq1i0OIlOqo8qC6cCFL523Vla
K8daCAon9DIt9O8y3Kle/JuqWs1EI9ZpRiDY33/c2V+DyKoLoqUU0/Qf7LWNoXLrN++NU46MAP18
MChAx3gfidCWWJPIfYhDYMA9QsCi79wlQ22tP1NoIEqXd/t6PVeUWs+ts+WtKfl6diRA0rEjDvYC
DLolNnyyBaYNW0Bw+U9gW573OxFxt9XE2FWt1W9rYAdkmk/HePa/3362kTlXufhPVTOFA1lDcNl1
grCLIiqzup2U+TE0krVxlf8NB0qt+sHJYer2a1wu66bjW5jNSwCENaFKgjPT2Fl+Tkq388OSD36u
55ye/rbU/Az3DQ53WlG1lxbG9MqnCiUXhXZonarnkXjoodvt1Uj9lwWRJqO5ZqqYZfRfs6o2wDb/
pX942Gr+B1Y/OkslirX4bjra5YcPygd2eSVBfxTphXdWkXqR7V4acnLO+crmpmQpYK4zcEFVz81v
JF4c87PGStALZv3TxwntISySip7vsJLoy6P92eSO+gR0oZSCE8tnPKAMlnD/jNiMvxzaex2quCIB
cpkYReo51KLfirQOJDDozx49t9RkgtOT7h7dDRFh9dKhoXKeLJmQhymfAZEKBp/Z5zdbfuy0ZDd7
o7RVt6hgztVANp8s3pBpxGL2Eyr9y/AteDKRzoTSwIoV6bdeDIt7L+daK6iO7V+cRIGFHXZtw4zE
7lz5DTTzKEHPZsd0DQwQwEBJ52p7NTu8S8/HnkKjkmouip+kKP9UWjKr7FVEKpe3oYhb4xdiqURw
6mzNVL9+lRiXkS27Bm4KtpQYfnZXdg5HHLsfKYLHSfWz7NnFTdqX3sDJodTYQW2BJvGBmuxlrsAL
R+6PVQcxYwzM8fuZAdCkQYldmUrjz1Slzns7vk+YaN8GqlrgLYbCSroaY+Uh/tVeIxO89Ggg2v5w
7gbdkV6UIuEkZZv3oTsO7MoI9FgOeSWxsrUEZP93N1+jkvJvqYuQheK5awtcdHI/yycjxp8mJ/Fd
uVZ/mGlC9kbRgijKFATdMakGi6p3DcZ8PJ40vSMFqzieyReDPDBqgRhzRiN/FvSAa/pHoL+EwUbb
RlbTOZOyFWUSD1eCmTTbZ5eK1aHS8kTknVRw9X9OjIZn1p22I5MorcZEWYPVKOgTdkiwyjVOQxNx
DZ+Dtx9s6gO9xiUGnVsBkAZ5CRtwsoNzvyD/R1z/JRd0A0RAh9x3LLJYPSh+B+c5D9ulZV85q0ff
rXp+H0EKTuFZd6I1T6FaYrgwNVtCZ8hcvkMKxEkxt9NvdLhchO1tOv5ey3+RuGUA4ArLmw8FD294
mzaXFy9QxyylNbGARuISPxepTwFWQK7qgmbqlHdkbVYgKtuzFhhV7KwXP9qLcvny6oQ9yhx/zywI
PaAwHYlA3e8ZFk6U8C9/w8t5t3BvnCQZDptKSWa8X/2TjXbffydlxctKWyW+akEOyssjqCkuphzu
aMXuejTki+DKr+eRsv1r4aR5EeLLVkBAHjXnLNTLsEVkpksiv2mQExAXpC6cSNodlAz5aTjKYPYP
8pcR+T7evGoyE5ygaffLQsIkTW17Xry6uL3pLjBNJFYUvWhd/k2x0kzcgWD5bWsbYjrI1mUeOZVV
9vMRDZMeMQZPMEGkmG2zM43Dh6INIhxGAwa1KuahUXq7M9pGPr8lvK+t42OzzwVgBtlQAg7cu25z
rwawIO7v1xjkxJo+UjBlRffN1Xem9eGknlFeSGCCklijtneHAcLsH/dUhHkVbzYMXP6P8DVLgkeS
+YLg4yMKxVzkckgmqjOXl3mrsLMSPl6HfpVbeEA5jHarIEENTRNWOSzYMpXtfWo5OcfEGHAW9/DC
/0MK42W1NnI54n+lO8kz2xTqZCfqTcxULqU/sy5RjV/XUdz6e2FKBpMxk7zwkf2yDn9l3YMpmKyq
NXQl3GrvwApSZ1g2//hyqCjtHk3EUBSwxKxwzSL2A81UYHmdBHPJyf1Y3ft83jvK+gs62a/mGXUm
w4OTmfR3RQf4ECmmOa3cm8lbefPH6ei+ujWD2bXDpuHCofd04yg0EQhEOaUva0Ey/5jEFaioMTGm
9R+V32R69QKuAOSbkrfJCaP6H85hEgBIsdw8OF2cyQp1kq5Dx6k9cZS1//CFQe7TEnqkpXPO+u1h
qfcMLr555usvO/UcerVyxNS7UN6nxtmlPeazFAl1srliBB4cy9EuZ0JmEHaDLrfbIJ4q0sTEG/Xv
FVDTgTtwEgDq3d/1de7aSAm+kxSh+3d+9KbWNLLd5RAIVzpEc6zgn6ximvxyGZ8qcf6YetEcDiAT
mByOvHXm39KjXYVukAVcfgyWmy3CGWAjZtjd1dvI8cxIoxc1YSjMlocLYeKR7CE1Gc892sVqCpWY
G1wE3SxPQS6gq6HjlvEB0hJQt9hN77V4SQwG+5l0M3LLdGGq0A99t96Eulx0y4Jz0kEYPl1Fs93N
8IDIchCxN/Ok+jeiw8Y/gDJJHjcLU1e5DU94zAenFUcUoWTTkNHQSRu0W6U7xJjnNTmOhB7ajcmh
wzbjacx0moaVQ8/VvrMsIIkWl6U4WZX3viNgfhFelWzDo+bT+FHBK3EyxkuNUf8PP8CFE6mpD9og
TTIUnD3l4YpzA1hgyJlFBiuUrc1tO5gvE/olDiDd2ZjNAvNemsiwk0POlaC+NjmTsiCa2dKGc4Wh
CNVcrwJUkyZi3ca4rsdWrH50XYdaexSdOjSGKATU+bEW6+27Yb894fbowWDajOVH+S4IfOSqnK7g
8Fw1ir5lAj3285hKzwZomUJMFr+UF3cf0F0w03d7s2Eufk+NJ8Jo+CzwsJ/iwo+Pjz7ILctSqqJa
1OBIhBTlEfqAyfpEIZPcMm2H6NDWkNyhqA2VECzsAndGVFxcU74uzNy9vJYPOBsBiGbmpxtgQOtV
q6zSYoMQEXtz1jYRM7rM07c8ugUnF5y/xA+8grxLTPWCNb6cHw7WoPOpil5n1yeMBNO8uwPPdPmE
9eNcbvcy5t455R9FiSoqZvl7zkQS6jeCuYsz5KAA5YfytvAJ1mHeedvf1RY62fRL4nU2m0A3GHwg
gdgeNG1qz4yZLfHNfN2tcKClcE0Pl4rJv7IasM/lz65m6r5WkoFytYkSVTb5ugt2Myu0v184wW2d
7FExzZn0c9YZE6SFIGwPAs9i1bIwNL4efpn6an6PfbJGpvylkSu8ML+pAaZYct5tX0+PxvhCUvLi
IwD4FPqpmCoA3XXpJKoMU/d8zrdMSFYNr1hK1cUp8oIyNqHVxnRsp4SdTcFe6Lmo3m88KOAdlqee
H8KAzJKc0FLynbQ394DRHGi2m7440NxcK/a1Rkipp9eYnxDU4qkXjwadlkd6s3Y4razDAipsz0iq
yXkZr5ZqgT0AzZMYBGO9tYX1x/dn49xDJVzEtkSPghrGMrvsoukoy1nx03wM7r3COT2C43XoCH9W
4yOlIMgQonVXssX3QmF/AuUwJK6kMkO62IOWwqG6eKmodF4mtssRbVjltGOYW3XzWp6JEkbZO+sH
yC4FunV2NoBOY6ohn86V66+775oOitYixAB7ZYkUV3v8B4CMVHKc6g5+MJhIbPNDrE7DFiDlYdhz
Sb6qOjQQCd/zaNQLKqiJ5TAJtdhNNUkCOy9PTi1FOJskq11VX3pFw61I71Ls8Ecmb8iIe5l8ccQt
xLpQ0VQMTmK7v18dJ77slg6quNK6zjdlamL59L68q0l3sGLxRxifdr3y0ywLHjWvWnVajjarjnl2
mwSVXlzvEAVD2JaXviOHRIPPjT+uY8xxamsWa56lzb/gUYgyj8TgpC+UryvO42FLF8V850pmuDAs
YMb8T/td9uLwD84sTrvF0F+GWkt3MbM8fxxG4Pcn52+njLJczetsu8se1QlGzlmTwFwtLIEeMruK
EviUhfD5ZcZ7y9Us6ccoM87gkZetBFd7P/oIO5ib2VWjgdCl+wYY+851I4n3D473+P4ijrv+nIrW
5SYzrCMcrvPupeLOq9CaGi0L9ctWHzhBcVk2aruKpoC9R1fAc18qZgaBTLpHAIMCGKoJCPOa9n96
bI3wj1nD5vUIf732oald+38aU+UUFHaXnSNudK+uifXnhaPgdLLxBoGDTf2+tMPssqTwXISiAl10
aEC/g3GCZONNLQIrMh8wsbN7QqSWPU46c/JmDpq05VsgJwhGhKECYOaNNviJHuCuS18HoAmH6aJj
S1ANumxPIEgRxBHe1q9/Pz5U5XHs6nDlDxTYnlcdINiLfHAW/YGFPTcqJz9DgkK9MoDxCvFiEYKr
iesmCG6HbiQOOpOe90CHtQQIHPJPk6KbIuSjPKcqmoPjW3NdYoJnVV2OMTBy9lp91WdSVixWEZ7o
o8y5xdKnOj8WT4ahzbVX/YNuA58QWE2wvnZ3uLHGqPyFZdR090B3kzwCkO5Vtf0Z/2cy7XRid0o5
n4F/+qOPNZqzJBlxN9laQyoaAiNrWtI8awuPAT+y5pibN/RwWd7jDpADfFk5gQMgcvmRMXPcv/mG
ooEgyvtTxmIU+Cf0sEH/fgo2mawINN4RoZT1RenK+tCsGjKVgYOAnKzGNoEiGL7VtJb+OIE2HqxQ
R2TZZ6+4AqoD2rps8lY+33F2jGNRHWbRr+CGNF4iqMeyUX5EUORHEuTTuDJ9n/skDWx+hdzbHYX/
V4RZVxw5xjS2oCH7XX61KVI48V25GOSamJWEWzheVEDFlILhdNVfx7TFgYot5dnDAGZp5jd6zueD
4ziHmQdDl0TDclx9PiCqC72/d4pivcwxGPf87cE7pXzVBQ3ofIZhN2lQw9+tCXUm3z9G1FUxJ+hB
ezQHDtuCeKwDHbJkp8tb7kpRwlsBuEFcxkSoje9kdcibnc3bbeLTGRff6rKi3XS5xtMWi+PQRTwa
1S29Q35SOaJvl/APqrXJIVh1O38o6w7ijyThpV5DRsgIP8ip52Ta1JD8kd/egALKaYy1JH9Gdpvi
Kj5MNjryDf0+LKanZZW9JvKt9mPkN3g86yCydvqs1Jwu6YuUCzU1FUn8CSRyZTndqCGozzzpzOVg
652dgE0YZ19ShyNGs29YQK20xUKOwPLjZoDO8j7TUTvXDdrkn1UlFuiKDYA6bvuoLIEKJGhdUVFj
5cAzeGkdFc+5PcE8vbV50uJHLmOhSthOBm4qokVsX2YsBQ32D+/FE/81ncVSOsxWVFIHnayEREbg
HiM1W+vohj8x7vTQ6qHDM6qn3yTM0I9MYzrG0TL1Ly6/kEtDRthcM1PM6iPXjqthz0mvGk7l+UYt
mQoJM/yQ1x4uycwnY54f3DljlHm2v4hGyFE7dFLKLGkK8BDslAaLkpmuPDzI2qWfCPnws665g8Rc
yl5+dgj22YDaULTY/t3Xwa9N/16NLLuq3fz4Klyj2YM+4saBp0VnlgDE2uquxVdP+ycrUC5hA9Tn
s1E/FZ9DJ5oWGAXelxIwTbTwtRv47nhPOt/NR/8tNBEuberXH6yr3Pf7FyVqEesmQtIckGMANzzX
wHAsRgz67BsDmZpfDT1DQvRY8nARO0LjfxJkRJa1/B/ncb7VL6ZoT8XHeHM1TJBQQoC28j4Bp/lG
8/KwSkLZVc9gFL0vP/xiIRVo/V/LRduA4xvU95ghFawMYxOW3uu43qH6UINJJKMBf8zCj2typdaj
ms0+hNvuVdT2sFSDsQqDLzEBZ6fVJFtHqaQKeNMNQ46WUZewdPXs8Yx+Wws8z/jYFoy6Cwue4hRk
BriSv3yx78bXsyo5vPb5T1oZ34I8EZ1KipRbrm+SQet/2wmLxMeIoWGSuxGz3ZvVfaiWj7bnzLLU
gXcp9MEznoRSvrAoRtZB+aY3j5HCQFVQ0G2RXhQQv7BJc3w6YDCGyfwybiX68CKEOKGsG0erjXjB
3yYkt0eJYdfYBK/IjI8opS18zoPESqNrxtzxHIvxcErzJTEEt4u86igd6ZB2B8rxePr9WA0Y/JNb
H+Dbo+fNVXlP1jCymhKe5WnTCUCKWydnVh8yeLZwQOtyx9nUvwVQ4RPU4Zcera08VStmwoGIirPA
95ebs0YbAEdK6OezKbRzu3gFoZtVLm9svfoFX17KzLtKmKC5NlnS1BK8/P/3B74GLxxD9ThmF0aD
zehi0XW4OPeVuo2Od6QV+62ejchhyhJJhYNBXqLUNVpA6V+kztq08p+EQhQaWUTTd4UlGTJm7Nvk
TlI57XiDZx/LoecdiuLFyBqd5aTZ7gK1WxS/XrlKY4V2JiLE8Tv/Hb8qh3BS+x8E9IZHaE44odcO
DhL6Ql2xzz0ypIOYzDp/TAyxxyFnfZNkgx1mwWmJ6M4GAfSJb9fPPEVlhDA+ZfVZAe4hBhKWrWxb
rn1gZhTNzwBm0FvjCAZnP8HOjNFlqz8p6bKOxHceav9KbtRraIFbyFL0qdS2vsOyGfaispdAqlpb
VE3Wm9Xil1+gYcFalutHGrDgyLYelygsi8JkmhVrdvJolTmALiQuJqn3pT9Y6bw/UCfrwZyx4dva
7D82twaH+sIVXHZOiWzu/KbX6HXiOM2dJIIoev7peF6fSebMrF43PwDmdGLwI+qcYzt/PdzIPEqj
DO6vA6n70lU3WGsCYCQwbRpiTJ27hPsmCFQTTWZgXEeL2Wup9iTxkh0d8qNjUMvTboYdDaJuNuv5
uMRiwgFmLZGPc8t49A2DyLrwtKVvs+W0lGzNlAO6TcEMdRWKGIB/oGBj8WUa9wRs4WZ6tWmf6Uem
aZ9O87F2Hs0/JthLV3mHWRuTC93aHbelvD2OkNKfFlvpWIGHwUTR97JHpO/xNOHUmK+AyJSkzJPy
R4+iseFjSkNWcCtwbwE4lZ+/yaPybpPUQBU9wlb7+J8M2wlcHMlmbnmzWEXPVp/q7t2UpNsJIWJq
sgN8eNlpU2XiYCB25XJ+F527Kt8LuvLUkxpQ/DPKU1Nru3aL/UKUNqRBbJTA5dU2SUFILwAc9rhH
l2yrNKDQNdWilkVCKOZo6M86T+1uIKOPk2do7w3jIU8dTTxkPWl1Doc8tMm6tBKpet4kGTUOWag2
gON6VzJJ9ccefqjxYGc+OCG5LnDMM6W5EgX/9WC8clwf8P+g7K7AVXZpCbKX93sRzYpoErFtrumK
d1FNQjmLY39oVUkiDpnY5FgghjlSSeU9TTGh3M0PqDmv8W3Kvu2Cwc+RAyvw2NFX4Bs0TmTL8NIW
qUuHO7tIG9YrHsxYitR0mPx4yseaurdE7XStqlwOBahfa1xkvzP7XL3yiKX8h4oQsjhfOxXMg8l5
HOl3nnjYf/2GPTM2HWplbqqBmvtTUFgC2ITDcoViVb9Uq1+ArtfiF+btBVN6cA1mDAfXJj+K9YT1
3BP3WZoPg/rPzLJZv6eucTx4ScSg5WkySRLErPh47WBc40ZiZxvu8sE/I0wKA4FbgvoXf53CVtid
cSX71UlL0RFPPlfOALmoDm4Gl2fGZFn14h/Tz/yxBQF5x9DOrhYvzVO6mh2piqUIESu3YjyF2hRx
CNgkGfCvqNZEOgA/O287KenId6+Ixc7WNRfHIGjkqFFub+ExMjOInSpPmm3V/PIvy0WeFQoVeZE/
oMhcDkEf/WT/14BFUt0iXPkaZPD1641Q+5IEAdWqP0/3I8W6K5JcWDmctEfvm8QKzOMhIL8l2hKw
oPTlRlRPgUB6bFU26ikS9uzR12RxnwleiYoxqlZ5Uz182R85n2ZJSNuMc8LIhwaeGHCx4/yp+ZCD
HIqdnq8vOZa2mqiYcySn+QobGOjRWSpyjm9ho+CRJVMlnpT2fHmgyeDdjxunP9RIPxEvNhxqe/F9
pyAipRepJ8oU9xaHgMTRf+qmXmK7JkOcYu2/qUQaAeF4YM0H38MX/OaHNo4J4Ooe8foaiV8uf2Mk
DxQXEVSZR8kvWgOLCYD9cphhfbDJYiuEoNylqpQBV9IzrmTEL1kiGA5GD3K7gz+u8YyHnL69Yybr
vQOMcbrfMHqt2JG9dw8ZH8set3ANGLYK4AcvvcsCTchm3al3di4CDpCGiZEWPwbKI/Px2CwhvX4t
u0N2Bp9Bh+m6i3G0gdrrLceUHr2WXOH4ZjIfvjTDqT8WS9+0YQDMEIKPPFTndjsFJ8QzvZVe5esI
0n55g0kphUPqEwL9TmfjxW22Nub+RybD++3OxpdKzLZMHfmNdaP0/CtEQUK5tUUuRdarR1bWkRw6
QZAzP47SLz/r9qLd4MxNzVTK9jxhq5uNbNdB7ooiGwD1HPXAN+j5EwwPFrJdSVSnOwMQCeznwvcZ
sqJJGpQs36SAguvTVB+cx92JMl7qFfoZnk5KFs+7sOSDlCTlnY1jRw6f80WZYla/9d4l025/Ruzq
OhBYydRh8gtDw7b9ivamaWbwDaWqPAlyADgbNIuqUAhLsX1WVe4MS11Dt5/inRo7Cqe6yCaOFujN
XRKGeTqLiHehctBVGvS9lw8yRvEsElGtJn8D0d+J28M7AS7XbWTCxR2dENhUu8FdT8LRz91085/1
pjfnYB8p4m7fRNji26ybRTFTTDk29HNfwkRhedYzPqE7vdDUB16nKphG9/orahHWh4UWAQOTGWZ1
EwflnBhULKvLhzrSS3sBvEpb8wcYnwhN7T+Ickt5F6HfWMuO7xEOGvkvSMePQSjqijeZVoLXANdm
XDMRKHQMtnVV1k/8W/WQLQy88K30f9v/wAANVJ76+sUrM949Fm7+dhyThydYg1SJflWyeMa+D/QJ
x9um5eWnxaIrEgzaHkV+yShSKRD+ugfi0EZx03WW+cXxgQQ7R5dmhkWaJ3OJZnQRNuyNC6kUjZBM
NmrC5k+7VgvvFektxkLtOKd5eR0HpOmCa8mOSMP2FU4kYI8QIZvzR6LjbYBpqk8ZvnsHWbW7O8S5
KGgKEBa+kr6dfkMwGO6yX5OxDNP/WBja9+7lC3t3nr1TeLdzdlVTb4Vme/ZIxJzdth6TGTki0Bpi
xA5qGq+gs1PajJlSYpzbUWU7DS7/3swvHHMQpy3BSADYbLJpNH0ZV9v7kr4o1V5mIGwBI/HpVT6X
7w2wiAl7RVatM07en18nQwhsVAAwUWeYORpL34J02flHGASkEie/nxR/3BQT/BgGdd6EQtiFAzbp
MnZO4pzwuTioHK95GB/H3GAM13RqhzkTBhiTvH9YHP+g/nOFijbu9ceFWaTXaNgcqkW97IUSbC6n
p/x53GBjiV96izR25W5jBpFga7Y+/umFiI0I+defmlM1rfsYcpt/0MMIaqRoZfNp7SstMIaN0Fv8
FfU3ySDwrywgG/HSBG43hA51O85OlkdgjXnWJ+rOznqZ/cYP4zbv3nzqE3pbyWm2/PLCDd1Ea331
ohn2I9C2aXWV6ewYcEO7zAbVQ/NxmNs/1wY9+lqS6OpSWrCOT2tWYGxYYhmt9btDgxJaBOF37Mcj
SVj7XVqs+qArtlWSwotQXnsUlAT39WjM9Gu7KDwYU/fWAdbrHPzKkmZlnaOraWwsB5/saui451li
ObEViETBVn+GbfmzOzSAn8/984u7i4lT5dwGj0xPAJUwEmYo4LvFh+hFs6p6pe1BOikwvgb1KZl/
5NAwgIQWiqnXSfJx2+8bWaFL0ArUGGiMxLt8/qjQv7/vvI5LBLt/FaSUNCRicG/GsLTCvZRMAaqN
418rr2GIA5dcwFpfWKoB+dega4ZucotFpEfWrNB5SN8/ByXrfusT7Iu2DFNUgzgtGjaLVNenvpkG
kMHPIHLAZDhnbigBQ8/XNzJtVJD9YgBkU5L0fRuCsZEvtfVtMjtYg6SIyZZe0JmmK7tCaCkPgrMD
Mq4pOxL3Fs48g5Hl3Xx++ei/33TSP4yQ9/WhDFbvACxTJpLKVySZy4nLycw4xw42oTcWJL8GO/WK
G8t5uXYbIwtcGG9YFlzpF4RTLu0J4uIecfZF1WuHzg0SyGXJJFDXjFRI5W6fMrVcSPNwIYdTopkN
fuZLPNHFVCTfOK/yn7GsCG3xXAvpGVg8OF9CfPehuSLSl6tqv4jDB6kjTJdmvKthqpfOOvRK6eP0
TKQYdNqzjV1B6H0GyeBgPpjDVCoMDaRNdGfnauiczBCnYLmVLyb5KwLGk0x//xBZrIbN3VaShw+9
6jKHESuNuUmtYhb+4I9FXpQYTxPHehdCJc8EEr+mN146zn1K64FVFsVN+JgASCoFxzOYofOVp5CE
dO8vw2hGyUzTUJvRVJ9Y4C7lDE6qj7PmPTl1PH/dFhyM1xA/mr1uUKcxiVP7Kx22RpfDdZc4dDX0
agw2ujS+pI7ACa23LoZnpkGwZdJRBtBhlcbkR8UTbMWFNnXdTFARvr84IUxqJQn+8zVmTRUPIuWJ
SIVQ2JJ94gefXDMUGcfoS+Pv6WOugikyla+k4V46gbKmEd0Oy+oHda/bT1PSO5ZWaHb38DYzxJE6
OndhMkVfCFmO4XwOwSxBVWCKDqwQIw6zu/pPfWmecStBPU30VdJ0QeTns3Dwgr9JTIfaiTHf1hUl
Q5G+bIrjnnm6xAdhIaDZUUFCawEHBRj1/nSezzJG3AczBXZwQe7XC2BjN/jjuu/jsfDRv/Xtr66N
2H0O5je7dVkTUAmIGyO5C6oDEF31VRZtk70tVLwZiRcPJxdK0AS/4UKgV05EPRqi57AKAJR8J7uq
D9Bq3JWLYQ3hLunOeSX3KkblvCpiCaptmBr+fDz7gMhc2pMsY8ununfYbb3yJgi9ikmB0O63hgTB
cfuok3MhrL79pDe3UdZzL4fblj+xmry2TnrsrOBw6eMnVODLavgm9xVBpI/60BxEHyaZvcUmUW5W
3OEOGwxHbn5haBVqAXVqChevbmEGDGRgPQoPU4ZArx4/T5+SpEmGRg2TUo0lHzHQG4Pcw1l2vEir
hYQEblO+bmY8WCvVkpkAgjC1Bpc3EXJYisfXd5oyU6drWUxZgd/VlUKj5b6qxdto2jwjpAylq+l+
LDz/sWb51piuKljBVD1OdWjjLA+8QgizZ3ldJTcJUUHfZhL1QejtuPb0+Z1QU59M1jJgxn4nZuqz
l5/jjMHufYOXhEupLvnzvVnEb12n3vhwnFWC+55go0L2M130kPPEDDlKTrEp+OsiE0K7T217qJqZ
467QTNbOi4BfKLP1sBhfTfZwJcNTn1/jz5v5sQqWqoSZUCVpIjcWEzVCbZY+7i5T5/5u4zB6b6QS
/uXEqsTnz/3l/CMUXHd2M/xXIgVF/41I/GV0l/zsxppTjlM2fZCyi9NmwLDhhFPyzFl05UaIDTG1
/3fVZb7mJUNzGtcKCfi1nYNlYGVpMRobXpk6LowD/zDwOq4EGZNLUH3JFdofvlNjgutizSn+rfKK
BBTuzJXCFRBW7/8P6mrT+g1GJeNMFxN/9tZdb8L3HTMNueC8vhKJyhfNP2pgacSB+gZ/YU1sjR6j
Ta6qROWqFE6H+Oi273geVhoUxDiR3OzV4iLZNtPCjlLiKQGtdeNDwlzG2SJm1ozaO2lREXBN4f3n
vEWaH9gsKQGzewIQL/4uIqs4mlGdgFTp3WpTshIm5We+Q5GVUOdEoCUgqxEnZ+EGFF5eObY5W+0m
U+/LbiL2VILQIQRXNqWBWZJFMu5xj0xX+bOkhHzOurbPUTz7Fg/DTYhr1rBFKX1I0y1GcC3KCuBH
+DsodcqI+N+iWp+VcDeAu78qfbloPQ1uZTQK3P+qbIDT85+7s2h0M3Cibkl22DVm/KUQ1Ir5HkOo
7xC/Ym3iXJpyOdR4A8jFxs2TYnTtXJepTmFgpemEcg0q7V5G6UkmzdQhRFM325NUGgUu93B0t+l1
pKFIpsicst47hUaJVDYRVAdUvTGJXgAbKJ0xy/EtpbPknOi61VFsDtpd07zOfFAA7DyX7CPG6Ibt
HUT+CDl0F7X0BMOkF9O89KOm0c8I2MS2QMVWhOUfclx7n9tJ3NnIj9YdycRad8zBIyhuJQUhCB1U
ffA1uMQ9k0GVId9a29uOYt0+3JFrNs0i3rInjwOFH4/YynJXmm5fLavf4hpBakCHt0/e47+ztixI
nXy50nevb9Z5te6DsffyKbgv8qWrcwN6E8pXYE98tKiPzB17qGOkj1tNhaDPIh+EWqhJ6iGEtwUu
RbqSDRbpwGvd/h3TrMge7F6pZQryrPl7OGzvqctOcCoLMSnpSyDP4YV3Ei1VpxfAwN+YJ1Q3Q3Xm
lXLoIZYR5u5mTYP1dwwdVfCScfgVIWgqGUt64oDxKlCh/PKrzJ8xjUXYlb1SBF/+7x6B3bnU1YMS
3zXwY94dVfz+bWYi6QZzU9JknqbvoyAVfIJO9Deavh6JuVBJuCCKdoo24SLg+7oBlVv32ok8YJ2K
WXAiXr7noM6sitYVnLrMGfMV23/KSFUWtpJP5PbdlwTpG0YLcK3HxP0GNWaqxwwICSCg9TXsRexP
4r69xG3nP9N9PckCZofGTgBNjsRZ+vIl3+olE1p4d26AdN5eRVi/uXZqOFijzFAxv8L8Rem7dguY
vI0dUsvVY4KpyR7ifIwH293tHMrBfFiGx8Xh49Bu5RHANBUkStURgLNj8A1CZQvD7Fgv03DLgrWS
HjOaiw1dg2M5tR4uLitEafnMwDSbNvHkXwXgNQruC8jXZoCIVqofdlS1Sk6N+sbHXwootKjBNmcU
dV0f17uRPjXFpyO/xDUCQqSCmu982jCuGwTIynD3GEVlmSGECeLfN0fQpQvQoJtyAXZVLOEgoSMy
fpccCHAoEiDxuuWoBN0Ib3LVcDJtG374akn0lvJ+JibVnM4INZgd39HqOjm4KdUjjZJs4pw6YZF3
6G8PAmZ3VKbIjkrW0aLNnkzOwSJ5ATapya+cH/orWnkmpNJo9d710de8dWKuPWfu5zOxnzr1tav+
4JCkKztaotYkM58Twrokb8vGnT96uvglkgeTenK3njhZTl9mZrxYt4WXDRKwLNBJdMu8fvsl4GrT
SuLffeKKi3G5E6P2u8e16hnAV3ymaqAx+z6khyGwUULq9NiLDDPx01e8EzZDU9WNQKFMXdPnvDiA
BcjToLNC3ZyGWbLBrlOFtDfdEJwM5h/zCyXSaRyn+iryJDYOc8mEPMAp32MB6sOXSjh0DtROIIQZ
MhoFwsQ02YW0ttZpX3pdsNgcEgwLeoNcsk1VfVm7NZwbZa5V+wYylZqYVPceOgDDb3fDcxVxzHn6
yrq3Di9XSU3G++sg/0pX/2pck0JxoxjPiK3MW2zNJsmfO/ZRTfmGWPUyR7tcR/DGLxbqQNXnciYb
cBk/1Sf9UE0yHl3lXgMI47uzmEUZONjEmOu4UexbaaPRL/cT3LsqCG00uK2rBHZrX3NY9C9Yqr2w
iYVHQ+KuDkkv/oVlaTjw7dQ4LSfmSVAXiPX69zaFj4hP6qFSu+21yY7pAUVYO5ubDF4bTcGcbbiR
27Reo/FLp5BPWEY++fl7uSvfqKVT4YnBocm2+lt6mg6jQyS/qLaF8eJkLldBTZ5QLAx8/lPlaW5e
es49+tnUN3boJQv7cMytU3//Ky1WpqqASgJMaH1MuaG/b27wxKCtnahRsgfedZMUMH+0WQr+pmNA
spHhmsaicOrEmAeJyDomMXmmuRPrbltBxg1z18kV4osGVDtLBFF1+nElujM8JPQQkAwRrgXVY/vo
6MtBcR0xn7E0NJt0fbe49/GbLCjZ/AbQQWIAUH/j5W/SCovPU8O6tey/RETe/z3ak7//4J1Rhai8
BtY6oYwLpC4TMjq24LCNNUbuwF6wFBuLbTi488MJ/srC8oQlJGJGejlUWVWoLlabbsX3YWVVApav
vxUtVf7h1hW7PD7ffL2rhVujbcu7RdwFPUJ9KpM2gA+a7heJBnXPCTmkU6TMkhVwCNCSEfZbSLUJ
U/v+wQ2OEj7ig+UYdo+bqBLe+VIcOjjoG3DS8cFfM+Z6o3ZG7rjlZKN9VxSfkE3wj+67UYadVeXn
5GZdp/cnj1kp5RyE1HC5mohxpxkBe1ElTaH+BA9UgBGPmhW/sH/hzH6Q9TO08HJ1Yc9JFnwjozZh
ruZh3aW8B6fdD2JLGohOLhyjZsLPaCziEk4v9GawiLuyc1Sa/rEGg0lMW7V+k97njDXoHYAXzGJB
1K37vJ7vBouzKETclCLsvjsgEY4wU32/XcavefTLRflwWVS0yD92Ev42oR2o5NYzyESjrUo3fwHa
e4qzOfALs4SrOyd1FEG+igL/ybONR5itKiG1GipTM58W+ZtfBwD0dkzyRFeKvkqG7S5DSe5H5id9
NNm3PrH78os86OLBwDmVg+ByF66M0sVqSUZA51mwFpZIXvDb5LHG5cmugqnCah91bFUn8mDnuQPd
NLXFzyKTX41zHSfwer1aWKOgAF/KZnp9EPylGM4UjpAgL4B7DpYS1/GDdfEkueeHLuWF5MHzSdwK
6YboQK+pEZ21pILi0DViWbDQ4wM+hNGik2S4WdQo9qUJXggAXCSGmB5pZTjlJvp94Jkh9zu1fzio
Lk26h+yOMjEYPs+KvmBDOgzDcEzUkSSA8sJ5KXMRRGzezFasyOUYu2QrWnG2uls/U1ktRfOwHCBu
gZz3g7+pDX2CCfOiINiqEO0UbrdmzANUAvK22Z/yw11dW4hpdvoO8ds8CDkvzPKArnpC+kfLhm5L
CPVcw+Gcex4s8tlg1+o4v9/JJ+kLjSA/cS1qHbq0pW0lnfE/rk50in2mRJqxC/21Uuku688pvbm/
9Fa4DrcTmXxvVp9+4wG1ffH/6v8X64UBVAhSdbdhr0GeqXklR3n67RuuZtVryUjNcHp0UoqYzziG
le8UMaobWPiKXX8hiT4YZ4CPCDhpJOru5EDdiQDnKB5F2PhEYDMo9llYLYorfJXAsyZ5cD7Bm2YP
xaAEN5qNxBoQERbLPENadF+6byCgPGgBmusZkDjl0gzZRmQ1F9yeS7UhVfkJWs+C4tyhVQCQXC1Q
hOoRIF1Pmg3UC5QyfrxItEqFXh0X+iKodKVK6tbr25SrNI35Is8ydbsKwbeKQCLAae0CB1OWZGB7
61Ffo2+SkMwjXNYqkD3MZlwXNxkbmZGxcjDbI3tpjBDTQEdZGToFIXTzkvAMSHWphsB8Bz1GrW65
sPn01FU7g4EegI/pt5vaL1xPjqjiR0py09f5vzi4Guss7X3O7Q5ZjSUJvBSTlvmaB5JtxW20mNA7
wJPkR8zJr4pRyZLJcubmY7gYoTJ+DKuISEgxSOB/R0QkEL8bqX77NQqEoYHOajnIDJSA4eS3UH3S
mPukW0BRLsYOaK2TWQhbdsMcUrZpgDdT7qFxLPoAeqwOwIbww1slQM0pVaaiwpWI9/K8lu7tCnRr
G9B898zu0FwSQ0CXd9MQ9dnXCWJ0oDlMYQs9jbBClaQPpGzfR2BHup0fMlBCDtRQwV0BV6fFMUmL
ZddcohLypufOIaPz1iRKeR9e+8WdjqHYP4PGElX7QJDIqfjFrFyC7Soc2TY7QI5Ox9ZYzPdHaasx
Q9K/lJdQ7sKL05Zxbf8v4k8/z+riHyYBFShVkJVgValW3aNrQIA/v3+eWyChKq/T4oxCP9f8AkQm
AbbovmNlkQuJprrugV+alqGna9Ub3m68vDmTmuP9DMZeez+6G+OkUzJbP8csCKfEd5CMMWpS1nOF
aY8sXyuxgFqzENzW8HWE+x0dW4e4n4R8aSocPxi7fcHPkXchCbwXUEUtDyw/duT7UKK9x4GVMSSZ
UKpOTD4SVGIvKxVMWfwywQ0z9fG4ArtFp6SacpBn5Yl3dcEvi6d9KFALrBmKIJXcxGzH4XD6XGAx
ILRWgR0a2HyZuxibBQlAKWXGnvkedGhjv4ikwyYYG41LCHawB0fTqCk6B3womcwTjLftqj8HqVx+
FYfm9qZmlqFK4insKubb8Ndr1PkNLj2xIA+j5LAIoI704p817XPVlZO4F0nnFESvrUgXRBvOQYzM
lazAcemkq8WmbtKf7czX4Jq0euZAbMZKBkJuy3SVoES1hqB/bFNwdmCwWayhpUTbeeHFXu0bvCsg
Ue70LrYF8YYJIJfJen7D9DzQdgjlfB5gWe9kxzshuvH1uEKFPNwQFqirQN8BCn1+xCWfOlfXGb3k
KLX3FLBr4nFbMfkK7IdF9fdnu7FHzkCPPgT3+JGQdbq3UETrpmAgVwdDWBz5qMKWShY0b2YcowUX
1+j4Il0jfKupL2qAcQw82HXIZXa3ga5879e2sB2b/2IxiNPSgqe+WdZANzx2Qr2UbKNwTTvOxIti
cUehJzzVK1UJ3imtwBKPUb87fU0yH9iqhE1YC1n9VCZve4mAi4xDyUPjH03eFvuGg58s9YDAgOXb
RXebMDw774eFvpB+9TFE/8W04sDeXcGUXI7ETIpBNoxqAD58CUxR3KPOQmFdvHrVCUoHIbGcFGdI
3Mf4EuGoaPsyxcyfRmkv5FMwZNugrl/wQE0UVFknQhyL0E0hosKz/AXDmNJnfyvJIdNSuGbWLghG
PC9V5ingb6ogRIPmPIOMev+XrE74dXyJACoUdZDB+sdORMiNqORMa95aj1MDo6wPlYcRDRj59gFL
hqaRlnb5wmsNPCEVJbshzOiJTwI+vfwQzKoqtKOOYvPqQzw+m/ZiQo10XomfVWfBbt1/bgiK1Lr6
82E68QSflQybrIHp4coQalEnJABacquxhOl2JtG3uqhL5kmM5Qc2yVQiHYetQanPHuU55Z7/wPEk
ReTgycYjJ9pLyTZbhbI6t9MGGYMGND+zawSmsHOhpkLXAYChthKlVvtVEkUSnMB8DLXFJa5sXkoZ
IiDUoGvtRf5OmYFZaa2Za+ZMcUJun4uI9tQ9ApOeAxNuGznBXoDCRO/i5LJ31upKHKYvlH/9u3BR
f6udgEven2g8PDNHYySw9ijFs0RfplPqAl/XEbR8UHGS4szVdJDYTK3jpSsYSjMrno0ycoyaNCtb
cDiQ686LC3b1WeggCwaiANVp59HsCBLsxECcmP3pIgxLjz2/4DAkWtXuNJpIHWcq+ZH+CwVg4+Yk
4EIv+fuRl4IIA49IZpy6lu0asSxfkqiXLTcO7fOptxl0KdTnj0ENG/mOGhGe8UqsGoBPE0VVVe88
jKRbNv8r0OeSAk8KuABKo20TmI+DMKKOBBxLS9Vks1mqPT/FdGndqhrfyAWGDBKScc82J0HWLOsW
IQvq2waD/9PBlOQ26pLWLCfdHY6IXZjJl/kKmEh+UQ1JWBpM2MIlf9VTBOCva0Z4NSOMre5D6lES
S/xEScaarcFRkubZizctBchRZgRBzclE9AudxmLsZ9P8lERBoJQxBsS2duuZC9NSCi35WgvXaaWV
hdI8wGCUcQhliWfJwXu3LWOaUNNYX9xSRrEAcctSqjrWLvSSYeinQ0FovlO8B3+PHt8kAmZPyy0V
aL0/Q7AG7Ik407BvgHPE1Yz1UII6CHDtyi91HWVV4/N4Ej/znA5sZxAYzbtP4bqYwUR5XhbRYmJc
VCaLusr0x19PnldRv5LFTCWLq5LUxWqomoH4oA9OOGF9vrz7h9VPoVkuTiUT3VOKu7phadkb/4ra
pRbrWLNzC8o8dpaAReGLty2G3E4466V63TWOD/k3Z/yBtpziteBOXmIj9qx1q6aZsT4C/KvXgzBv
KMu2q9ikCP1eqewIh+jcsxgfOMBh+qw3vHA0XaNtHxGL6HNpYwUEFRMbMiHlkDQcfq2aHCSUF1M4
cnTopanXTM/kf9++zHPWpson5wOFqUv1DIkAylFj4P3ndtQce2BrBzttdOeVlh9yqECGEUK7/KX3
uZyHQFFKbRZ/S7G5huaY6KRQaFBgm90fP/2b2Pjj1BB/qAs6SqVtN7YJH/i0b2zSGahLWzfEYHAl
BLY82I+/didOUo40eFsqmAR5l9zfxIb59UzufRVY2ZZw1K2cwOiNfWurb2UPcasqV5b7ywb6r3X4
wt9WcwrkDCiuMbwJ31mrjBd8+TBEFDXJGC3Dw9y9cG39E5nF0nqHFiVdu6farEKtovZ5Hp9fdxfb
9nmiGZPAy+qJjiY9SM07DmSl1i+zKEACZPvqI4Yaj5UwCI89XVjNayt3iLROO63NqucQTYYgqF/X
qBUGSsaHOz4HcQUxJdCsmgsBOnf9AtH/a7Yma8CVVeQhulTE6EsTCNKgTUoc3jAW4/fjnNbw48CM
TaGlorra0tQDdM2FEH1JqWnPpmzkKLdqJ//2Hp6k6vyVYir3rb+Pqbp8Vc92iRu0YPx8cz/FYEoy
M7dgIxurU/hofmot9y+xePjvKIDMIzIZNjVGRN+rZZrEQ8eNkKZ24+311L7/tkIi8v6LeZP2OH6u
e2DXxP82EZ+p95TOof7vWP+/aR2it6APIMBKhKWeW6yL8R9m2zwpUWhJXmWS99lGii0pP+OgLukd
1LWvt/tylSf3vO+W39k2TXL2ty++FBXJns9PWQp1L14YW41wiv/YTh+ynCuqNqnQKoGnmGBGe3Fi
jM7iCZE6hti/KRbqUDBK/54ZWYNW7o0J0fszIA7vudnkR4Uh7CzNGQZlJWM4YPSbmZT0xQ7O0sf/
CtsxQ6y0vmsPlCh/sRq58PqZQqi7EEXWyCMpUXTjXdK723qFaj2YUekA8uat79LZHcujNXEPNAE6
xOdiiJiNWVcNgGr8RCY6C61DVeAlnprmGra+mIScGTI/KsmCo7bTkaz1+Res7I76oNfs8+zmXmPF
dYUFEcdcJNIiQfaanKn71Uym4r04sCMKCwI6u19wEbDbiqxVxC/onm2ufRbliGi/xpaP/ypiBMBy
2zD3tcrHBl8XXbPMmuYjTrdIZZ1zNT0sf2GKCV1Dd7WRdT/oz9sIhKAmQDE/pHuAZNDblR2kFwwS
Z82xgSd5sJifGvbHk9PLTa7mIyD7BH2ITHxTDTUrWQlzgO8K9pwBmd1Wt5X3BsnZw01WUGvObSfQ
wrN8uRN0PjH7OZjj2UvCig5tN0MrwD0LVrEjsTQ19jlK7AATc/3slfQ2LET6Of9pfHvkbPjqzoGF
Jb9Ahwx9NNS3OvRaOkFVCna4D1KAUGTwQB/2A9pYp6myYS1g58JmY6SS8EEkDoBGEBq3DW2ErmU2
oZ30rZnJwJczeoKQbbAba0S5+6kdTEADgEIaqtCj5chIBvKIj+pGrzYARus74CNWdARk51zn1N9j
jIF/3aN+ox3PldeUWlIbzl2SYmwKcyYwdDMY4oCzQg2ZH2q6/s3o5JG5unoButqsGsIfP4RBP4xn
ztxhM6SWgXjo7V8YPlAerAD8piUuSOuNrQkktGssAVwWg0cM2CQjutK1SmuW/nnoaFJVkixjK14S
XfrTEUVHS6BhDEsHERtToiuuEP0qiSe3Xzy/w9Og7PX0TclkafpHwdCUZDbn9T4QaMuhY9Gr9nwF
r8GMaKf/0d4d6VUj5QyuIxiKALd33Ea71YgcJQRvxIlytVpySvuoGZNUv6YMwK7p0I2G7kaGeNTf
CSMASD3RCCww2bx39Zl++6QZ6v9Dxlg2JqKRUKwSwA8ELRu8PKqT1C5OW+GVQfmyaGBJRV7mHA+t
DHjaREbZFSjmubNgjXBiZluJhLWCPjgKDKy9STpczD4VxFauZG5D6DIFtmt82t2n8jpBFUNe9p8K
TIeDEULXmnzi+2q+swm8qsmBGqm4BvW5Qb7yBbE+iTlKnysVmhSe9H4w+lxiPHBk/T+2n6iyVLD4
kNxO5e8t+aH6yazsNK13GTyrXtlaWVGSKTzlKUeYCqsqCqJb6ZZri4Tc6Bkn/CPIWlr/l3iqPu/u
FvhrMHwEHmCvL2RFRCJDTV3CJSDQo3J5sMbqCVZQwyUGfzuOe9Bfvj+jE/v5nkFZAXEQSSflCb/8
ji+URf5owFCM74seZVxTRg72qhK/gwtIPL4WHbnIRrJMcCzolOS6rQTkyHar9f1kkUNvH16SCGz1
arS+0qz+VXqD5acmwT0OeM22n21iTzQmZ2VzYl0AAAYKBv5yz3Y55y/YSU0gRVmtKjpCfLBMNXNy
o5mGO6cIbtiSxNlZCFGBs6N+shIzjtt21CoKLiR9EoOo/SXCj0Oc/0/oq4B3iGauzxvMRLFRkdwR
sUkQXAKBuv1SJ3rAOgoag4NEfQaNxTbOBanC7oQBE0jjfRbmprw0ZoijNiaK16oXiGT7KlriXpR0
2W0yxrCa8VfG1xWvT/AWflJPY5HWOUnkxiq8FeR8/WLpANyMxXoZDO0dSMAAeV+iTYDjCaqFDSZP
X2HtQ81ePimPcuktcOy8TkCuh8zO7xzVxsy8d/SDs0YXzW/0zxUNs2pbAo8xBsrq8T+pXkBzQKDB
QajMQ1NOJnMJ3T7Lvi4FkJrrTHswtX9mUS7li+tP4quVbdKWlPf9tlr/NeKSF/XRONpVJyy2gE5D
b50b+ajVfsErW5wD3Iu5V+IoK3SRvRus+U0T/lDtFFA8113xag4XqQiQwUgS5Xlmmqte+xt1G8MV
eHXsuYihcpifdUKXy6GWZPDINTAJnglXDx7cXAgdlr+GFezmxxuCq2rflQ+uoZPVuxA0ewtxDR7c
E8AHq3LC/N4Do9aRofODxbBF1hh0xvR3Zfc+d8JldnnvGPWYNqBxqal8EQiHze77aJBziYtC1JSp
UhT03Hgk/5bg688L+gd5R5Un/JfmEi5sog28M/B4tIxt/QLcm5vZWOZ/vwrh84CragFS7M1jD9li
kryZsFmFqIUBLgOP2feDCK17Ed/w28rre0j/CE75Lm//MNBIxx3yyOF5HDhaAuJgOI1Icjg8aVZv
Gt6j9InBXT7JEM/29n7pZ6RfVKoxiNYseLiLw2NdL4fBlDNZoiTUwi0UvEygtUF/zJQ46ZP9OdXC
maLL+RddaSZBEjPp4b3kmu0SULbncvBWH9VC4J2l8JIJ+Vdb95Bmsa1J/UdGEuH02Leg2yVgvFyx
rVeEUp7e50BdFu0sG49aZwFYLXVHQ97GIpWXepgChwNOFSr+hMERpj4nzIWawpzm88APgrI8yNC3
H4IKqSH8p3QnmhW8axpT83yAeNpoZGqPQvp/lrxTYLyIMmxowoRshH3hv1m1BZbLO8ZsxQzPAVih
WuQaucWD8I8BxQioERK2RrtHPxhFshE0VQIw5pNUSGu+tPOK++QHSyrxlxsiLW/YvQkKU9CfOrG0
TMhfDzm6VihfLaWWF4mqbv0yFH5DJet0CzaLahym0/prNoYLMLQHQgQZFAUaTZ6XBYRygFRWTKcd
FFWQ6oIEXg/XmHbIEHEDqESng3QqiDsKYL0vH9Qc3xz6hQgUekaKvsHqtbhBqf+uKoMC4CFIZ9Ag
lKDfsM+prAACcsC340YhS/dpX6Kk1zkGJes+ixv6rtIxa+25Cg7C7Ux2cjqG3ZYn/p0PIUtwLtOe
9bG/9uM9JYreCCLF2Qi6hA1B+G4yqAZkclqamrRhfiW59r5U4fFv9USamGlq9fGKXOxkimHOVjl4
gUIGnIRKx/S6r/YGOD9pjqtaU4JW8AKRzg5EDnigyXlJzYCB7SP6+YA0GhgAl4yEGXP/nVKnoofm
7PURyZ0MXRh73UW9AA3bWz2Kygkv71FFCXXLNTHVM7R0rdZjAsVX7zj8YMw5oxQGRO22ZyxRfH+n
kLWC1nESRdDB5VGQPmJ73kg+rR6PBgv+SC591oIs1hmoROAosRs5er6bVko/fCIb3F6lMwRW2muM
Fx6d11u4uq3U+8ks+D6TavkSJeTsMKK0NdLjX29QCpLO1qEMXbS8eyEkjZt7/kUgsG/e7kQ1wGOi
hpPWNgoS3gnAGPbWTOY9ZvY+QXqRV4JCLCIDT3aRry00k9pBPzESCYpWuO9ZLFSjddtD6ofwBFnf
KrgBEY6Jx85p7QwSYKDqm55LYrzwjOf8p9MP1sTwsTjW0EplqHFlY6OIPaI6fNw9FLwPxwy2myRh
eDjA1TnMNhTGecVtA9mIqdCwndx37mjj18dKXMh9zokgNfox5Knal2XfrM4LdFXTol0URCFigQzf
Rd9mW4RY5VLTvezDpCQwtYsPXvfST9UAvfwY7v3vblfEY3VSxGCl2WeW8IqRSGgTj2x+4t8WXCwL
To/dTDPhwVQhTvpkyAGlMZFDk2+ZXOhPcvU540IqcBigdddbdKWgfNV4Wq4VszcRlZqOZSQzBKn4
aZ680kIsoNgYpKfUQnvdgOwPtkl58E55z6jnOqvrU6/8hP0TcDZXoZBYK1hjKDfX/SFgnDxx+yHR
kDJXIXHbeCgc0KUQZyL2Fkr2pwqLi91dTsRL9QarkgeQXs4WnSx12PHCRuyDKX1BRPj+cIAj8Ywc
5hLt+mENLi/IIoTV0CqkBWRknyR5UwC/59HrUqvQbrjpHP+l3b5w7CgsiP/Thybqd47w6WG92agE
c2F2xLHgjXPzgb5fMWw1TrMgjAcnszXlklZcb0lKcZ/xiKXlTNxqNFEHbIoM2ExV4jJLPvWWJFxO
yTdto8G2OWbnHzMDx7pFw4vv+6W3kRciYCt8JmHRy4Cu6boHrjV8PvC6+PGPWVyn0yfw5pAdOwUu
/HpDG4nYynDpeq/ky1ox3Jh1O1Zw8Jv9csWmBrbjwrMtDAnL0HbK4SJyfukvjwbrDv8dd/HUqiUs
N38BhMk5w6p5mgxiLwIowOb0l0oV7ytnZr2+ZzXctjr4xewYnhWN2jExr7l5Ga6AO8zX2fsEnSm1
n9eP4EZqdDCePpibWAJ3Dv6Ze5A8grR+TK1u7j/om/cDxTuHCo/0eL+gXOYWFDgcvjelDGqOrwdy
Plg/XJrghdYTWZTCeA9e+uPTbd+h8ovIPAjyl/CElEdgJWxaneUUs56INXK1b5/muYXsdUESnNYk
LbAPlb0urMEoUlUjytuUzY3u84wl93W3SO6jAvOJebtMKiNtT9CL6xrz5fzJM1CbwH0GQ2cEPNZR
bbdyirnv4OmE+ZUKqHv1EtvXJxUuPkNAnt5T5ut5avKK+bHSsT8eV3/ZhVnP48Z5qyjRsnh8V0mp
f9U+kPGcln61RAKPxv01JEc50DOyyvJMZ+f8mF3owFVFqE4Q5XonYiQhsrq4pALPoFBGKo0OUsjC
lU9SN7bqOBQNPZz8HrNW59SalT9O1dV/HPvp3ZDs3Mauo1zqwvTdAFfoqem144TAEXa2CEjFRTdp
45kxRjLX8wrnm/E7eK1fExOZTOnpVS4X5Cg6iz/dh/ID2YhvujOIC+Cr3MAGT6FowlTsgrE10M63
zKlcfdsROXb8MSVkZsLWBhN9QvjENEqW1lxeoHvkj8PelxQ9ypGnIe8TrFiYnZwsXQewvgqFnHJo
UtyHBeGvxHhBUbs7EAcIrbuxB3ROg70PfrT7nCG+1UirlqOJSmlxReojzv1gb1IjtOQrEwIwFAO6
nuHUFYv5pf4GqbIN6xYMUHRR/oggRWAYshhZ6s9DwK5X67q9sNGi0clD99bR91LjZavGj6F8xTry
9TxeTgfkisOtZ8Hn/FqiEYCOpbyVdWdDqW8h4TUWsexkraZiKtBpaeERvq+NKAVRkiVDPUWq9vMw
hHqDH78DVMRWIWbmDsvn0J+l1SQUyATul3vYRovT6xzNiScRlk17b/r4ywpRGwqwTiw/VZbpJfuR
HWWngeqL4rYBTbf9RALCv6kmiIfbl14zIpkyF+72c7yXsA0FYO1UNfbX0g/wWpp9v+OcaKLoYDDC
eOKUHvJJgF3QB6awFs40UZtC374BMwvdWkaGvwPFX1Abh3jqnRywkmqwq//CttDevECSmkvGrCBc
VvB0ZO3WKFS9Rk2ILp2JBdSmTtUbJBp52Yu8gQHcUmV8iH7qYtW8DnDaqMQrNyd1n1DLfi2q450b
Y/Pgy+XOnT/dgw4/1OFCLyITSiYFrpPnTiV2VnTeljXY3WW0CQrY4ncaWGtHquW6zIEhqm18JCnz
9jYliJ5yUdeBz5Q0eov1CAydJ/N5svkOXj+bFy3Pn20/nCFDIi0yQA5BwnRFzJ8Glj7aO7ziM4ZI
FZUtuXbIn6F5Hor0R/kNHNg4xjOhUz7d3jdQzPdTkMXhyCBwCo7EtqNGKw0TEqoR3BlD30saROYR
vTKAYIbPH3J7CsIVpx5kIROFSlRz7kPsCCduotWsuhewvaw1qQbYQnQbQbRWcwVro7+2YZigMASu
1p5laH3bvV7eEDxNkN33GeJBJMQYI3LY/3H24itoaHJSXV6nUo1xzRjkdiS/YeywLQNAsl/YXYhj
o4ARHOGEoQvIf4fYHEgLHuxn5GeH7rSulxdtjpaMCoYIeGaqry2l6rfpR0z+BZzx2PO+SboztypS
aUwchVdb9U797hcLVFsLOK8LUVZPecU3xJkJZyU9RCsguZcicP+vTs+YGXB/OHhFL6zfriVXWcDu
JtuqKdl46ktNymlUh2YvNotTFYv5WG3qb4S/pSR32kEhOFavRF+H+OaAdVyDyUk82dTbqTdME5QX
Jwdp8TBsTqymu7DsXSmfzYKGsqe4kYe5W0YTOM5Rki2RvJxw2o/3YOWF+W1zkPevABONCUNor6MY
/CrleEBp+lq8RfiUdLLsQh1mM2iFp8ca7kXntoSMqUTpwoBiQIjRj/UMg5319UPAKKcsrWUoINci
fFZfnrEgI+zbLL2QqASprX2Ah9nIhkaMsPWJSCCaTwajriMvXVVdM2mkLniHxooRuz/Iw324PUfp
OiYuy7kfOVcYakWQPzthfM2hahBXSCaygPI7Xl9VB+UVDPMjxCFFVxLymASpfHCiA4M2PLhEtGr0
o7JzF5RWCEj5ojRoNwpcWUDKdEaMvbFWNHYd4i89ozVsX/XWpye4BaeKddsoA38c6U1hbvat6neZ
bWjovVoLkhwu/1V1CrZm//ers52fxtAUlj3+9G4ocVVUOgP36XR+pwpfx8FaP1nRNJByErJIB3cm
U9Tj+Pv3Mb6oHYdKi8oHWrSw3INVNnnkgQmAzNlWGUUNdjaf8I4n23lBeFjbaD8mBkdFEiLg1u4G
qWeLa4Eud9ul+EuUAJAZExXKRXQToLfnAuNqzs8+R5hZp4eAUedENOyp+s8JVObdWjDFFw+KEuNF
jio1K2E01/OTlXc6wpFQmFBvPDWDaZCqRYW4q/w7ZUSChMq+HcDqERof7zCSKhble6PfEF4S+ccp
G6sST6aTlWmbA8y0/IOdV/S9hMmDnGT5KZJfOQUWRsrHnBiKLjoj7YcTDzJ4R7cYL5+tGjalXNB/
JKb6n+zof8l0ZlkoJw3vNI3oNaKs5PoZrJe5eKQWENIoT7VBgYsfNPvrYFsjOASs1WB7aU6zrkxI
buzQ1A4iSv1x3gxEpHVScwFCvd9eQxZyeKKw8zaTxJcmxUJQuOUwBuptRLtu6OHslb0UEcMdeEnF
d9/XI80cSAsJNwliZn8oNtTezO+GiTYDaPXuSzkBH4bKAPUGCuXeEk1N8OyCAhr6o8YedBrBiGxd
+Cj68/OuDbvV/eFekbgdrcN1vgTzYswGIh5il93fqKMVFdnsW6vLelhZDdmdKUK/OU+R3uXfUMNJ
tQn5fOPlY4IpGTzh29KfSELtxDRm2t0UfFwmOpliyPNNSY5tYPPB3JzCIRWlx9+FoUQ1371euvDw
e8uFhyfM8rUUxuKoOjTiJmJ4A/ecoGGh1HcZuMmQ5BnMfvaia1TCU6awNRcysiZVayzt9WBcz1zQ
gaYMNNIHqgIFCIhZvAyqUuyPJKNA/fVrhslnnoDgpS9vd0DV80n7mKm3be0NtOSDg84xSugdGtmN
FJyjWt+QsMTyDJPmfR6N9kd0vBemRBVr4+G4ytTJqWY8OeqvaEn19wEZ18sauVCDkpuCX8EaH89J
iX42TlirlFCBcG+8jKOyBqG8lTPkpflfcXy4Hxbb62VjuLfIeEOC+iUwoX0xD+wUqFAB98g8Giwu
Rxj8ON984q9KpD7N0HynD7BW6VaYb+tJBMUSgsCaEIdxeOX5RfIrFmVAcSao882g1T6Jgr0ZsQ0P
iPsSZExpv4z83mQSp4CjnbhbVeWPRJoJYDUt0/TvrrDbS2A7nY9/ynqNv+H/BF71rSowgEhuDETz
L7vZiVBV1XFBLuEY/ADcjQrf8kD+/ZIQYuqD68PTUiyAQn6nvGqUcHyC+Sx5OnVP6SsRyoJBAKJz
z4wleqOtrJ0LRujfLFpQbMsefRSP60+F+buTyH2MjM0kZFVcpQ1A9pl9mebLJdvIbSejgffcfUiW
hcVzR6MrzMVNyEzh0Bjy6qJb84bAt8oeAmbFpepwEbesE53xy8CRNMSSDD/G6p/nZaajuCnKw37O
Yh0MSMWBweLnqmbptOYU4JCNaZl+MEFv8aIXRLrTKFWqyO145UDcOlTmfaRoqworBeSjhFVpQVZq
R+ouU0/wROVoxAfJiWrz+dSZiKe/qnm4JHFE3zQniTviOZ28QHWSbpeBMZ2yvKB0TCrq4yd69w3Z
QXIOCZKqBzACShL/zEvexmvqpuZXpvV6RCkMrNHzq1yQq8eOk36JvaosYsal9hnalQ89omsojOPZ
pdKks56JJ5m1u1X091bDevPJHc6/x63nq8m8mKFUSGo1C/g352DCKLNOy+n3XflAdL8PmEBdZC0N
r8G8bZs8ZNQbOddYbcq8G3Rozo5abipjwNlpGvQIkAp5NiTichM5EFvfF6pZBZ7jXfpdOTW80ThQ
GNTufo8O1/mj4oDIIfS4lHSyj26QzmKVZ/cpN535yYNruRKHaS5z1ZSg59FqHbyMnBuhgsOKlBHb
KtsGx/HeWdvYHAeNKaDN/fCAJNq2vdSYu76Mx+XkvldUOsIJAvtIdG8AIo3PkfyXxNxm6wV3S4hm
vTt9OhOeEMKKGhAvgztLuS+8Ojzop1e/bIeRhsVlPGadTI4VorLkmMXMt8zSeAb1Zovj7CfteRJT
4Nm/MLge7FjSnhxI9kCwMVqpKxOsJ+GUi0V9nW1mcAwt7eep1hLdwt2P1wxEX6a6J4CH/mHUiPB+
Ln6maayQQhVskFjGjOgMuFjtFLp2c0F2EX8PkKQLY58+AKQm248QVPTQqUZ7IFNwDZQZBW89rIT9
23QgUWPtn5Pv+qpFKowLBUrRxW9QFKlZWoHyowkblQzYUrs8QIZ5SEY4NsG2XsUDsTyfkVTQGMKz
vPSCMLZyxMuFOJEyaBNThXk1qLnGU4fEpfYHaVgnJCYpei+eHV4S4smqr3V7/xtgGuTFHtsY5mdi
7h7aPPRYUYghnQfH5Nc7WtcQd2iSd8V7xfIUpd5kNVFBY6ijJjsWj5ymR9hjGUdo73JLLXmp2hqU
HeQ2mQuKbi/OabXc/S1ndsUEjCmd8F/ROPND59abELjYRHohE4QF2cuas3BsCkXc2iw7kKyFQr2t
ZKeGqpnCO23YczLPOUJG9MecrC+XRRlAqCJWVBpB6MKpttJUxP0FmVT5x3MaQaK+fZjk54IIX3qq
X8iy1LJoclL0XLfAXDMiBfvVRtly5YAhr1mlxYjAanT+tFJXb3VAy8oeplbdVarSEAallqPI1X73
Faix8PHdRTGxLRYXNez7fptqYvL2foiUCIWrqfYqTDqX8UEn4VH5Usb6yv2HBvXLIWS/8sl9zz8U
imRYwo38aANHRGRCsS5TfXOk41CXtEORPoIOvWENhuM6caXC5lWQv54/PPpjE5S7SOo7fUPUL3BU
JoO+aHo5uMeLe0d44SRDwZhBqBDYrL65FIpskok8jT9lGdRrqWul+qsyRbHNQJyPOPliIojEAQkL
Uaro20odFuP4S73gWqlOo8ac9tCUYOJTt4rWRRfHuuHAY3l0YSBLkvsDr5qVRm632xhxHpEZhyze
R41v2BMBQilsniMKhNQwpJPgHhL0RhAqoqcoNM1bMm2m0syhVL1eh7kKco4FoWuOdtZlJo89Q6Lj
+mlskKEOtbhykJXqZvAfmGNtYn5ians5LOjRUS3a8QAxk6hmrEJyurdSCT+sCdlBpd7gB1ft0S93
LzxTm9nZ4t6Hvg6B6CKJ3rox0tMycvYGNjfn8UqkwkWx3ni9NbHUyAWCrSXFB7n2f+fRuFiWQNLn
hItF9g1TBU7cWAlpoJIXwJYfq9CaQ5i+2PerYVId2vRAqbLiFzlDgxdmwO+U0m1mjdMjTBP6Sr5P
LdOYfJAXzi+96T+EYlNjMeJEZiGKf6Bm4ZSIUptUeayRt+RcQCOZaOEzBDdhUc4CPeQaSgKliy5u
bT4EJ/l3KRfPY/Wkx4kHyqQdteDfZbi01gSUo2FJ+xx5mKeOjqJZ+42LjFjKwESHETQ3XMeJHdHt
cqgBEi3Ha0OLL5OAhPBEo75RQqMIiA61k3AzyiJ28BK0MXp0dBn+UyuXKj+1+MYI1AU/g7AS+20g
boHagKs5ofjTE5Ka6WjmDqnH8ONRo07rGo//4NBpch9w4op3q2HsJOR61VsLDXZEogdnrDibNo3w
DhdpRM6Fk4NbaX7tAsP6oFTEG5Yw7xjMytWG9tTBWyZwwetIl0/9DfHDIeIKy4ANe7g0QR9f6cqq
WihyQuR0F4pYroYOSGjBa5la4079HiLauc96AKLUI7oMA4KJ12h2Rr8ScwzqEtNruTCpHfCGMTr+
8zH5skcS9NYvvqm8ATAavmuWCOv6cy0sGLSNuU+RF9eVO2xm5l7JeB/23YK8wP8KT4XNFSl0aBbi
xTMD9grkqNii/h7+sD03jHwzVaruX+vkxQ2cydBPjOEWieHOg0dYzJMvxZEgvyVwqh2VDHXVwbwf
Nt3TCyY/masybne1bvhsV34ylPUxPdI6KaSnZSgKxG3bmsIdJhuSaG+JhWkYvypdcdAHADA4ejmp
xb9VhT5kTqqzUdVZce6SKCrLgr4FcXITuIOlcxgo5sgFW9deS+eB0QDUTeSIo9GItBV587aM3U0Q
NbyEgyJBnkUaevA8oHintxp+fA8wnhxboHuKoz6QUWAxxfyNT1v/LJesRhyfMu/A4lfcP7NG8gFW
XVMScNHCZjS/RTiDIlNiIz0SBjhOxOEZCMXX93gnvdqtw9VGKZ1pK7Ls0htcIlLkyRNHZZff4twP
cQY86jQmG3dX6WqN8ZdXseS5bUeRhhh7TU+isaRF1gDDCxawsWf2VmPWzvevMagowpigUdjoP5Lf
iEOPq5wixv5i6oSCNu0Ss35RynoBOOwNP86G9yEr+G5BkZxEjE/ZkVw/G6MtUzXI6Ah/ZTAC2H+X
5wstVhbNaz9ERM1sIgW8iIkWvcXTb77RSZhFpiqhwZt0iht7/IXQIyxOnEBHIwnLMNwyF9Vja6Ou
xlu+xbneq48PccDEkcOBELDeajHPgCJ0gw4JHOKjsOZmbkb2bdZ49GCImFzFsarwo209gt7HSXkA
oY6hTtvJkwiFtcSIizadm6wPX3Sw/EDVK/BbzWsk8FawV53O+Y1VvK/AQ/eND9fwEEZXA5H66H9w
4p3DIlDZYCYDCPonwdE/0eKFwTKU3uI4TvbND3CEHETn14uGSeJmzTlJFVKU1XNhKonZnIQvvly5
Re2DJquAMcpHLZlvlElEEo/+MbcfZuei7WCTAum1nmxo/AzSlLR5iJpUwnTWIoniVweiKZBIjSsB
YQt1yZ3r2V/QVH2OIykOwv01BSFl0w2a+bG1NcMhbj5w6kaBJMnc6sBfqc6Zm42ed8vYbk6dQ4kN
6whuBPHv5NNbshLB9y4A61wDWyODBb+WuQN49NcSzEy3Lvo7DN5VM9qdvcIwL6HzSdfXFkkfW2vf
NIvSBuR+ttd/xxr5S75OmcSWvbHHx7qRsAJE7CEmZXqnL3qPOE3C9m8asx1dhdYIEyNk5feZzoYg
Q+0Nq4TYM9erAxNPd6PguVR2RJ+dSHI5guY125dlTR4mNnBNAEju195wAIKCy2o6da3yU5bqHWBv
SsTXCJxy9iO9+qw0IqqUHw4tGKAgcHVITJHmCq3WdFSQbIrzKb+5WvspajU9volXwHglNt+sdVC2
FY5zCcadoZY/39utVsCJ5aGvfSVwJ3q7kVV0SMcKQm50FAl61GVge7pcyPlEKwPf+L5NIeoRxWS7
USvYfPl+KD/qVQ3jLLAOIwwIXXuvP1yqAH7381II/bgGpPR59w1JIdek1BWyFr6lbdOc+EDjK6xw
C65Pq/vwp9WoMyoYy/fNCTeyYOw4bMfLb6VPx6yMsMVCgw9xO2KVk/s2W+j2XlKVpe2aQ5kf68AP
Jxwpk9FPmk1gsiGG7BEG/ukybmkcyfQVMo1RKxDm3ofAzR5p4szSfiUnV2KTWL7IrijsTHU2Jp5B
QPLJZIpnUnPfzIL7v5zo9ChbIva0zFdOYLVUcO+gYXGCrL4ns9scGYJggM6je4kuVPt1jUx0ANVp
re1jp7N/FRgtnUQOOfBXvy1YXiKDXOBYm4QN3DteEKYwKGhbLSaHHiic7GQvT1tjCLQzFH8a2Z8b
hdBSitdLRn07wW9R5UqTOjC3/dgok1Xs+V/8QXFMrlc/rN5Z7VBGoFh3nHqpypxhsNMQkUQC63+b
HwvRZ1nnWok5lieO0PhpUUA+Jl7zb/m25BCeIYzgUS/uqmiK/L4AkzmZILH/NrfEqYALPacUJdmb
WXiqsau9QcbgFWRPjMqXg51ESxWJlXHiNCjwtZSc7a/miMdiwrgK95NtVuYrPmdETOcObBTzH2Ny
mgmu2NjNuPqwdbusLltHv6wgaZg5gHLgd3K+zdg60OROtR7w94lM1bgeSq2U5pnrlUoVbVIGAZpJ
yOpfPDW00Fdnc8XFVTJ3EAQK6Uk05kUM70RJRBnzatGqZLCdKJS5xMZbfxBeKnqLNiuVFP/Nhf6C
vE+QiWFxQpWsh4BME/eww+/MvuPa0m7rP+dKhEWrXc6ajnGiwdr1uf53XN45YNAtqugaVTWzSbvm
H5Lgd8Bc1xkvUbnkBFr/Ln2oz2Xz3rZw6VCfngfALs7K37I8Q3H7ttqKhDrVWpOnv1DeGJ1RXeFv
E2/fBnsZ3uxlHd/7K3R/zlFB7MJvig9uDEMAzX7SZ5huKyIrqZ1QRPN8Sqky5RVm8rj65rmDHV2I
k9i1RrJp8JBTOXd4WQvvHUduxnS+tCs5GIBnVoEWiTH99GU+XeaO5Sr61k6sfxaDDuyvsXrI0b85
OOL6OL9JI0S059Htww+UmAvGDMO1Jao3zZlY/hwLnA65aqr2SgqqKc6IHjzK0n1DKBmYFpSaiYiQ
80xNvZLUsA9EMxnUfAM32/GRnm5DqXVZUt5ZxwXy9wf4hjugj9eDQOt2EDX9xBHEvzu+IAo3SWIY
poYNT00IdQOR0DpGqrwL0IVgRYxRmjsKp340HCVBoigSugPSEMnRBXkHoi3mq1ONjel6wC9gqFFb
zlonMhPYMgpURTaW3OHrqEgCsUzlz445hNnYyXJoYdSGIS3TLAY7VjktZAG4speAuKeRpIt2eY43
W09S1aneBH1bhiI1lJpEW3lZ1hOU/8M8uKB7Zuho+sNrQNAlaqBbPDKwFR6lkcOk4evAmU9dmcW7
URHLCmPCUm75PNmdBUuUmQElfA8sbx6F9FYBPd/Bs7uztBjh/WOAcz+SGkYFLuE2om9YoyWPs5zO
D96Thyk7lzhX4Zfc8dAk9gXJsyIdB4oZj7Kb+dl78N0w3zcPl76tVoBB5zlmNwx2v/UvQ7U4aHgP
7Ylnp3HTUO8iAJl/vbS0M7Mep75oMdyrj76hBvSNScrmkdx+wwlLoaYiBki6VHXlSWpiMaPCtMzR
OgYDdaIw/WPL37af9ej7WNSlrI+bpmAOBe3CdsZxJ5XhoTFN91RGiQDgzs1wpO0Sw1n2Vpkx9llc
qAzptC+LCgO/UJ52jUy285qvpT1jNpk636ta4/cBg+J4mh+wVHY+aW9BQv8HYSxxOwpffjWoQfDM
mtxPPGpQjaQ9HlTJw+q5YQjM7v7yvYQq0BmXi4jU5HlVPMSh9c4Rnju3KvKUTtiS0QhB9vRr4KsG
z0ZWBiGdV9yp+hYr/Ad1VIwmOMtZoXkq+4qhmadmUCOleyLvWj1r0Ah4KCJ20CMbor1tS86fq6xp
diwhDAog4DQiVU8kU3Eka/oGzlEluVP7hsZ6BCx6SHGBDbb7Bl+9ns7OA20oBkDmEJFvVxN+SpFi
CMtvjOb3uUGBG3gGphQmYSZHN9viNNnikCPo8y+mZ8ZgTFhH//uZKhRZWOj0pZitMivW4fSWui3q
GER7YZID0yk2YDvCoWcRM/Whw7uXAgiDrhvuVefiAtVLJN9EyRO5Ot85fogCyxkhcUjiZ8lJfy/+
t6xtoHM4qAfS8jjMcn+M/NYVUzMpRVVC3HIa/YXMtFP98Sa6eaVoUAJkqfpT0qqqu9TaWhUOS+8r
scbjOs/ADcceU2kvx1vX9fNp4wbA+pTfUC/bEHLOy2XczXT61bvNIV/Eyt31k/szAdadhzrN2d3P
p2bnhUz98UG+PwJ/YjN2+NbJDykp1plVzcKjHW2QYwRVXxzHTb5IP0OTinLXPUbvyZfsuy54Rr/D
CY3OBqdYxpXgX1vkHZKvtbcdTLeygiRi1opAnPjtWjaCjL6RQSsYuCoc3XrV32+3z8L0WtG8VVff
tBU6Tc4V8dweD5i136LCVE/r7wYlBKBWTS3RIZzC+yGXn4wiJUNTtXqvPwvMI628qipnfyXJlBZk
e8ofV1Nldgeb14n7sdF6SUaJ7ML8/+5YnnTryLjbvsX065wXrG/f17ZMbmed9HneYGzy8XDEdYZy
gpU4fDCiNZaJaj9DhIzpVxiW9MmO6Sw5XeGwwOyDR05XJawOZsrefZYmAzNw6vauGLgVYO/pw/6d
p64qa3CdXlmL3tEdXaq1OQvx9/NR/GEhVucmNUobLM0hzRBIDyvOTE1nlG92/kttReOLAqLRRpPb
KzSaQGXvW3dPmUndYJzOHd3+7doBTt/2M1KgC3+iNizg79XcEYVn5qyvgieR5ko74KRCVJvGFAlF
tuI8SufjU+beIvXEW/UpvU+Qtb0FdHOhDRwHku3sMrwbr+S9xXUvPTgQ4pC0ngldRjn7ZLvayzs0
pHAi7vHgz0P8z/gkgDdzvstTBHEDhCeuZi/W+vN+Mh7aQwEeP/qcNjDvjgz+UL1hDzjcIw1AMpoo
Z0+7mQ8dqJLWtnwvDVbQUY7flnm9qaktUlt5mK+CDGMfvvDevrobzbg4Cby7i+R02Qt5MXpV78pD
a1u33ZDlFo8S9G8Yw52K1ZNBrBNJKj8re+nPBrRaEn/iTpvXPFbcALuKU7ImOpRtPquYwSorpcP+
n8702r3E6WkO6cpPyCLTwJn2QrI89wANSGH0eKSGJGwdVjvQxxq6nM1n9ICsv89wdoXluFj1X4hD
h5fGji6FzMPaBmXhlwuisYOzeQ09S9vamXAr4pExkpLxpddD4I/Xn0v69gdYU3FOeRoSLBEoTyVK
TAay+U6HB8ERc1oz+hVmVr7JT3MnXtYvit4dT3uSWjSmnx81yzoat2Bdgma9UBWL1jaNCRHnKRtW
V9+muGBdd4ieRBjeSRisidWJ//ha4T4ThSiR7WYKleW83B50LhST2AXBItSSxUCNV94hHCgyZUw+
Nl5/uQUSWUueXSpsLPY1lXHIHbkpZMSkuPh5xFBJKFIPfXbAiaqvQNZaDQ+wHESEzBHdjkp2Vflq
XAJOGzRWijv/tmrhrwPnOWHaI2i0fhl5xaZmg19SdU57rdUWGGMuRQrW2aL8o5PJw/9ppj5L4y4a
HPhlN3EZGWmxLTdrjQan53BvNam1jyEHtKIx3/TBzgOze777qVzyzk4mI4q/wgui2+gwwNcRcP++
Hz2YqfgfwTGazsYGE0HOXsvHIDr3yMtOtvn1uiO030R98aPUUcyQNCnGeZjCYN9BaJLxvDeoD/Vv
uMavUC8g7PusUE0GkP9zSk6+5fkzGTEk+UWKCFIb3jJRZjAkgOp5QLwRmOSP7wFqU5pUAdY3EYtu
E0dxIfejJvCb52CHhE8knrcaDq1sJa5ZU3sbkBsH9pSLbtZfAqqT1V4RDQqk/PZIUTk35gAFWYD+
zogtpuR1PRVf4luGhw+hJP49rP2sZ89a3kjsyflFeljFQWiTzuOfuHOudRr3vl0x8zD2ngWbJx0K
ZF/6R14aAydiia7ALePxCMfPZb8uaWMM1FOLeoP/D0dWseTXQlflAWbdetvp4+HHrUVWFlT3Fn19
oItXS+Vo6oxE0V+Kgz4yIhbbz0qWZFTYLOrW2knGC0ZIiBLcSbvxiivYqNp2dZ19romqkeBwSoCb
wz+y+yxDACa9VzRBVvuZiztMP9eh+ynNVqYdnYHO9pF4u148ENew2FUkrZ0zubAOeEDXfnwL/55s
aUWYIrZh/pIiDV9p1bfPGHmdIgmsHisnt6nxqSH+LN5eIcwwJJv15nljjW/U7XSMAcVJr8Dd+yp7
2F7cvqV9hdXt8Kw88sLwIqxsU3LEH0Nm6TosQLcR6+79/0LvK6VqGOjZvj7ZhoiFiEz/Ga8SOza6
z3mtb8OTnr2rLX1WIFmyjgozrpc3uZAwlgxXLL1rM3lYk1jI5ObI/ElMbtZyoSNhqInbp0RR6haR
r8qYQuhYIIJZWrmE2gzlz278XPSyNgQylZLfLi5JPjdgG8cMFljX0r1y9ElqP1e0+sFX+uT0e142
vrTIYWMy6PTCETh+cnu/+lCPkZH0GHo+ZlUnfkdETXgnCZHpSJ6x+Lu9tW40ILLpdALaRj64gXaD
ArDFebR07cRSWG5rt4o2rrTMs7e38kp8+iZfieBbYoZYy8H/oGUbvPgC0gfymtTAQiFa/JFasvmw
3OGFt75FQCGu5s5doVvfD0JxmX7bdVdV7xPU3gn+8e4zPs5tvoGDJZhe7IS/lSnxbYRgqs/HWquw
bFWrHbWoeXq9gCbF6L99sKkPVkqG5H9ZS0BI6VH+vIjd0wFgb3aKhpt09H5/9APjnx3wPC83t5OU
HvLyYU1v3fcrhezC6rzJCApgazxvIVhGPz73ODzY6/Zzjrt4bGB7kTZVmMEGslW1K9wC2xqF6xHm
Ud3bkQdmYTjON9Q/t8UqkzaV+8Dpr5aSVpWRAQw34iuwjlUnH3YEeVVTlbUUF7GLN2g8q/H1SchA
OA9GqebaUtFLuqYyvF8kxcrkHcCVpeS30jqBElJNmiNtMuUMC3zCMMMIn7KuS4vFdQrW/SAr0b3V
mba5uyE0kHjXGimh2v8puxB682KPdmqipu23ZerNXuDDk32G3S6cQQVpLLVzNoS1qxINywzaHacC
y0tfRPJcTVvZVBVunujTufZgMuce+MiLzlhYYf5pkuUJDXHt2HPVQa58Y3n6uMXdIaQ4y7OFJVKt
0EAyqiC/UMpQw93ZYdTZXeALDwUTpRy2plsovrEfJRI2neDd2Ou4v+Lkl7bdzpOMpEerPLq5nkcU
eIi0qQudxgClBpih6OMP1HFVr4mp7CykVQSwP/28K5jmigh56fdLVrLlfAGpDi1I6XaOO9KX2FYj
pz9SH4LxjD7yA0n2E+Xi1VbOJJNOw9/1mF82vhyhhdjmBYo7mBKVsVSL4ITez0rBBrx30Yne0PeP
PfdefGZPlFebYjojS7xKCy0eDY3cPRIDaPw2cxV7lkVtUdylWfmDJb0z69T+OIefq5XDJNpO98/3
K5dm3dVatWpd0H/GfEQ2ziZMWSRElJoynJ1JyhNukrZYjPzsLx88UjETGrDRgtFr4iHXtV9bQx8o
s429YzOXTm/+zgB54BveHQX5oUGo21jTDJA5Tu32F0Cm1wXbO2W27/MURPzSA1tn7GOxcgP+dY6K
LWfF7bWeleHlXzHLLycstNu5htBWRwzGKSOz4UNfHeuxYIKqMUhnqKTdZCMX1m89NK5rXw62yJSV
CD2Z+yuPmVHhPV3d/r2S3r95RJEC/jF64Qarlo5XvUAnRVvCkMnbnUSyOENLoxlChH/f8WGTMI4K
FIx4lYyxeHp5A7A2RLOWVWz+PinNs/kluN8eqlBQL31W5bG0RHRvIs01aESqu77W1lBaradXZHY9
iUw7kluIZDAR7QSp+aaYgWXKbHzMc7W4/5Poq6Tc8HdCEOPNdv160ejlv2MGs1RREZXbwabvxF+Y
qvfuVwUbCm9RRHhrmIz5HXC9Z/BnOgUwDmlUzO/sdRptc0dYb8I3oK5xsWafX4CLl7Wro8d0R0sf
eiSTbvKCBFe8d3Q7vC8/sFLiuOncJ/phvM+E32f8g0RG5Umvt5iz910D1w6Ed25Iq+MEavpexJTt
pEss3mZV+DARFDNjC1kQYTn89NCzKnpjUjaPw6N3c4Je1ESKoTg/oobXyHuwBRjWAybwju4B9eru
/c1gZVChvB0zDLFLANvdwplBGm+5YyVTMKMEF8gedIDTJl6171Qd/FgzJJ37ZaYMuvy6wuBah/6z
2Yvp9NFyHnWXU8INWxvypr6yAUQuPhMduYUJ5PdrW7z4vst4iNpMguqbu/0ojNycyu7V83riuWLL
QQ9JqcKHtw2vLh16LG2xAU5VHuDJzgGRrnGhPD6Ul9UQ8c751Mwm2giIQarqq48MKmzQBcdj21+n
Rz06XFZzocZ1SSnmjh7mvBY9QNcNZkApqsRkGSJfxj6BLqC/hwGdwLohu/fbjXIoSL1DgCJLI+F9
978I0w9lar7s8oDESxlxI3JEB1oWrRZFgebnTZVr5QncyTqO6RILXxRB5KHyaGI6YMb6xeSEJ69y
yLEsgOucxRhpn45w5klBPcRea8gsmVy/+2Um12XdTZSuw11Y4fVxRnG9hj1VcuAJmoyZxAob2fuH
WQWzhJ9bzf57YhKHLWls/yKAtcrIw8hc6uD9327KU8BSxl86Ir0p/lCz8qB6Ojc6nyiiY6pCgbYO
FZ+bI+Fq+tg+WhVT/JcWgWAt2c9dtNAJsYnn9QtXSI8HCGeFPk/FkT3KbvS00NpsFOEUnDHJZ4Vp
XnnsAnjxqBh3zFG1XVx2NqvjPe56fR80dvVSxU3EIFY66caypiajAA3PU7YnHZZSXiyod1Ag/q0q
/vDvDIclkcH9qQFhQgfCYhxkpWkK3JWqwpzX7db2F9FBcpYN95ekNjmK2UbFw1B2EsJ+PzqclApo
b+BAxuwizRUR2AOnQ8w4OYK+3cVYkAcikF7A1CEgh1Kg/VhEptqGyj148aQ+/vH6veGqbQuMs3NM
Gereqz8Zx8SkEfPbUSHp7AQYH5+B37HeC7j0lKVbSHTpj5s5y3DCgLWNEDYCYr1ORw07joe8rmLC
CpTPP+pLAith5v3PWTF/hHAFTAtsG+5bhCiTEZbg4E8DgkMq2GkbJJ8udyjpzuMzHe/uLE8NnBYi
zxjpJcbZ/0aB/xaDxXDYc2RgF+dx7Nr1FoyoPoBYDvBDG+od4fMh6xTMxBlrhDry0Btm3rCmVmPm
kidmn8LepdqiKWbLmLisycxdOol0s7LWA1i24/bflyl1JHplN1700kVkuJxXssJwr/QSUev5p6YB
K1y2drjOM0UOaLSG8e+lVN/I0PG2ovtAOeAqxiS+tGrHJ9x0I590OUjssEPZX/SB/PpfcNM6JZNl
E8lOxCL9T6HkG1cCffD9bSg/WuBkl1WjzkZ/ZTtrC5III8BnzuuSTqmQXMIAOQHNs32A3fU4QMQ6
zjxNOQNlkbAPZl2aR1MB29NlceYYimqPwd6LyqqOtcPDIFlNXGISX1qDSwiyEVwuG79iIrnmIUBq
x/b3kFFrL8LD2fhk/OfTXa11sz+JUyCvoVsDt18Y15Hknty6IkIFf/SjByO9T1+F8PDi6erxjBTy
z5wMByYo2BAD2ucTTeHEN625nApAmmZH5dbhFim9aKRFhwwVkkid27TE6lRCg2gbsGBv8LWQ7SLE
VqFDWppAhM+eupp0KimJSNxw/MFMmtLqaFqdGb5jy6H9R6eyt7ffm2zBnU8HFaTNvXoM+JaWTapI
mozCp223LO07BptQDHvU5EzzKfQK5Zbpiwqf/8Zfk4Yk7xAZb0XnpJxnh5Y+w4x8v4a5labgY60f
jlwKs/4rk+SdGrhq2nG4mEq714louLHMycfW08AfadtL4VKM7eDu7Sq+XE9I9W+84zRd5UywYpTw
iARSTUMTLAJb5MVc+vLElNUsmboDcz2QgY9KM2cUO2H6cKIBP1pUvbpg9N1liPPEg3ter4dUlTOF
3AMwgkS/iLrlsUedY0DYZ5xlxVkVUi0c5d5eEBCXLqO1gtAfDskPfAV/m8Zma3efG2M+ZfJ6gEM2
io89y2k+NU0Wmj+9fPOyBkKBrdqIaWkdNikv4C9/O8tQjz3B4Do2dS3SK16nFQPAEB9hDNEA/odq
X4FALw0fmP1MjLUqa5u3iysx7SPKSoxHcBQlt5q2cbJEV1UUvbHjE5417ZEuD0w0H0OuB0ogflNc
COwaNw9xPlHwnZZ9Y1Knkwg3wVR2P3U1vvaRfNcbWF3nMxf/69pXgKXQR4GkG8w3ESqjhtte9Cx5
Xv2MhjQCEvbDmGyQ96D0x+ZIOlmOstnOaMX28W+osqSTLTdyDoKg6QUgEMWeWtgfYGc434uCEjpi
OE9jOxqAmyL1VuKnUQEihLzAw2lGFa6gBfrGEtvyvTpSQ2i4O4oXoLdlc9QDi46KmMIEJmiE7CFV
v/WDxBtMxs1jG5ctqtQBdRWcN1tBBz4eVpB+YYukpbOCCmTHGyF0sEdyGNFd6INqi8r/yWCn0lrS
8cY+jzD6bz85IM8M1MHWbkWdRu4n9v1CrY1hkSTwsh6tLNRw+jjvb1kREUys6hU+La2DsM/aZso7
3QdvJt2sTULIQm6HP+9I56WkyHldJzfY/tmGvaC0KvhpvFJ2dvhi/wKw2Gv1a+T4NxG1QC7Cwa7x
vF3hYx2+ppJRyZOndkpaXfHmrBjGI+0bJsfsR6PpbzGSeqbluHWYlWq17FXXkca84JHwgEeqrF/O
FHqd835/hC2Uoeu+b2wKjyhdTwAz/MpxHIGH2QNIN1/w+2DyueIphdmWeyda7tkQb4LUV1kUfKgP
ZxnrPjhpxAbOCPfEkx/1PXqC1zutmSP34BRXjxp0rOBV+BN+BwdCYcQzduYu/MnA0bOcFzZk5ZFK
DDF7iSJbk60gMpmx68/zQpDpdybJPbXLG6vsThGn60JN3f7UXoPJFTvw3cIulacMYSxKTnyFziCL
4VOc4P9HBTlLqO2QbgXKH2dNIMCDOoo5306xp7qmPKitCU68lNiNUOPlpJ4smmyenas4UOFuU6V2
nWrBJeGJJjPJRPoKt6JX0MUrGy/Wgxc3fI9Qn1EfyhbZWf8LaIXpyI2lRgvTaITIrGStbMynhWgV
hKbD3EgN7gM2Hxtkod1PaTqmmhVcaTZ6zzkksSijT9pc32mv94sLJR+xVRAs+4AGT7FlldvIWaK2
E9Z5vW9nm0qgb2MLO8llzdLDSXOChGqx0I2TVGMa6P30iEfMs5AH4BLu/31fvRF7OFpzZyqsTzMM
K+deWH89w6Tg3mtGarjRSs4NkhKGOhcqWtgCWyemRUEWt4tTqk3KuGRpgY0cGGDC2Vrw2Prtl5Nk
pcoyuW4Ei8B0AePLSj1ZJVRtDWlPl8cYp3FRwSElR1FoK+z0tvzxf6pGKtsZPgAMTOO4Rf9eN2ZU
8lE72/WZ/B8Sny3DYdQBlJSxCaJb9sSFtJN0owzmb6ItFBd5IL+T+Dlfy9Jp6WDRbocbyp7jCGuP
QBzCdKgPZ1hoeoPHFEwRdfd7hGoPV/IGWeIwTd6HalfOYjDadd70Ow6q4Y5DWlI7Xlwp0/I1YvUt
czYkgv9p0jsjGespPzHCEX+OZ7JKI0bFIgm3MNMntDBsezS+YM1eNSRxFN7ZMo/Iz8irV/sJD/Qj
IAFSAK1KKYiAERPBKxtMbDUbY9g31vv69Dx41R+pln0jfF94pRxm5oXxfTQvxLDuzltWq2ddpWom
F6tGhbwtIVJQ6MXPMivu+e6Ym5r9gZqfd7v+dkRY8pc+c7L1ZUFJiuX48xF4bb9Bqmir7P6vN741
2r0SjVVgA+xZO/oOxt2ZIsz24ni4pJ9xFvALMUaLv17OqOWU1p7ZUFM68brVS2fXf5OKp4wiz17p
jqo4l/RZLAgTec6v0VBDX9kX5t6Q9WbuwRfzMyfNcPGZMWmDDCuWS5Fa4MO1lhQEqA0j1jCxpkBV
p2JhodZdzjtlVxQ1dVFONpvZxZ4vuc6nv4QSg60+8fbHT7x0jYOa8gh6j7BAOS9327vm8gPtLatl
UlPdOgqQtFpMLN3HTbHS5ShmCPX8UGSQ/6X2ZOiU+Uqjds6RBs8YjPvswIZ4a1Jfk1RI1BsixCeM
fg0WFytwVCCVZ6tzscKC907hbzULIC9Hca4hLjjzjB07ejk8HjQLHVTzsvKEYqTEGMNCZgWQNapE
iX45QBfBoBnNGC/jsz/iCXeGeaijJ20W1fknlHoYjv5VsGczHjCBnd0SDtwBMug4O/LYV0ECAVdz
QBG6Yl9p4U1Cjr3ZVZqMho7gZcVvCZTcmORmN04RUSwZujzcB6VPW/GetNHm/fcHYle2pgiXXdGo
rFW1VdlsoY2jjHfGnhgDSvczZRoytOlI9tj2P1iKVawPj784vvtQooGtq7Z32fn9GDyQ26KaoFO4
8cmIajoNQ0oLGeDwtKpxsfFiGWYDpF6dzjQtY/HVlY+eZzOgT1/h5ZGwid1/Uvf8CcjXbmNqWU2I
WxYTMy/xQ6L8mftFHoxHtInXhP4vvK1YcQM+Th+xFVhsNtXNgagjV4iLogSqMZD8jUQCmtKj1qzx
oPaJK0pVwhcY437w8JylfKQjX7XGu03RaR1P9XZHdc/1CqNfF7I3T2npm3P4Zw1D16DxgXquMbAo
/pilFf8jAp8sfpci0MBkR8LnjHaccXIckTvvqyofiS8Wdkk6p5dPOoxM/V69znI6Puq5fEr2GRn8
YVtIFdR5Y4C0kELJCl3FvBjqRELGdcmWQRI/OlfPrEFj4tjNQy16wOVIhEibEIOWwr67rqR4ZfzG
RAmqK5rkn5TrxKNdfz97YlhmJQQ9SRWrzzU0APuhBJJXLgjhxrr83HK6cHgWO04D/OpZvKVc3bGA
/qRKMt8pGqTkardWw0aITRxjT8zbVeEVCxwveZZxeB90SM1CuozXXWiOElhXuC2G0+1MiWvpUUu+
He2WaYymNA+YYcil+MQPKjWsP/ddDXmC2Tkznw2VgeZnQgUzqzkNUAHXmZevcjYWx+S4ianZs41Q
ESLv8iAwTbeZVBDy+hCeKlbr5JX+gAhKmK69M13jt2bCo7f3xwg5yHbdmdX+toslcrqgQJ/wixXL
HSfo9nc+xJrs0tshNKtZMkGwLIQBtGW/Qumca9j0YdPO3DnzR9dLgxWO0jYaKR3W83PBCM5oG4jn
YqPuw3aU4H1vxC9nZfNV71S2AEU0wFSGN2hDnnbPGUZ5f4rV1HrPtj0ESwM510r01Tk7aN/z1SRe
K8d2xpqEOiLL1h7ISa6RvUqH75MepA48OewDLsJ333lsCmA+QUPm3S+5AZodUkDWzAsS8GsMhf4v
XbzYDlfjz9Am83odd2sUR2Yb5a8njputI3RuCEnWC4oZkaDRNd1+ymOgAgRAecTeykD/hBuVOC8R
Foqq51rHwEXoS59/d0gJsmi8FHxVMQz0MtxNfHZlRJMVLvuW3rZ9UdwBcE3Vl/0kMngRtomzoRY3
TuU2K1l/T/p+5SbnDVSQxAiG76YgLiK0xxHzcDnfPcG12GL2UUSM3iPPgXkfJPZ2WLBhiaZS6oko
8RyA33McbhhLFBs4VXAR5tunplph7LVeLQXm2ryC1V70Di33BBwLie8GMWGQR241CJ/fAHkONaIp
Bknac2YOBEL2pF+GHaOlUv7LKjBw3uzGb1JpMoETizk4afY4AG6B+AIWrxPrqSPA5t3v7G9AtPO/
+Qd/dObtvmbT7vESCNLEQ/jsL0QOVn+e97ZYfv6Pgq/sdngfrPSYOLVsTSdCzDjtCyLrBjlt7Bk9
MSz7xbVcLJLKPciwHKiFpG9cggGxo2Z+uisejomWcLVh3iKPF4TKrXIHZ4RDjALlkM9uA6DvgESq
XZtkz9CquWYqgfA39w9bmv4Eg/9SPex+nsk2LgqOPKmOSB88xlRbULeqgVE0eAqIOBMQ07hP7l2K
yIERK9e6AeW5jpmJuoXOGOIXnp0IAI/xtYUSxJcUfqawQ/PS6vfs/hzmtTXvYAhBt/gxkPS1CiLb
f05Fv4crypqf7n82/DWKsOpmGMVd3aPSR0qMc25dt5vEplsXSYlrFUqBTYthhEDMPvX+McLCSMsK
RIHbxd59c5Fx0VBs5yekhpqVN72GyA7XaDRR+8/ZPLglE5YDXUfWz8DqivtHNCQuYrPGQbaOTDq5
+myz1l+tX5O5Obeocuuyq3owkkfbUS7M4wL5dg8h/RLyguLiP5MSE+fEPnjko5h7UVWlHzerUl2Y
d1RT2X458mUjLz3NksFCFsKW80rtsVyUNV66lF2+cqhzbXDmnyZM4SR4MEjpZmaJdoF5CuC2tDCL
UuN6NCE5GOgssIjhkPBvaI5p5rgvEdlhX35AAk7pTDP+PgeKGTLFWGLJm7TJyG0zvm4+bj0LThNB
s5niQhwMTZzgLmZy8YRHn4iYb0t8qcPIF82QX6nHDmGhINL0G6fTfL2QmqbPdYc6GJyTHE8Sn7RF
hEiO8OhKHG8hRb8hB17m7O/mhBOzyqD2rgvTKju+e3wdOCRqc1We+Jfc5I+GBnVZZmn2ZyOJsmUJ
97eiBC9FIckGBwzCnw6wBLAM0gKSrtDyxNdv2RpI2vmHWuM3j3NGQFsmyPsXVwgI0lcu5Q83MBXq
OhRU2y/QAWJl0EER/oOPpRkL87yyk/QvfsffCwaHKHu9odYVQRf/PvBtWb3/JmapYpCOZmONJU1H
LIKEtLls9wSLpRVMDvGyIwTa7W/o+tyGDeGShpy41xdOe0w2iMWhX+uwGK9d+WuLgRumVQcmbwtX
kgqoYn+5XC+kMGdkyLUFRbH58MtvWtDCU3UX9ENyqo12tG2ilC/aCqMsXKqcT7nAHGeOPJpp3/oe
TeOunwr7i5+zzcFlWlAHwaGi6mDs7JuNSdPgFc+1JtsqagK+DcmwNKWN/S9yDZFCMcPquTXORWlF
KEHvqmT/By4fjolSRZoV73VJiVZ3gwufPkpyfi6fNalnE8ip62nTJCYtoaDSoSxKXo6CUFf00wDV
cbdkTsckXzLB8qt2SwV3Hrm6bjM9Js8Infk7+v6myyJaPr0GieQ/ayjcnoWXTI3A2LmoLWdDIZu/
XsLHZul9x/oi56RDUzOyp+GKnEGyN6au6QeJ+4kPUjaaKQhiMdCscwVxjE867daGbbK6j7/oKOGk
KvXtvD6kxUlJDEnAEPKGNSZAsP8biRifCMgFK1DxyQsRWob0T2FfldPlTqRU15/ggWYi1f6cQKfn
uYjMOqTufszR6sTgmu/hY9m/lcpPti7XTbo2IRD6lm/KUyxGY9KlZ6U0nIpnPoIQzwoI+0HlmXtc
PKUvvsNkkOogl3h1QmD5p/VvxuGT2Gvl/NNKFwDB3lw4L8Pfx0jn39aBeibDNa3z7HglnFalj8dL
w2biYWEHxkFtFBk2V0/oqVrXuzXDAa5nm6263TOds8yWuJuqluqTRtYmC5z1GtJrDDa3RPlbw++x
eeusnNCVaVBZrSUxB85iX15DteirFLzMSNoYiZV1Sa7S6LvP2k+qTw91EcdP65jXp0Vj3hqcwItX
Rp+7BesyG8Ndj9ZPXrZWBgUh51PPTuBWOlGSbujqw6een1Wx3g+w2zMHx+HZ0Ki+300sX8Jg7EqU
i+B0pshnYeu/xU6Ae5bu7Aeh6OZE4AKC2GWiabw7xWA9UEuy1gzmpDxB97mEtpDbbIl9nefk24IR
DugdlQ8fdDr6nxSZzCaWxuyvhkX1v2VuGAc+OyKMPY8w7NBGDTeIygDn5oatnB6ULysxYDZmua0s
9gQ7dI+B5h4gduORWDe/B1DYfjrQ+2YQLskUQLT07nLLNr3SjC0KoEkYgHuK/V3dVd5jKWwVcz4P
p9fXEIGYfMu/Ny5h2yu/u8tSXtkwhvt1R1V0JwaMp72xXtO+h6T6xvk24u0VoM2dPRTtxQc92ZFV
gFZxZtw/tWejGipEL7LgwTxRxB4PK3+ELLjT3GN6+y/kb3Z2+o18vRHEhVQK/NG9tth7InAJQd7/
pDkVqbEcviNAcgpD7SlSjhCtIODDJd13dsrS0Qq9E745d1Ii3BsSyGFkrW2W46VMzqDZ7aCMxh5I
rX09ywEZsW2UUFFfC43awzwr+RJc1zruIYmdgwd5WrMR+oQIWnzneB+H6UyNUOfZMJudDA9U8EZc
G6OhjoENS1+or4DOe4EHsUD4Wk6FlVV8/cmv9x6BLblTsGKNF7OTkfB8WiLKuAASYmdAczRgH3Nm
EC1aye0gieACBp7Xp+ajEPRyPiPN5z+9UxOcNNVMl+D0N0dtiSWDTGgQPfEoPURvp72VEjrAErRQ
poRAPfiSQedgeJWQYIBqDs/y4y9XOcsSz7LAdego4Rv4x57pWS3zs/r5wQAO2PY7L1aoxH8J3N9c
sJWr6dKWifFWuvB6AQ8U0UGYwEPfmjUVVJSkCeVel6EVslF6OTHaH5GiPFnvp1xs8DSZslIcqYxU
MFi1lqJF9iVtc5ce+HbpCRQK/wdHOXUgLKram0nnE1sqbraiL3J/tG20TGFhUtqDmf7mzKvAPJsH
VmR9UCsiwPvTkvGKxY18IdhGX9DAGnYi4dmd27jZW71Ue30twG4WpBchwUeutuoE+F7z/BHJWZVn
vIs4K3cz9kJ+IF5Li9V61wFlYOOFiksZuWiPdLzwzfRihFqYHf04cSiFiiEawEAvuJApI0U4XxRK
30hXkURGqmZrsZtQD1rf7IW/cU4DK555oHnyft42KaLPm7Ofpyx8I7OPCmGDWmchkUePD3k6xX1w
i6PfC4m7ECPz780K5eNKAjeZyk7EtQe7QZEowrW6nPoUiueR+P9lHk0502YNwC9guUDjZysDYJwA
6j8dl9x+nw9rVZeApku8j1X7+1/r1GitNdOkqbh2wLrSU4pm/6BtwnvwIQiFSg0Zc0qf8EZ2x2mK
2zI9OhZEi5L5JSPmxDNwm7YJpk72NV3+IkUtFmOkzwQrcQ4rC9kMfDcTFkxqcwGnZ2Opa1jxmZ4h
xmLqv4wDVljw4inB0gwx8FC5217eqnBxxG1V8tpK83rRslZ3RI/vBAoTsOLQCplg4CE113n1sCzj
5/ay19loofn5ZyBl74Z3a1+4txzyUcBLlKTfp1+v0B/0vqwfWIEmYd1fdTCZQypT6rsD+QUFsUGb
1aMa8o2KgGxx45tftAmnfzCuCIiaeulz2lA+wPbv0oah0j3h0sEZqxDaAMrDTEqiUsFJAqWpvo9C
dytzmLraVeCJwZCaM4oQIue6SLrYVlLvVXvXCn+LhX1PQkNMWn3dVY5oX2sCNx/mgu7MRiXBppT4
kLHvznPwG6CXYk8ueHqjesdoDElMsa4z26Fximc5rOoKLO6R36tMb3vOZwjFyffyTWR2g5YQ7bB6
mAl9imOM96l0mNjd3Upxw08j2iBKUikyf6RP0LDDCOOGTT+bDCEnd/VQN1da93A+foYfKU9qZZ1H
1bHhTIic+PoP8G81jkqxAOn3nSuyXlWsgAmNxg1QRTJW8F75jrtxFLwzH+lINFm93oLZCw1zi2Ri
LtZl8yr1FqgDrl7mKfLwKGyW30e6CQzYkaH9RYmMPcwiSCB+/wsQEVBGHy2eWMS12Rr9wS+qVoad
m/Qqz0mreXhukP7NeA38A4WZWqzedeCUJvbbSmySrwGOTrEVE+NllyKrSaXe0taDblhtQjGUGXSN
N24D302lPOePm4g2W/pdWY/ib9pfBggcY6vK5GnJ9V6cW14RcAIv2Ex8Rt1Us+4dBUGphsbqYQ6w
v+0zogcK8NSuRTY6/QM3dzTaMHcpbRKQ7HrjW2dzMwkj+csUBF1E+iDI8uauZDz3+sTXMnaT4/Q6
r5Q00ru5RtiHO5fbATXDsJMoil3iF5N9NWEyXA22PpgPO/sqeJwvXka+5YYynhu9UM7EbEcWpyXq
nV6P+AEa0xTKaMPU8ujkas1KXE3Talp9xWilMqUD60ZCh3RBKy2xHuFevsbqfwr/aLzh237GGgwH
blaEpWlowYEHs94nNqLpV9/sTGKSRtvC3fy+Nr4VBo+Ofv7GRV9pBPTlokejE5uDQnW4EsdhH5oh
iscwzc5WuhlEzlj2utN6N78xDLQcco7otYHr7qpk3kN5j0Vea8aI7YfvQWPSwC8tCBG8tj2MvIYd
jq++OLh75rXdw5u/7CzGyOqQ0FVqeaqajeNS/AxkTM39dJ0CUeTklZr4gG3Z4/Yo88sFZ6IFBFbf
Yu97tAnJDRI2aasVyn7HehE4QJ0ENugeJ3IgMj9LIanjVmVZn6PJVBND5ZR08XfvYAnNigNsq90Z
7mMvWfwQxiNmMCxIYHl9M/rXBFnlVB+RkEOwJfWdsKSo4ObhN6TTgxFinl58fPZ41/pUM7tmgxw4
i+L5ZQTuHeVnIbCDAzdxwZ+o/k1aKSeg8bHqjcPRONHh4aSRb3ti2dBrUlifmv1s92EI0WOOvlSb
tsSBw6wyv+Jf6l4bJYh5fjKptwgqrq4CWSg1S7ka4elh+dVJYDWQQKd57C0/o5ezyVKP9KXTbSdR
pIledwMpnn+hCKPlPiN0vt8R8wvGJmnt7tOh21cZwHidFcTnaE/8MNRi8TVevtdxZ6O7AW/l0LsW
qS7baXLvUHfhal2VaAFFr8VJtzY2EdPflAg1nZ6Ndk2RGaXITYH2IbSkHBYCEr7mAUE4wXODu/Tz
fmTLd2+AclMzbyVsFIqA1vPHMhdj+vP+DBi+5njXp7+uubZppVzc3hskySOSEclPgFrPRDI9YBiA
8+sIPu7R+KZwSpDaH452hM3CG0vVG3ROVyOekoevZjqGBTZku3rGK/o1zmnOJsXbN1ACkxwVEVOT
dcld4UbACQPeacgmUDwzrhmgeb0qebmp1bzMVEg+zYWlaSInH/o0kifup35NmiEnDJekzVtUuyH2
ER38nL4r+zoR2zsE0KpKjQtDnwdBTXU+yh9MTcgDjGW85kyktOPI3saUYq8TdqZztjG5YyPDN2+m
xpyZ2ZEkArOPuOXMcYTSn/RUq9Z4hdhcxCvrhwK4EcYNu7f3+dWUivGC40lERfMpl1SqP9DFBFXx
Zn27AAXi/LAKTusM8r5lW5HXMX2yc4ydqOC8MBvo4KlykNwXtnrO07vYNj75VQcDsdl11eMUCwRi
ViTCcyp2aSkneI4sWkRqmNcj0JZuG9M5YCcoRGLqEE8GszTkmL2C0JwlwY0yFB+sRHz00AP8q10b
iInpf78gGK6M1oda9Diug/NsWBBr2+HnErQ1Y3OQTCtENDBFoWOMq8CkOTg2Q4XagIbtKy7P7N9i
wnQQpAFCP5abWUtct4+P7y+b2B6tYxPjknVedGEcN3NTiFKGhCLBj1hJtaINpfTOCAt9I2g80V3Q
FX+qIIC7LWYsXrEHMmuq3LAS+LcP79OJ6YEKg8dF4MRg+5fDQEv5kNf/YEEHb8ijaiB8SGOgmkYx
ld6FqlydXRW8FpEIOEvSMMkC6t3OUMfrnqiIvaGQaq7AgJAThXDc2E/FcRI6sFHxPPcZ4O+1tYpE
rcr+rgypuVlOLpNt2kncY/l/d+TEU6bVAk8WC09bEbB3czh7IxAXw993ey4W8asOq9xOvdyJ7Pxm
hDrDlMiuK5BTN0U0lzeUWitX4O4J8mQKz6YBfihCs3W2V8hh5qlThkcK19b2jWp/m5uxZNxj7NqG
YiWcy+K49qZYnsUEEervAGa5+r+zUllYXPBWPLF3cu+XRIEocCz7QzTV3pzF1CDLtaBDC9jwr95f
EUr6JGUU380fLxnAvXXoOrWQJ0y+OHL2Ttc4l/LrBkTthq2nbo/p7JmnjbJZYqHfu5mcNyn2Nr1Q
hue8kUMn537FDR2SmLNp8mMPlVD25jph6Z1uWGUuS2qwU8dLGKLfykKQZ5gwfDFaHB8FS/ZfaxJ6
T3ueHjYDclOy9/BT124bTj2tOJXmmTzDszRHwujeEItSjYPM9ENTMqNNIP5vB/wntHlJE//zQ0Xo
3X2HvNQj4LLjc8JXFm2DBt8Nl9X3jPho8f2Aiv5nYYyPDu66nZN05IpJcje5xUY+KJ6vkqZdTOFP
37AZwuHBOcOsQS6ALMWewRKf7sXnW0EvlDtpTnRbrtVa77VIgvbWqzoG14gtXC+XCPpf9W/k8sgh
NdoJbAcPjH8NIWm1u4VAgoSHra9yxpBCJH9Y20gTODRSE0Hhz1N1W7aSECoLlOswzmDxSfMDntOj
QsihEjCiznVvTq3akF7wJ+2ERcxjwRdJy9virwnsHhnrmjk/vQyeVoGUkwtVItyulg4nxLI6kV8j
+AW7gcY7HzlcyrPy4D7kznfJE6ndU0+lg5rtiWprunNw1zXnCkjhPG2i5JzC2kh2xvReFT+iuJfN
Cm9IcXdECFvIg9WU8ppzQE8pSGllUBycJm7YVVKfe/rCPDHLip+8sTcVvVq6M9xINzN2LeUqA1H+
ZISCTDlDibFVCBSsjWrFeRpCp/ZJoheCNABruPU1v2kJH6ZIcfWpeY4opVeoDvkogchdzFPlu/WK
jSHzRCt8ucaP8tj/FLVP79J4XSVHr+zjk9APyMkexGhYDTkqkbJ/m+uY2FelxNAibyugphk7VDWu
sXvoztF19gYw3OAOIjtp0bFTAuesGAez2EgA+c6dbTL+pbE3wkW4UASrqoXQfN7b82LnnOeEH2Db
yBTSYC6TEcP4KaINRTBAUWv3IwcrdCln2GwvIyBwNtU5WkdS1tS+Rl6dcDzIGq19B65KzAdxt03x
qj0zgXst8g3dtI6NXltus2EMArbuqBMzmH14lBD1mwJ0K7LR4clQcAnJ5u37/8dImU5OM079YRDn
bBF+l19PWaZ+wawdFCdxJKaYQxV5TCC9BEqH1CamSQlszcz4xq6/qnY+smotT+grxUpiVHMHITKU
z2xqcLW2UZ12/ZyIhhhVyMwT1Zq7QgMj7uBzdHlN6ILXTv3d4m36IvbJemrne2Ys66JsuXFjjSkg
3hSOT2sSSxHkTDz8OBObbKlrixOSfDAzRqpiLxjra1K79l53VdvTueJcAnzxu5uOHCpzokxNArlS
STpcwb6GMsSpa1mnWkiAqZ4DvnDEm7rMCIzpzbU7t8QW5elVinIhc0krFahyf4iNK5foTRIbnZOa
erNRLnydpQ3q6x9DsXatbCG1AZlilGVthgzLxXXmNi4qiyM9AdFxC7JJkmqcvjHXc6Ki2Lbi7Hgs
eB7mnRu4JwXdrN1LcLx/hxEeRH8FpQr2iIMz7ytDVO5eQfeHSiRjDr99UfAF/2SixlSr7CbGJGZV
caJnIaUhSiO3Bg5BFjubB6tAWpWHHi98Bilfd7nZgAMq1EFN5iw6qguG+590nlHwyx5IezTVlYs7
LTo0neDCETeSJrG9oskWKPoxb2Cs6kmIodS65Rv9H+gR0wCKZ5UPOq3YRgh8QD3mDvSKBi2xU/gX
5ALCe/udlchCa3XKqcOWtV4WVLqJnKLV6ZVw+V0bcYahJ1EtgfftpOSUuT5F1MT4OWM9L5abnP+9
DWLLzJZsyHtKM+L1mKAv49tYNfaYROsMbYJjwZHLuOvk/FFQ8yClwo1l3jtBZpsjxCsXHk2zyg4Q
QWeG4PQmZdC2GkRr4GVToVDTu0kEUgSM5ERE0Py9KtYp0y6cVVPf6sh+l/0ofwTp5+tG63F2f2dH
qjUsytEmqbolIbU/AMU7KulTYKDYzp+0PJkvOREl+OO4po+7cQ9R5ldiq4tgo6YRDaBiECSHOCpU
6HI9MoeuQE7cdgNjVo8naTPKdfdlQL2LliO+l4lWlAvpJwuGXdn+AO/Y80mHLuDbEGxDM7Ug6gEu
5JtH5UPlnpPsfv8lzsBVUgXUPouCSA2UYERqLC8i5AMXQHGoqCHdAXXSAXPWEHAHZ5H2rof/ilEg
v5uGCny5vOiKBPcPZTPRyQSTwisNpx+7lF39GorZ1x3w49dL7IVptiKqMAsAlwlGHM2UyhdNZW55
ZCxaV6EUv/b6erKoui3O3uVdUefNLB8AGsIJdex9BlNObN2HTTL4cHA4sGGUdn+r9DJPJ1HlOPAW
XtgxeZiz99YSaDzOiRZXDyYtnanbwn0t+nFubx1Z/i9a6HwxaNzf1ZP+IDby6bLkU0LuwqRAqmUn
GJelCd/JYHfhaL0FS2psFnHhG+N/69LgkXmmu4zIexDzlYOEApAdp+vdFfm+0DyPY/4x82e8d2E6
4vchV6UcSDzP8UwBORKcNDg57mma0pFQh8LfwzmrB/uL+FTWaoBt1sBoWGR63fI5d28kaj0qo3w2
BwmTc78wcXSRos2piqk+3v0f/fUBQfT+zKeh7nluGRVCoaHRxwJwCSHbIJehAluIR7UZrMODVe8b
mturW7UJN2XGA5x/w6HFetRz2uPAsyFzxp6BPvgXTvc8dSJJfmXtLP1WMqJRnWHwosyQAtAABGQX
QNHUBtQNu1WICis1tViIg48exnMLMIWXO+GFt5GpICSNTRGkuRszFrp/tArRYQpF1h8pQVTugT5+
TcMvsE1ZctJvUZCAmDKHrW9MpDfVqjDGDdFs3QhQ4+hCq1o2l+E3L8ojGRuIHc0cWFAGpTMnmYKz
l2oLhTZ94/itVUbsHznsmEZmeklpnTAqi1nFuWYlkSmMf8523/2xtMOhfmQpBlZ0AJRddfWrcQW0
HvdjYecLEcDEtWjqDBmTAyPDeWdGhNSd6gQT2a5gLpf5zwHaWdKBILpuXKfu3sHDqXkzx42lm5fc
8+I+dZbaEhf1l4cEZwyqhdyYHbLFGb4Fo3gxnA8+IE8LEIkmmEIbTb+eR06RUL+F7KY41bWo1eBc
GvGIFmxk3nczyyfiYdHuW/hCt7cbuQYn2704VHgmokyZz6NLWzs5efeBmIzahwljt7rmbgelq8Q4
XUWg08xhoEmJkTZuWCQRR0nCZzxu/3oS2hWbm0ULRFQPcbkl5zCSH0WZvGlerhKMMMwJ/rUVbGNe
kj1mWsLaU5hz3fgtDFTbJlOxAJDpWr5RUpk2gXKEp6YRm7TLX/0Xzmmc5qPDT8yB7NxBTQVMk46B
YW2DCRVsxy0hIXB+TjWBaIMseOcgFqSn922ji7T4dsfeK4pD4IiKC7RjqNPADxJ6eZfohWcQd8lJ
owVgytsDpPVFO0Q1gHnRoLrS5GBZj6qJefHvxE2pZwjCny043zL+/fufqUDaUFGsgcJqZbqTi71U
svH5c8qctK0AnTvUHPJRRbunC9OdIvMKPIOS8p7xEysMAImxT0hvMDgadxn3XmAKgu14NwG9rbVZ
u4c7T/AroWUSARqt6BiBmgTui97fiFhRmf+QptxjAFApXCgTgSsDgawuRbq6eYwBMjYcq+T0U5BX
fS9ExeXFuKtfzxZ+Zzr1cF4OnxKuMJCdoRuUGv7+FM2fiA5aOEDL/aYIW7DfxtQCeiePISprnUJX
+QtYS+rpP8KBH/hFEKgycsIZvPFq/M+IMsP9bAZoi3nvnqeZGsgm1QTbDQIgZvZCNyiMRTo4K43t
6LgiVovhrvPQeyZIrRXbsxfBialiNaDhUUNw8wINsmz3XtCb0RmDbqteDeNqTBWGbN81k/TUWnFr
5LpscXrqTYRnOXg8vgJz/STXjDaRDCfLXdSxENbRT3Bf2TkQLPDYc5WpZWsQ5bMjIJqT47NbNdcQ
JGYkR2TYWG6GXQzmUf+Bd2Fs/++/9imTdqvPv+dKsCzub7Lwqcw7Nfh2gmYdIUUgpPqCpxzYHNs7
bqkPeCx4MG0FF8C2ls3kCnbnUaS045xiekyBLOKNbjrdz/THMuOEzyATUlKboHLjAqLf8x4OskKw
GG6sxFrjmfJ8oldaohVDVEF5aVwfmC+hDI+F9aVJg4Oa0oSsUwtaW2JK6sa+9q6HcStCX0OUAsEM
uP+ZPEfv7lOHtOvjwbMSwDgF4I4CxTxlpMwpupE1ebxvogFzod8E2oG4NYh9qEu6yKhBTEf4ZJQ0
EpecgY6ZZGKL7YcbLzq4QxBJ47NZX85ooo+g/wWdzRIIu/fQNxoFFqkQtiAljpheXGsSQolK+Xpa
LP3dd+M2lkiHVC1hXC+S+hjPNjbZ4MbtnA4Tlh60D6xDe5d0Kp4GkxZaAn2qaw5Un5jco/eFVXXB
6UfW0UDYuzoFsYuo/2U0u0FnHRHGAHEok7B/WvdAHgrHeuCqemiN6ILjLhNX7mDbanJWG9yj9EUS
gNxBO7r/Q3ebwdIqJ+TyQdb1JS0a6u0bYIhfAp7RxxQ+hAD23mNO0CFxYUR3OsKctwS8HIVzf/Xi
OR9Iv3JoZYcT20RKfDQhMDvC6q6UozdcDHzxUAns09lAGpkrZuCWaXkqiyEKrH/769kX+vCIDOC7
RUPansWMZwzhYFwsNV7MXtXrqMo8JupmbzyNd21PL0mqOmHijYfJv+gbcUx+jl5B+qihSyNqrTFO
HRgZqhEwLvBn3nrcnvIRY9VgGUieHVuCz880tyqr/V2Iesr7kL8YsMqt/3oN1lsJAIjLqigJIdla
jvEnCfG4Ov+nb30nP747KAvEPChc042ZHXOaD+1OreEDPWfixbcrLlt6Za3048n0iMJpv+Rk92cE
zN6eNfzXpsy1RX7HmZRikUYj8pXwofTeDz6TxmH5hPVIf/iG2r+GQXuL42tvNoItbxr1tAbwERHi
oVhhY3piC21bPxvx5ZkVk5XYvo3GdEt+tXTR1MIFnmMztiZPDvXv6N2cr/woh3YaHzv0a0cj/98u
mv6T1AsLcmccqBEmqHfcSwQn73A8gmtOK9GXUDG8lOqx/HJN6vEXZHSwshZFM3qQO0UKCHzRoJmW
+KnBDw6LZEKqqd3Wykz+a6AuaSIRxjVdffyX3A9r4FetYTMi4rlq5QQ51TM2mlx0o/k8nkLuJOP8
iR8DzUUVNYjI4QrFCoWdMG/Wm8vmwDvBrv6cVpz08v+x3JSmIn3ZtL791p/7hXru0QcPQ4Zz+ibp
B0Y3tXt3ANm+Nzn2IWo6GILu6SEXIpmoyOW9ZuYaALVE4Op//A03jiO40PCgR3QSCWyu+txwbFkG
bnpQ6S8fLgJj1+ajRZwblhGnF9MQzNcD6HwWNsQM6y6EZ3iQ/fxFvK8mjjacFPEB4Ut5UtnceKG2
EUOu9wQKvyCrxARkCsdImlJzpXhxOwPhRaq3FddjvYBoMu/UeJb3EggdnM1ZTcKLD5VCQhSavq6C
0Z4R10o3OgUGpGdb95WRace2T874K3FH0WHXAlIZ0JCDLkJm+X29/WtkHruPO0dkB3oF1cNjq3ZZ
crhY3ONRBKHCwHZWVPtQz+CPfkzReFtt5R6A4TAkjJAEKgHcgA7G+tAP012sZcWv//cns8VZc6c8
YWkKAJYwgVlloCEj7yIYzwLpbDFMh82+RGtJnO2btpZUVkPdfOlqzpdtFNWBCzpfFbNDjY5OyMpX
mvNnG44EWSdqKxxk2yFGifUtCbHYXsrWe9bpUrRMJjAxejJHkss9nnuuLB3JL23/9eCW7JT2+N6r
XlVGCn3O90Eo4LfUckZNDPYRp07UCeWtwQ7C8O5qiY6oxPfbLtns2O7inaJFdgojiFXv5istjECi
SFNMftuDb2jwKtX8d4Mjlv1/b3HynH5sDnrO7KdenGdwab8zD4fuQwAobcC8OxYdgl4foPkGlY6f
2d53boN9rIO8ycSGH9+VBIzOczemD6Q3uW3W3qPHRNSP2QGxLb8n9gd3hrFfW2eUqm7L/R8Nd0oI
y0KLlE8OAEsdNliUFRRJU7fFEn83I54jdxtfVKn7P0pxwfd4xJrWHgL7E+xx9PVkUvVEPdMCoIeC
xY8kw99vog5ktvq8Nc6kAQWmBbKwMzLBYJPpZx1KhwgAgV8MKnm/iPhrx5yhIOTYmlJtrecsdjaL
h/XMxEohSMMpMQBFoYPxCXVnIljisH6nKVMa4z5vjaafceJ7K19HZY7LoRJQxL7m63jjIdRzkco7
PqavvzlLTHSGlTizFzN3uOS4rUNaBzpcrwhhOLNh33rJGGADIMDzQbdldwnrLV349bgdhr599muZ
3MatvNt2CnpBJNbMG6jcQxDdhZBE3GcqqBVhnaIBvcn47hUUQU6g+dx3jBTgbu7Oy/PfHvj6GJRa
Xr2SgTQLiBD0LwVNVgx1BJ3xTJnsFkgXMeI8PkdGDHch8fUktwoZ34YHBpeoqwTYOmwNeBZMzeo6
eO6zfp/PFpx+NzzCQjtl2Q5d8I4cdy3tRPnwGvvdpeJI/RREu1KowywRNOJH1+/J5neDj5MxUq7J
BxvSvPxtZaRgqN8cDRiwKaIWaUuCtNmYoiV2QKPQeXswHLT1z/5z8gB2ud7iprlFQ6IouF6LS58w
/88C0KI7hIdqdF+lfQ8tm+JD/MoHJ7D840AByuWqNEYBOHMvOAVQy+1y9QHTA5DY+lsp7xD1TFEx
qfgzPBEfySn35M+jKd4w2SW9+rINFUUskp1tqRFSEhRg+LnXP9RJ8m7MeKLjWexRm2069SfsQuM0
KulbYQhq0AHfHG9FQ3xLlKNCzfvkVXGHtfH2spmXfKmy71+zTSF3DXbPgVew0hxNc54bXNvLGrhw
HxbKcFX2v+z8PBkFMqvUhYlrLVSUBB6FjsmoIKcXpcwowC7dXZ0Qw9SmLBhFvp3QOL2A/2ZrZL0k
jWj83prT+GY7Kuce0TpzrYbq3zABDXbqcD9786l77sxFPoBZJdKT2ry0fnVMilUE7YDDlspgw8eq
/wHuMcp+AXrLPX8EGiUUdt2ofmpqH4oyAFeNMEc12prph5oQVZMNny5eoNUaYZt26eG3j+ZdqypD
3dkgsa29W1slu2NLE4+IzKiXmQWbE4Iy4ehbaCleaV5bYqF2OYubPxWWMqYGgxfJ+aGD1h1H5wg+
f56A6i6VUKfl7bKALi4OWTnaayz+bgu2R5vEbZrsEP8vBCZU42FMe9Lde90Y4GpGEalb+B9an+J6
e0p5jvJw8IWvVR985kzUW2mA3zXFGSlVnov8dkpDQ7GfTr/dJeOk2btnIIK42ZZz/zQWvNIUwZbF
Do9zqspZirMfCyN6WwBTaz/gW3UAd9hatvKtl6UeutjRD5ncsbSb6G4oktfts1/OiaM6XabBrF51
5F2sd2H0q9DitBT3jvhqa+99gw4gZbGNH+wLz34E2otjJ48lw4Z9cQ2YdCNmHsUg2F0aD2Z0wFLy
uJ8MY5Hptxky/MEVCMqwfKhs/oKkktWJbxJUKm+/eR+Ou/dir8ve8eHLuaPaslZCU7SxEDudk1IO
DHhClKI11Kgds8C61iikjxDCYnYEElrYL6VRr8blC3+drIF9Px4zLZnpIjXgTiDlooXyIHvNU9bl
e6Vti6KsLwxjTWxz84p7s+AG2hL5VL3ChXTZYTXVHcbeNSlGi0UGmrfPpNdqkodFypSxEB43641S
9J4FplSKY1PWfYVgRnpMlYGKwwNWIVvmE6z7A/KStZAfTglEbqoRMCwJw2DQq8UTEg47PAXlKE+h
oW4sODaRZl2OBFfNaBjW9TLOT3dMH4GRMMQAa9wUbUj5eMSLShyqUieZXZd95hNrK/1QyE7dsU1a
XEFC3r3NznDjG38wliUsAICsNv+Jb8Hzb9WHnCK7oJ8szO/4L4WZfZk66cYBbiM4vOI6Z4irt/1O
bU4aVHppJ+dKctqy/DcujAKWUMApQ1GCZxCK6vE5idmoVeYQANsh+bgJmTipytc8nWnUJ7WrDYc1
+XlJHYzs7GYJClrqt4noayUCw5xj2J4A7zdierQ9anJbWBFmJpDFtXGJhZbLLI6tayOnwKxmY80b
Y5yyWqc5R7VtwkUeNrT1kR5qJ1sRyL0uLQmObN+n16XREva/c9sjeIoqe3YOebB3yJEAIyB6sukD
pMlE1NCeP+bOOMxZgWn3eGYrtYmA60DsXakJuQmJo/Vs2nN3YcN2l2Y5bBMN4DQqypNIwrGleiSd
THY5LFMVk92vjot2z9110zeULqr3OjWW6UiqnNNr0I0NEAnx9mSorMYeZrzEZN7+L+BBkA5tDdJY
qiRBaS//g/rDGpwpgmU49YS/kpNOICDVS57ZjbVzsLdiZccoSOYTnGk0ZTtGObMm689v9jUgHUo0
5Fd2RhZTtLSqZb4GK1DrE7rgUAwsDA5Ul0pvvheqW5TZ7NboaD0iP6jV2tBq4Qp3b7pKE/AkdvwJ
eeGqC58pMQw4GUvXwgR6yRJQ6G24v4IqYoxBgMOzBb4Uvd/XJxYgMhz5WCFn3HzH4MuvzbNEteHx
IWmOuC2ZLtY64ftofI415xtiKd4LjEAaQAlRSMB/UMyZgM71LOmPV+OPKmRWhfDgW7582YdOzDHa
qw6a+PmTRKclXkVS3qe/k55anPfAmr/3EM4XKpxGLO7Yulm8ZEkTDW1TwyMY9V0GNhqizKi9rNZv
xC5tVH/K1ICbcsVznGUrDIylaW+7yBvc1qLMVEfLMFjmciAAjK80+p0MCbNzE5r87jsbxGy/xbDS
qzZJjLd68qpoG01eyQtNm5rlQWA5lw94h6cqeN8LlqM9VngFJA5wW1asObzxoW61vZ9Kl0eNfIRh
1Nv4VE5ULVh6QAYuJwQw74BfiBBB+xxZoyT+u8OyJol3rdX9adddXpS2Z7ARd3m0RG/JwfeKLLkM
fwQ499q4GZQlxSg3e8x1kTcAQnHurWX8FxR6duTl/grInOPVCZc/qCE55u6Y7HcNgCj73eiHcP9W
MhieFWx4/6LWMqY+rgBJD4EQ95ctNN+HdgTIsF2sr7kKSsjHWlfW18ug7azI0UDEbqwWts5JpTJT
dtelHL63jX2R33XL0lnetEpkHvyyvfVAPz0SJxbtwjOyuhVBDOxO5Dh3ay+Xj5wiY2+YzX+wqgpf
dbigo4yC++cXlJ2e7aLe9Z5oSkvfipuFsthjgqakhhTlwJGEEyGlML2hJIKxjuZgEx85nfH0TsPi
pLCHe7/CiIKokynJCyz7DWa8qM+/v57OmfmF9Zufkm7WAAR6dtsrWXWk1Ogil6x63zYxVy1a+fQo
XFJtG1nKOAV3rcurJiratS4PjMvg5lp6lx9ILsswbc3mX5IgOLt7MrcjYavCLgm41vUJxMM2sePS
7or2GXl2KcqKc6OXgVqy+W5JNjKgmLGd8P7e4I0OGimujm2ScvKa67OY0jchYnYYdyLeaS2mLFFE
F3xsRvK9+r1xMQ6JKNOl9swDVP2vIbZ646XrOnYVSLqWygSJNH66Qm+vLdTdkB7WvmbHIYhhpdlB
9iUZR2VhpT8DzhHTUk0G4cH+TVPgQyNY/VtjG3sVUhbyAheembNh5EX600WC26JRHZ8r+tk8lbQI
PuDDfd1rMzKIUvbaX0DG7UHiWnSsT4azjuvwCG4Wie3fOmGurCJfPmairJHXgIHfzoFwiQzpd5O0
GV0xxGMENM0l/MvZ3LtFR4/hIwiSHn21He7Og4yOOIz+1cTLqEfS7BOECzAno20pPSdi8YfCB7l/
Emc+T3jpedej2hF9v+em+39JpTr5zA34M3KTw38LLDOwqExm/nJZPJ2wT6xVpAFSBF2FagBkFzaK
9DNjHE1tJtAsTHfyIX/C0gDzjZxCJuoBoc5EsPikmIqJHnpgpfl5pewS1BjnhqTghWLrzn/R0rBK
NQvA+lLFucqjI3VhrLenJuKw355s0bDR3S1HLbKAB1gB8vRMizNV+17ftmIB+pf2rMJJFLkRGZpE
OkplyW2TdAbgVLt1Vv/kFeEdavPbX1GAkOPCD8e+P5okoKiVq7QgqhlD2s6hxacIbTJCbQuWVYpU
TwDvNZr9V+4s+uzQKTNXw5i0mApI0b0TjpbG4XO3o85FyjeoxlP1amTXU2BDXa7+nI/UX5jrKuHd
BxV9ngYU0APLN/F2lDxE49+Eo99mRxBqmLnM0vkwMr43V/7/e3EewqnewoEIvklvNjNIX5fPcKSw
D2o3rDFu+9egLwH+vcKncJp2xDVUgzwe1Sp34OTOmFkRulcxbkZXOyrVOJsUgA+TbPsXnk27z1Jw
CsknocKfRvBjL5JJMkVbN1ELz0ptNDP51H3RcAimh4RyMC1y3/o/ALqyI4xF0DI039J3v8xhcanX
enxxFMHkKFrrZ8TfoeUJ4sDpYBdvDt8gXIqZhtyLET1HXFUihPNJzet0usXBc32LN3yxOwP0Md2R
7OMLOnwlshrMafhiyM1XBDfj5igymBkWfE4G0EpyYBVrHJttI27TuWvdKdcXGo7IpO/vhFKWGIFF
sOMo0nHA9ihZ6Tpk4OJ4cH4fxK3gwDCVXadNGbt14r9eoxhfdju9GeDyQgEvdTYXINhr+GtndQWo
ojv+s/fki256qxZaN/Rc5nI4hxOtAFobaC2JiscRVkB1UIHn4FgOPZ2veBUoKXvRM1yGtIlKRyd0
3x5jid4DHHjm7XHhHJTKINPo1wU2odUieJwNV4D5lLz2cV5IcE3fBU+NXEDYtwLTrCeBpUaLC17x
EIfp5kXTcNI9KI823O2oj0Pju8Gm8mA0PhPtf8lSOVn6+7nGdxnrr+R562QZ/ncVQlq1V/Xb07aA
OWUC6FpuL9b6tzdQAAlAV78j+rhYsVwAFbJj/dmatTb0Pq6ArP7v+gY/CTKHzuYGhgzEpZzb0ZNv
iJI5V9JK1TbFURDoWIPiXLOXRRygeQWFHCVYQpG6PMfZMtsSHgtVLMaBXEb4+Sjl9VPzEhoxik8e
EwwYWslH7sn6LqyTRbDSt8ps6HfgVaJBZmHMstX7CEPLwDiSSBgD6b7O8hOenP0tCdS2Le36KOAO
lW+8XUmDzFzNbnL5KV2f3FdlT8KnFfSbwQZD2YU03GntqszCJ4OsTdAGY7lVqpCYwC9i8PEoT/tK
1/uvJyI8hv1ZjRt7MQPqaYi3BlpAMM+ulS9+IY4QKhl/UcINrc//AIjf8A9Cpu2+BjpwHthbkuAw
j4/2pQEN7e3hFUeHzqeyVpwJxzI1yoLaAovdrYGDzCS6HYZTiWvVunHbiiJb25VvuqchkKGotvPH
9eNMbZ0ea+J8VWPbvaBDhe+0MR8lL09WONCQ7MCQHLarfIIvK9dgvIma0VD3YAG+2VDTwv30GLDz
mvmQzqurf+jshZouYmg/fTxspZm3bJ5PEFEy8VZJmhwGD0xYWCmywS5/d8kZA6oTsqiotwTBcPsM
d0MSQO0aMpTAvcKA9A0zwThxvxCQkLLXCW0XU4ue4A7ctBUY0LCj8UXS0iWeaSejViGZVAesZpuz
sX9xCbk87KQvQt773v46mQMxCeqG85hwpgjl1AxUZALvhNfhf3WLadv+XwTYLuPSfCZiJOWGkw7l
z6EaQhIlc0+nYQEve22YySwpq+qe1b9uwOldurQDvBCOWR3q9XOxNEdZgTvbOGUnTyRAs4DDDF18
rdugOYoMUlAiD3iac6NCObmgLpgdRBpiCfVFnZ0ylinLgT31rjzMXp5Iw8LKM+n5s4HUXzfdzbCP
1obAuS+Rbb1Z0MwwMS0kz7hSagicZvnhoZ2ee4TW/DlFxek8EfDsgAht6l6xRczMTGiC5wGu9kL6
yeisiJw+/ohaZQ8mbuDSnHiDAKKM8boAT/IQrBeC5s5Du+Tx0vgIaSvaJU54G16BS5o9PTxJElrp
JbXgM3YSh68awAY32L1fwwjLhbYeqkcSBtHec74ol/i4kxeTTFoEbDaK6ZUIYQ1pVbgs1dVeAw74
Ji7iqP7/BxHrpLMVp1bgyFHnITkXm10y9Ue+a8LCVDdy7Mkv+LZrRZpTbPibd/L4UHK3QLOh0uaK
Cb6jSsDG+qPd3PaRj5iP76CIq1ZaE5vQtBLXA5kfAtQOhgSELMVRsKxMcC1B7jEhvcEWo1U9WemF
+N/hqKnUfoHUSE/ERlXniREE7Ed9sAKhfrU2QwHowtsjWhcCIl1H6IVy263wGBatbxuzDHJGs3jp
g767aG5Gvozz965pO6xN3ZwIqJXh21npEW5frQWetzw1ZyYRHhduV3Q7ZEenb4PySWmlPK/mPQys
iZGnCRAzGOKDcvfnp7+iayJWQwyEFvyYvkRwxsk189DYgBC6jpR3JRPRP/t+mInGdbvoHb7z5oEv
t76bIaHyaTjCtT756N0P0ncU2fY51ZL3cQUENzPdMgeCnSNR96/DyUfxMhn4PNU4YsmXwQ1Oh/Wv
d8n2snmZ9x3MGImLavKI5U+WsTH5O4KdC2rqKQJ0qv+450T1pomGsrz4QESWB2zyqwW6TAC6y1oi
uzg0o2TrtmqULI49cLSApKOMMRIkATD1jwBzqtb9gp+1veg4Lj3WEqSkwn/4a9ezCDfIvRSBwg8Q
xTqWy5++51lpx/4UfLICuNC/k5CvsiHbiEh5zDYp6FC5Xw35fGk/tCkBzjnMYB1yPXHQ0RBNV9Jt
9rnRbqvrNvAhTPSHRLisjVOe8G+PVHmTo3MSlm7TOGhye/+Hf1fi0Hh28Xo8Kxy72cdq40nSD7e6
jTFdArLp6nJLFdIz2NUrxtQ5DOsT4gWeXb32+pHKVWWVxrbIQkwg3Ibaa9siUfWWWjo6dyryB+Jl
1vCWeM36qjiBCWNaaR0tL56Gd4teJIRxdQOixhucJU8QgOgp5PXW9k7fEnKtJUYso7wMBQmxunrQ
hTFZMMFYYTZPamF8ZkN+/ALBMdFNWLRWCLdWwAw7P8iGc3vKXNWkZE82CrFUXE1TaPeRQ4XLc4Kx
+KJ1ftqOHWCdL9+ltR1KSjHcKyPBK3L2baSm4wOPuMEwgYnaKkIkkdeHDhYTqM7aQ7OYocfT1TJz
Yos0+/F7SVzWqfic8SWQBTg1FH4GmzlwrxDdYD9eHw6RtMFhi+JTIYQgov9MS/ukjxnNyJ6kUsFC
tbuTz0VOiVWxWCdtRDxLSx3j6Y4W9BUF6MkIsQPSPZfijpOaKHxISkJaYAM38NXu4diGK+LxaBoM
g+8+lSmrc9XalRHqcAVcGVzb6+eYLLHHYjDcoZodvNjnG+rhznT9iYmyqmbvDXmsS+zlE3nFWgwf
5EBz9mUzIk3h8LWcSSMSmnQsHxYNbNbqGNsHJ8pvOeiU4fZRcOSrs4rJWpn3dbqPs/ZvUJJPhW3q
VH+LM+5ElUtVJFfQtrVtbe8HQadTd906IRN/f45ZR++hTsyjZ1IALmdltYrwF6ED6K2w5ZpmWVJ7
aiivSh+0NmIcYW+9X04wvdhw6U3MJiJfwIYQIjlxMPnihuR2CSi4vIwJOaes/vllaM3AzOWotXA7
2BrkuoUcXJ1rAAGlfikU2LSvaIMoBqi4Jlm5f2gSepC6Pm+HYRAw8N4Pi1mHIv0SBAIe/pHJcDzn
dCQYy9RWODxzXZPcT0WyL0DNAhDymK0BCeC53bgTim/auTerATx5AhwunBwSKzU+/1C+5954klSa
TcwaPz9LECDap00ySB9cL/EWjHiC1E3TzWgPAoBjdjEwoQtW4WC9kdo9eqE0DlNl9KVkYQQ+e9I6
f4szMYrHNSEYW7KMpPXVNjkk4DNL644H0CAvkVCBfp6tsC2QLtPBkg4jVEOjz9mMfxDItW2Mh048
E/MTTvj5ybZ7ngoJbraOzCCPYubOMEXfP0JSsngnCtQXB4pxWeEzAAy9Vv0YMfXjNYTdfP7V5J7v
JkQHVPCyYyueSIFClvK25t/aay8d4eUJZDhla7/fmHO3lCsDsVbMW89CYpKAEHS8ThtSilaQwwAG
3jfRc6YZBTttAeEgp9EntjeMfs2Pj0VH6Em9Wav9wIiby1D0jvC8ReY917KAXA5BmAHt4rZuNXQw
rTRrh9CBXVGe1GiF1uWvteh4iRTNfR3zppjjNKbR6XcEmjc+ZVGzkhUOU2aOPRcyZLL+5RjyRKuy
ojB0INrAnX/eLtamjo3g+Fj895I0BmDldGh5ocIOZQZ25wc48NKCs+G8TuOy2E/xPbEinb3zrnIC
S/YiaOb48rfWqXshWOjg0ivjizZVwJSIMDdL6cHPe3+xerULCggpwrimjDr/u8tdv1Ypwz6x1h91
t8Ww4fc0WAATe+1+Gg/YsOpgpfxIers4JMuzebkeOXUb5C+Wj8KxP9Ih25Y4OBjK9uY+0oEFpd70
IE+envRCczyE5ADLVpxe8j/tpZA+t61QgzchbvooDjhhG2WoBUCgDqAmAQT3lRg4k51ySXkdrr16
BySI+Qesn6brtZLxC8RKqU7Yzrd1+zuGgn6Wb69u32l716llBa98Zzt0//ZbGlvkdXEXqrTJyRtA
C0LNgLTJyK1J5IIVtzsbvhQmWjYIGqP+75qSSU3+cVoy3QcUBKah6McjFMNCq0SLBWXpUsD3E+AK
bvcv+sieIxpdJdVkgQdP3poFBdwt7k/J9jcIq/PqwrpUZvT8ydgL5lWqDt8KDK8kiHJVcdbGtkGP
B+yCF2Hgbgk39OQCcjRxAi0hG6dxqPY37SCI8bbP5OhAafG3WfsxkfHt/71x+nmlvMFcY7F8T/YI
HnXuoWIJmGIPOaMi86ORm/7y2kCPxidbXZsSC0dbSmH7j2LDqRvEgW0lJK3Z6byXw5hu9t5KErYk
0ceKQZ9od54lCz8yiIFv9b0AF/wS5m2cnSKpQXYlRMpxVfTSa4yGPeBL3N3d+Jt/dxA2Ri1b9SzD
aA4R6teBYU3fJ+4J0PHBSG52gqQm6+liHI4vlFs/LlmXry8DgEQvJAncGyZCQRY9J4u/2xLB8gFz
X6ftqIBmIyq7lhIiGqqM4LFPp+HciNRyAnOi4HuyPX8ai+Nn1RqS6XrX+lLFpyQl99A8juZLkn//
CyR26+zeQdnIbTY5ZN8Vxnb3Be5Mk+eakpVBNhhwvp4If4ip1DEDjXN+oUEIqsGhm6Go0ftSEnHQ
Lc3uj0GndlKKSzrECtEKEdW1/g5gPIu1DrbvzYWObUuBYGl4PcT410fHbcYXMtgW2TsZqLR0bfBM
C4+MRlxwxe/LsRLs7hic2SJeJWQbq1hFBLP0rBDE4asvs1vXPrumOLyCnw+NW+Nf+EOZ+sV1OLmO
6/V/NfvYFmrBpxfNLTv98md4B6Us2bY56IuyNzfOErqiCSmJAoG4XEILZpnDCIZwLwnhEjhwdig7
Gcwdyoezn44+UxLnSaBdGv/I6TSjOpR6FD450BW1GQUOIXl6jbMitt5g5tLUwu27lebS044iDC5Q
AbpRtHjx82OdMkGslHcVesHALf3NGMWb/P+QFhA7OGiordhADCVRKfVi2u9rZ5837VgDifshldyh
WkI3P+hies6UkT7V7rkB1lNlUUk37A7E/LRJWgCuyNHkysA7Q82cae++W9vmrUeVGJpRhRWw6sU2
sn/lvX3WcdZyxBz8xxOdGvDTCAyWbGAw+0icNtEyxWXgncMRBFu4jkb3QoTuRjy5knoLKO2q7kL9
rgiFGk+PpJQ1kCQ9hprWXxp/SeIghFR0g94XpKkFFO2cVnwqCse5AfAXLeLAVr9OfpVxtVy7QcNJ
C+huryv4EN70LEtx8fW4TWXGTLQhdBo/oAH9HcE+9gKZbNTswGEzT7XpTwPi5nIq3x0gjmQka8y7
dPvlclOsxdpeWfym1wCgXwJZjpifnX2qFBu+ei/9zbCwKoTWGRHm5nPSzqrH5SlE6JjNHJN3U103
Yhcfh0tOnh/Vi3TAWK7b8f/LZ0XE3Ch2+DEsRNDMHxUXMJkOTckoUwSHxG8WtQpDHh2adwdBHu+6
VvRY6MP3ZUFiIAs3URmK3BlwT9O3+DBx677I9nY+0zItuKXsn53NQxtSQdUA2NJdQKdr8MZlMTuE
3VwC3vCCTsMdjhZ+2g133MzAk8i4fwpQVSqzEFt/lBct9dtTBUj+cN7SS5FCnw0gVGLADv9I9IjR
XwnOgBtXmHJpaYiaEREXv0T4m8swzLY1YFYxY9nupqVh1gkbANCDuRH7WnLRGrkzpOnban9fwxFX
NAjictkaLCsWQWuys9B9Jg2KUUaewCWryYD0bHjQ/Apgwgf0CaBNhDgc6J0opwKm7uLP7e6/WmWd
de0Y4MaPV9w2JHpDPWEkCtwVsdOFTpVPZpD+Ipqz+X+nJp9Vje3ZF8WQJvw/QN+ZW3/Mc13bGbLz
fsBa+fL2ufcQxXGJfWA7CAcsHa5MNaP1QFTMID1egfV7HZb2uk8gm9mbOSfSs4HZEFaM1ElpgH3z
t+QLBa19G6dBYOZbLZ5v9ZQ7wVZ6q6SWGddMrPGJOriKG7izOsGnhn1d33cjFJMpli+x4kaXP+DO
jvR4Sr6meLqlbueYftOGzByozdswadEqk7vTay4xfDs5OqP+iF/lMusfncjyAXYJDyGlkaRhCXDC
3RST98LCyeZNbXtbDTrElxElI0FQgtzOrQsFwr4M4OxdhDy8/D/Pj19tAtxwg3Nmxau1HXeFGGyM
30zTGJSSlDRIxGHoyfx0GjFKVjie1GcDpDZZANwu0+VOufZgFTmukq/GyQLylO/dOGP8xhwWK7Ri
El3jbe1aKXnCNpVdPQ0wbByxbjrR+vQ6gMnjKjxI0Uhz3PFIPI3IByFqw+WLI1KSwDZqHpZNd+CF
GLhCtUN7ibwbiHLxtnzhll3veNJZSjOfOnzRREVn4SZdUmBQOSC0meJhfms2hdxovzzjo9JcbREp
P4Xsmkr9WHAGK6uKjBYFhaIjuG/Pq6PuQ/FDKsXGD4S0ieOM0KHmx4j9VrHcY0BqQe/chwOQRUiP
bojycRGBshr9dIwoMYtssVLTT3UqV/xLs5lSpmGgSr0no7Te4KULjnJnvgH7osCteuJzfYOd731e
wJPtwKHCJ3X14fOl3PvFNTISSEkRBO2SOtRaUpXqv+TTsNqSwAeKVK5Xx9fvmZ/a1uQdV2cO/sYn
WbhhQIGQKUXm6KI02Yv4S5UK1blqeYX3tOmbSBPtnlBYZzi+OooZBFoihnq+j6LwDG9axQoHf5tj
6yekv/osVnPhExKkfG6Hg4GNeYpZsGTvsVjgAvdEnGAYA5fxyMsOrXB8kEk8vUilzT/iRm7KPhDd
nNT5rmOTF+BrKaogAwu3WAGtrXfC2oe+cZHNUwuLGk377nEyfZw9Fs/NS5e5xhZ2wLI8siAKv/yh
LVastSjIRfyrZLpyzBsDShMtHtuACHDJDFojUNxx6gGerY/QPtBAuotr68A//YV1PLPETaXqQosf
hVB9BTY/BQmSMrisYdmrjpQJp4Z98q0pDWg+3L2i3C/X7sXRIeVadzoUM2QazU+vx4LNagpNgMSk
IQFiShrVI9RxxSCKdHsk6KFZs1Z4YFdqa6mtORfnRRpxBZjFmZSu1OOluFmj1zubIIsFCb+5ir/d
DI7K6whbM54MxFM52IKf4j1QSUqC552xEg1WJRdyfwkDnYu652s+cdGWqYyo4TE73GPwJU2FLj4r
VzR5oV+NrPAg8LmmX6dwkxy++pSkONyzfvfXPXhXzoF7DH4ak3uGtiW1rt4kopm37NlxhEwBnr5L
lQc5XtDLiC06S86YS2aoxHqGK0eO2g30rDGSJEbzRghd9gGI5NqkoFdGw50BORG8u2XCgGK+2M1o
SUJqS5+k9UI6yjGy+YZF/R0kdsM8XkXm6Pp26AreJvg84AovBlaKThlAhfY4PTnccmFkL2/KL23w
Iq2y4rEWsEBmZXUp7eFLjdqh/Sb1MnNY3nNQacf37YuxVpYxFKos/C9aOQABsDQaCOXO+FEn2PG/
kPCt01GTEL63e0z+SzMHnxtiYzKNRYyiht2mpMUba+1sB7ZJMR+z86BsuJL5te3d+Js4dL/r5HvK
S5C04hfLKM+A6kME+9I5HJA/wLETCFTAQhI/vKVN6F76QuItYy2eoUXJlA9WSO+6wHuRagMvDSNK
8/C5OrIxu77rLJ4TGbR4WdS7218UPE+oGatUicnUeOfeRGgPxCYH9GbEl/LYieb5pxe88ajRW1Tv
QrNDp9eCerh+ruw6xZ9vbt1X1oa0RjuL40Dtwi9uK6s2RBrlCsC4GmI+3UNrnHFnV4CZGH/vNKLI
yby8r80K8q8XXVj5JOKU6dq0gi49rA+D57AVr4pv0TQeI7zup7v/jaj10jWuo6z9ZaELcVyTovcr
e29+qKDXoJmy+j2bqmo7n5BStGgCzR+IG0LBVB+LZNTmdNhOa4262ag1wUVrnNRGHrVcLkzpj9hE
JlgbLkniP02YHBBj7Iy9/UclmC/zklAqEgsFqhUfiVETfyXcYF+xBNvPBD3wKN6i8ZgIOz9MUpBh
Sdk8rane/uuNjZYOk1wWUVWPY4xzKYVlcAPw4sZ3ZVuZhWYjkUFTZeYThauoeSU/Zn6VK1bfdEkk
4wL+MsuYME/ArDNMi/f2jG5H4/xZZlQu28WDayzNq6hzJ9e7JLU/BAxrjzv3fEQv75+Aex2Yh0kz
BynAbOiyS1GweFlj9wRdkkO3fPUuSqupn0iUV97lmwxZCi3dAVMdTGXiHbS6sz0EWohyE8cGhzxd
txGzXW5rX2LHV/PczFRtMdLTy+0ULVi5SLJ7YqB8/xcLqfHhMf0DuFVohXeQGrfUMx7sranjmokb
mz11S4sy2teU6IDjocaD0rXpm8oEr6myAb8b1yufhcRnDxA2rFbj++lel3wvx9C66R31lxMWYIAT
geRxwNsWg1PD0iqzo1/FTfNwsiwM5LcxuNutkWDv4pPMM1dKZl0qXftnEV+mBpvPJTD0PxbtGXpp
mxl40lpJFlUOnzQlH0GDqmwy54dFkrTGbAf0UiSBOPnAGcnpiByVmkDfzWThS6sU+lf7I8uRC53k
fZXDK+eiDtNnEJ2lV0SyChabDIOmOS3XcGQhljgIIMuTOjb4HUS/GbIQmv/hCKGi0QZrxQvd5DbV
b78RtyNXnkjXJiPq1ewauOl/uH0EfTW2hhzQX2Jp1mAgp9dTfoKkiFhtLzKc1cCF0FGmKQcshe/n
ZUZV5rlxblAhyMx5jyZylAPs6/i2sJxAsGvXJPP9X4JWxphOZMNYWIHJlF0+LsxBZJb3QywaQqeR
nw0JpNCTj5kZD6InFDL+aWzO0u6Hcy7/y++oVYuUS/gEIOA8121scF3GTT2e09G2KsbfuJ4LrInY
+JmVoTmZ0E+SODxTAahivHGqN+mWAL4IMX4eDHXpffd+laIyXsTqS5RKYVv3K55yHJ+sb/RzbsUJ
cGyMHSK27hAwf4hwdEQfpkePLXunm67+dHVZQnmhY5HaKD1C2xit86aWTuozQ2eVB2kTbB+L6mHX
0uowd2aOeKpP7qKS5TtTzja4RSThFcJkcCHNXAB9HeXT2f13DENREujmHjespTdRZcN1fNt+dP/t
3aOy3bpML+Dce07nMCOPb1zmM63XhKEhcjY8nas7UA3GPpv/1eLTXTROu6HeQpmn6Jx4wYXkymF0
iNVH/1dKlA2YwfextNJhqMqZAp5RLgEFhMVJKpnH2UMmGpjaQWvFSNbTpj44OfgbhCSfaDKTExUR
51Rj75CL0uXblOJfndynPy58PvERsypEG2tDt4hJGo6GXCFITRsPDWCHiXX2+FN++rEJf5kxwSVD
vO0HMY4Mxlla4hTLVEg3fJHYl8WnNCW/p+ksy3O9TPlODzG/YbOP3TX9JHam4OqcxbL58f8jgnzm
CdnMZAnZ77JW7Gk9KL+iglUg8Q2cWoTuuEScSo3NptGxqQadBnZcno6KocVK91JzzcqNuBwBqu3O
weMhUpLxq5hiwIRoZK5kaRgaFPWE+u5Bzrf/2Lz84PHwDOaJo8FuwXpvC9c2bkISgB4lCe1DrDL/
knkOtoBeObmzmwdw/GRS84AjCeS9Znzl8fFzqSMBhA7i8KUU80MxGzvyBKdCOIqdEmtVg0hzMfPg
f2EccfRPaPNsz8r5EzhWILsTQF6GzhTTAufB6JGVhxvF3lT9rbg2fNDiV1cjxEZFti3algMYvZUx
/CGmDz8Vl266Qfs+2cYOFuc1TXMl+PXVTnIPQv85d+q25xHTx9Jv9Qdd5BJwFJGnHD8BcgXjrCx5
kuSc0OEj4mVoIUP6V0pVKCSjmCvfMmQPhNFui8PH35ywkPYM4xGcBltsKYQg0TnS0o6wgorLIj4m
6ZJUZi4H4aX9/8NPp9rzFuJ/yleqxF/vNrjDTQBBOEwchUBQA+Iy0sKhGhJhq9S7W+sq8S6YG1YG
dnwvSW1oXLy992Dymsj9JFdBMq2ss2663pp1XGu3V8oZg3DKvuC52iHtHoDlXKAlZo64PDmnJjj3
7O5EaV0LbT1VZCl8AXZ+0u+baDx6KJ06AUohevAJ71BDt49mP5Yk7o8TuqTDKxDv2D5Sykiphvck
G2DC8kaSdBpcMsKjiIBeYDaK3OJwl6XMbFjT0pI9NtO1EA4jXWqPrlp2O07H1NQQZoZZz+cM6Lgj
nBmbp/hjOvF2MBw65JJvNUcsWupw06l6eqM+Ajo46KGUGT+R7DYFCmRMrbx58zJqP/KZpDXj9/W9
jdX1nQO4hlRwaSLdWfdfh34TLhm6oxh0Lb/DXQsL0lXHjbpOqWy8gYMlVBNsNHcyTSGCKwYVFvMl
zQTXQBxQ6koAbqi015Pm4sGbDDo0dd+hUknqjbPG+RayTBmgZ4TJ6GaFAPgJQeWfiqqeZq/a15mN
mVwkXXrZ/mhKf/WKX2Xqj6gG+GkyriooloOYVnrd9VJb2mYRNWCtnEZWl+97FPrZVI4o6V6KRWZm
ZpnDMHNN5GSA4O6U6uDhUeaE7+sxmOI9wPTIY2142UzjSA/bbd+dznGIAAvddon0ro7fldd43XX8
71tlIl3FJwDRZpZW2dttVLpp+yiHDDSirSvcDxT7wKy2U+9CTvCn9bm5CCbI2JZLCvK2qp0hCpe3
BNPP9P0gYmqX8yuWwuNpsvewtu5/ECM5tWWGU9X5PDiR1GInyc/w+wP2pUEoKWkU75ntlGZVHEou
lN7RDnEF8u4fxTG8S3vLvgZAjMtI25YY98tBU8Wyr6yaB51Gwp4O/nPKDb9ZWZ0h52LTJMHoulbY
KuV6w2TZrIM1XKJzvck98Lb9/fN4wpIx7OD92P1MQ+/e2YenaCqUydyeRKa4G5cmmR6uX1+2YCMx
TVNHEALj93I2qMJ4VwPL2gAIImUJWVgTOkHZDL677n+n1w6l3ZkXef8VzR0+lc8xlSwkXadTW13I
KkufAmdupqAZjkgO0WLAWJuPJlR3CJ3JnwI5EVeot1zCfOl4ipc+xH7Oo/6jqfdBrLVkZ2nZYlTI
ryY36UJEriIgbnqCxz1+Hr1+RrXIKPAx1o4WS95HstviqmlTTH+i/uzpez4o+lZ5RBqYKQgqt7Y+
xLeJU98SAM8wd5mFn0lEjtf9sqGvTDpm7onQAYKV4PGp8O8IeVTJJWAYpx+KnrZ6zBeam/kAEG23
Hzm3VN88MtHRYaP9eKfm5dM4WSageO1eqaTehVJdgbX1ciUSEaBurrTgoiNsaWDm0iRS+VblA1SU
nintKcgdWCgeflV1hlk+bg9qL1bRSI7QMjxl34JIVOFNDZ+AtcQ1eDd0sof5uhQhX93bqEYrgAmq
RsNvXZBCFQZeiOu8n9XqU8/y2fpAobXtSUlzAXzz5zNG6rDLgEb7axf6cCv6x9K/1yYkGXBy7aK2
zfSc/F5d0B+C1Q9e1FiCan60fuIv7cd1Ex+z+7Xy86hiZ4UAWJOAmn4ZejlcO3eA+UscTb8ieVB3
uzEZ50fXLz82/7iHTNlAz0Gij+qyAnhnDo8UOp/clFzeqNTG1qY3/p3qPdQpgCaeQUEsSE/XRq0W
OCRdjhF2BlfDcDmWwgomKaRyu+SJP2vE7z6Y7yDBuITt/suQSqPQu3lA1YZhy6EOeeJVbcjJrRZw
PLIOl39lS1G7xm9InIyahlE5euX76iPoXI51uAW92zvmrh6aKABGihSujRvClfpsGtO2AScQxw4f
RMX8VxrQ23beiYME6RxHwKuSeHd/KMLZ+yPCpDuet7linvB6BKzk2Li9Ica1u6u8d+wqfckn+fvI
Bo3eBnOOwtiNbbwKKhjuoYujKlgej1vwU0kOi/qaaM3oxu9L55dWl7GYfPrUJL35ZPqGuU89he8/
680HqJVKGxukJlNTntjRF7u3IUTElqZ+1DUqIDOU4DhdR/FqWrTHvToZsFeY0KwuA79hpV+LezXf
IN+V8Tv17luzFeTg7o1GUEihctFLJoHW9a+tUWeLaHOgX4AemWzgXxiqtaRz+hemtEHm+ZQLuDIS
Kyha3kFeYedn8hEC+RDJhp+hjM45fbgCr5OOBtYHQy1T1/mja6PV74ll+MPZIpL6XZdGUYrRIAOH
7l5GSWpITNnOXT1ju6jsNKFHThpf0QuWvywUhhhHPolkxHschLhiXYQ51lm9EyE8BsftShzJ3FK0
X7yrl5kep712ctVe7TGWadd29ym4WegNdWqMH6nl/3vQ8sfurcpMlJ7v+Hsfjn+3Nvy/SBCdn0K9
n84h/FsZxDRHWMa9N9xJWw+Z2MO/u0lBY7GPUXHlPkQf/XeCzGF5j94RSHfjRCAeHBXrZAqhaz3Y
Y2AtbdS0YRBwUcgkhJOf7HEAs9TtFwEA2ed5+mUaEW6ups/y/ofcopGyy6m4WOd5+1iImddiS2mk
bIlDerEEl8lewISZls0wmH6P/c97iRBwu2gqtgmmldLWjLtUrkl7jTdnImSCGU0WH9v0rqq7ir5E
oKGjio5fJ2wYfyiGrNPNF7uricA8yezMq4i4V+/wPZ51hQAn2RsxV5OF/Rsj65I0ORqllZlGaLy6
/JwPbuqK9lF9TCoILw/tk88WbjT2dUsaXndvbmhCsmYDeZKb+SvKk7kLIVyT8UKoeML9G/Cycyt1
3pCqVH5XyPKK2+ORhHa3tEJBhg4dAeKYiOQQTsoDfsP4OZrIJ2J8SRJfVu7rr04WHXQeUQ8ogDNB
2aWgSGIVFqHuM+PlIuD4OUTnNXYdGZNWi4vgub3cp+4lwi+R2KD6UwNGVot8APgsPlR58tQnuFhj
TKcL5tK8zl0s1naQtEtH6b4ki8ILBJUTryYzzQCuf3h/aTGI8TefeQqMob3NWM8uNXnDYcB29X9/
3wT4CCcNlg2DX+3GCA+zt0XmFVbMo81NYb25x95UHNumgj25fbvf5sYSriqXPu/EBRjaRQnOt1vs
+WuVzbNeY++kLst59e/bLmCWtwb9pfYPGs5xi7M1Q00Nuhl2YDzVZHaATsjz7RwV/55w3Ne+FqHA
UdD36UiGmzHBGJRO1tAS9P+DPss3c/MhL2oEdeH7RkUCdq91GbmoQee+w8nhjw+ZtSyKRqqCUJj0
8flmLfPKihamWV0U4Qt7IsGr94+ox30/9ckPJFcpYDoPTcPcqq3HEVJIzApynTzGr1GyBJY7nyHF
wle5mg+X5NxATcWg2wWqyisIFj8DnLAERe+eI1tnReJkwq3QxoVEY1dHVmRLaK62i9yzdHSYfOqF
GD0sUNswAF/3HrkF1LtXOxiK3Mg0u/ygKwn66l/iSIR7EXjda3TVU5MU2KNPWrx5YMYJNDkCOTnk
138vt3ray2GPI9fhyQ4y4t7S3Ta5ZO3kTFV970/VmCA/wFhiL69bxK2OOi3i8/QfuP3nNsD9VXos
aw/lyiXfk7aAqo3cfcMzbrTtys0Z87SleaSbIPm64IiFkiaCxdP9tgu893Z8Ge+JZ2KOWhu21i/u
5TupwV/0cLH5mtiXaNhyrVIcOj3ofRrs2VGvMuI3CDFs8O6TipcaZL91eggGmrpdPlUZvLTC1sYB
UVzZWTmgy8HyzH2//bnqrSx8n1PChyIiZrZ+Jo4nLZpIoVfPhgx+zeSyE8B6QJpVhSWCHg1JC37g
+wyx/uSVI/HTpDBOG2hp3t0Y/pqBUNLl6U2Oy80ZwG8xOjY+YCDo4SCrMwjgMSf5jim235KyBdJZ
dbuYaifLM790TgGR5caOhOS1FC1QwUqxM8RzshE+0mLkSdrGXqey+mnfg/aDzK9LHjj4Y27HyKcl
uXsWWzizUwQI/zjGOeTblX+hdRVPMsVx1sTNFVmeYJao1PWPmweZqpoSCFLZSv7Y1DidILNubxu1
BWVVHf+4Bb4oolp5qqsXvMwkdU/gK124Sm06+MkJnovKbIcSJpZRGkLiuQnn5/s4PE49NlwENcFD
eF9xMTUzMxo6mIf2Y46WrMDpiPK8G/gBuCXAZptY0f9m/Vby6sd3lfwtDFgSpsl44F51l2zEsQNk
ix/hLp0Jf+Glebr+bzyEy6Hzai0wnPxJybtiimDH7DwHnuotFI1OTTAklZaF6JM4iVOYMYt9uQSA
1RzOlN1UJUCgnfrtOJnkJl8ASwDtQmqRxQGaMYcSp2S5xAjXZbQhaU1B1cza8T/Zdl+DTjpoOmdy
/PyilBYg19hp2OsvTMgRyRqDxBMer19n1oFRUueLVytvoU4/hcjQcDw2vev1KXLK3aCbRkpccmXH
QDCW3FJLB3Dly7LWCanD1oRkix92U2sGzWl17r/CQ9TNX61y/XtVNhl5cGKQMY3mkrtLLxQT6knj
jtiHF2klPx1Z9JAvZR+Rj54rlQ8QxWGq9WAlHWuW/gzicjMU7kHlho0xX/hWz3AnZRjrZQrnDuHT
cf4sf2Vr2IofIACdxtZQ4FF1F0JWAktxHNW3f0LO/Rg3JkKFIpjx7BgswTnKol1nHQIdN91HcdbF
uhoVC/jWxMELwG/eDftB2JZVw2taaPDMj3gbca8HlfNNdejDGivPDlQ0G2cElnc8ooAMUfwRMt9I
UR/bMscpGHKhqdfPoskq7W+c8Y3EBUmJtUonsda5+rjlh5JoIRjM4Y1RRnMPh1GWccXpfe2lBDjM
sQRLWu19a+4vYKnPf6l2tulrhvwYI4lhagNmK3QFsykO74gLgFQlqDLLV2yy2IN1gS9+j2/bkLc3
OeMnSTr/NUcb6GdaZBdkA8V2giZrJfDRRlwdm8LMbPeG2Vo3Qiq3O0I6fZrFmLuxUxhvEKZBWQJb
Yk1xDMNX+nr75xInfLFLCqu7XctfOz+8tYcn32JOYYWxAuZGHQ27I59TOZ73d205AAWW7IY/FbqG
4Kha8t7+8bcgLQRLH2zAw/zKBMRTYHIofUmRKY+yUXDXchMZA8B18ACz2+HtqaJ1+sR3fZ2BUKTd
ZZlP4jVtAIx+RxWpES6zAMO4eoZKoi6n4dAAY38jBBMNQWH0D81V0n0DjAdHyhmYgY2QjPILbRAI
J4RW0DJ0yI5oK7yg1usQFSmqTWzk9/etUBsmCOglOS+tV4i4CGfH+jvun4AAZTVxu1aszIPbHb7/
WStJKzPh00bpbRk4It20b/gCe3+sqgfEi4aXsbvc3JJSfqs6nMHG62nKZpVGann20oVCJ/r2+veH
pTiyRl7WkFebVDW2NzGRQ3Ld5ph4sS5RhnL4TrA03pDkYv+byGe2ePaYbDMX/S/VqNcKKyM/uxYS
tpPlTM/zRdfQCiA5JVlr/TzoQU0pfmqsLS9MjnIPJ8OU5s6rJ3L3BXMEg4zK18TXJwWk7AG0zaO6
5UyNFdu/FoN5djnAARmSRHBo7OEJggNdQV0vXU1t6Jipk0aKPM7K4S885LvqvaEpBOnNjLW2A9kp
DpVd3xotHwz8V8P/gAEwGCtVHQv57hh4XeXQjRvPOfh9OLnmaeij8v6Csb6LsAix6ZUUi4ytxTay
UVHECEQ7bE3twMUNVm14bFLanUPmztCmZefgH/BvsKagXVO2M2FysxXwjp2ZVZg0NyWNfSjOinJD
VmIuM3H+pZcbD2BZWDemz0SicO9vkVuRhbRgeUxN9ih7GN25P5HGoHWm9+VplUoPB0KXqW3Jye/1
LHtn9x7d5KPn+shKQMB/mwddPzpjQWINZ7Rb1eXutTbbAjar2u81d+MO9GMeO8D0QlPWPetSzR4b
Cegocf+GwQPmiy59LNn2gsNU9G2N9CQakYbFhTtbhZK9nQkOQW0QhiaBdGsJu7ULFFWCCC8Ou+E0
cWWsz3MCz4TjJoWCu325Gn9ffyRlmj+1N2WBbD3ZMoxRV/7DF3PXInYPXvPcCr4UlmKnI8cYdB/d
0b/eqWwcCSoA5Q48XGsLDb9BFsVmYJlwvqFVuxexpqxkBD0M8hW2nAa4jM/hm8bcbqVRBfGDv5gP
l1a9A327xofLzG4lUJg45Q2gYi4i3TAIlEqD8C98tD6YjThunjT81bLoNq+hoediwpoPn5VBHwA9
hKqbC56ayn9C51BPXRf3slclnKjyk6+68002SPlq8lQcpjNVdSZddLQrNwzhsYBfR0Amu8vqec8n
KAq5K19v+RVoqb8mPytNVvPjnAGSI2Z9va0CrWnAdvsA+ABWKozWzZKMbD8X4NzimuD8nWNDMdb7
Pan4uSomLH5mZidBI5rsDzk+Ot1oZmqcbmKfQxqTd4QjVCZMtePM03j2otckccHEs1BGnfZktkq3
wDGeK8l3O0t0pwj/KQldnif2HB1H42PWN4Qd5S4bNKCUN342HR1JEbIDHEZGBMHG6/nYCtGEMIhP
c3toaCv8bSiuEG5LkcM+z54jEHW7VoBcFECcaOljTAAk2SzvgGG38n2Ndh2tcN8v835wngDIWUam
Bd+P2LIPVdKAnCry0cse2452Z/KDSgTNiVUEBMWiUwRKIjxi6DUwdK4LQHbEBcuq193PycdT0o3x
wvbihgP0wMHsnB1KL3VpNq1VJEpZ0zDiWqdkeMBwbDPvh/8batVaapvQVG7qPfLAjWTayyYfVHVE
Kh45K1Gg9S75CyVHnUk+BuHHqQegmwyCzFL1fHPuIQr2LQQchCNRMcZ2TTS/BezBFSPWSL4FJKAc
jXzNV2XuPp3j8yUZGjCVoh2yz5yA30oyLyoFfM37Bk1QG+iTjuNaKG30q4cGTRfwe0efvXtsWSd3
T3E+SVvOfgFGhXCZwgJHxd4JpjEavWLrHsTSC4zlhqPro+zTKVUinTUizzAGO/wpo+TCui+C/AkN
xYSsFyCTKB0+dtRuV/oOFzCZscIKkgkySL1c7EXBe/W+U6+nmFqd45HUL3dxd7hFXNTkFCQNSs+5
/JbwrMC95pkxGC+Mfyd5QfnfgpmQH2/ekM21CGdG0KTv41lCvyAitZar/N5mbVMr08LaXHsVpycn
upDQxTpj71+DicNJTTl1NF/D6nV2c0RwMm5NWc9iYBQx7g07plJEX+n444tI+87OnbLF3oLIBEJN
1WVroGblTtrHGu4kFoAJlIK+wxoQAIJiQf6IYzv3Hf5i1lGmjOHQrqS3FDPIdhEyXZ+NIp+aStLw
6cnJ6x3wDereN9d835RF4abF2noDvv4mTNv/VI8cb9Ptfp3S6uYd/e04rfw79gnv0gty3uZxHe18
Wq+ayvrib3ktflNeIG4SazKMvdorbmqOeVWfemQzP+ufhcNykgDbAHmZSlGWIp8LlRZ/hhNLFEmU
dsoC23lF/h67a79ZfbXJjvMgR+iOWPH9ZFnL/GVzdNiiNrQGOUh6tkmejH/L5OqZICobKq3tUDDK
upnnURV1d980XQIL30FKYdwtOmCYHm9WCJ4chiucN6CLu7/wsF7hxy0mwspknYrFTSDmbv+iLO/L
DvQacCDKCtoAuT0kfXhKu9SUsxtb+ocAsmrzJiGOwkOorVCpnS6eKdbcAYa8sU16d9QdVyX/pgwl
7G7pJhGOi6u6YaQNZKrzFwvgp0E6vIEqHHFAcD/xhyMWkc6vx3P8DZ4bY0ICbuaTOEe2VKUUZVWR
PWsNdI7v/CCf8UiCkFBNC+0ZyDvQKJ76+Nx/hSW1NGpIZpBjOEnpcI2RyVusDV8HKkqcwN1vq67o
DGYxuT7+7I+FFUKkAvgr0rzZLBhNgp+x/QJICczOEHa4BfBRluhq4DAOW9elq2V6M/jBLnJafkIu
HS6ZcEU8IGMLD6WGqFiIyzZmKwPbDcjZ+G8epo3hjxIQXFw+zBUCz/GVMQv2F+yBIz4d+cVuOQMq
69I+pSdYe8QW/b2+fv8BAOz+dxKc0Bs2oZjmT+8ubZY27Oqphl4LiBa1cGNDNiJFwvROUvyguUb+
NcXkk+kYZsd19kPJPPou+onhlrfwnkU9HDxuijrIP85/Lq+4GbLemsZgWlAng4Oea/82+xDpLKzR
ATLiMMT9xAv+hjQg4ANZapzeoBsgGyxNOHo2YcEw9VHdTzlJiqXJZxAlGJTy5+ulB4ZSQgIcbOOv
VQlCaEB3OML3+yr/v9zcg53avJ11gYu9VmWSswg02eqdG/KxSyq/+KgHjkj8gp8w3WD5FcmCC8xh
Zx74bXUkyGhkqtk3s5Lmrhf+Xy8+Ja//Iu7a4QN3zUkjvMHHtlvSCKQwx6wFqc3BDj6udDCutCyq
pKEqzIhGjo6byqLjBG+EuLwZo5u5w6HD/PzBxwIxRdftOzVGgjlP6C6YeSvtG7ysLNXEIG2ltTfN
9XtkN1XomuusJ5EjaBUF0srE8/3bMeuorfHFblm4Fl+94u6qos3Ex3fnDWoKGkmyPykekuADDo+5
m/M/MJNG4qvL7Bwr2fIYPOU5r89xrfk4CYXgmtXwOC0rWy8DEiXZDdhuoyZqJIt8ekoKtMa6L+dp
q2YXNUSaY622vVEzk/DvPkdpvyou0NNt++CCOKrKf/yrXd9kF0OnJ3bzphM9Uj8otsRaZEXN/iRl
fKD+5jE7mnN+eFbIKLa6pRw1WnGZKDWimCzyt5f6MorfgiOflIvtjvgaOQ1w3CRFMZ1v/ti2ZpTG
7a5+ZPhEs8KLTnPpZfRmo4h85cbtxVk8e2BXFT45RwhBJfTFCs60LhPYIGb09MXwm8BupdxD8YXK
jEhW3E0oPSlpEingg6ZMkHw7UtVH+6JFw8T5pksVJZZWwYC81YpMq4bdqLxeslgBPPbgKgEk5GKt
ciNIREC4FILPn2WrRK6cCEvZt8SmkmFLWNtiq8jk2vcIm4EPUyk4UwCt+l+ASKnaJeYSIS0LIaEc
35bWK1uGUiM43UG4A1dp8EniuPVa0lluC7MkZXYyrDztkpZyQCItxM3y38o8ka0DsW06A146Lh70
4ptylS38wC8fapsqvMo/aR/m2KZlwFeMN88AVLCdZBwkJb3VEOmK+G1v+nry2pqexK2Kiy+yF1Nu
/OLIy/BRIqsR2MQCnuN+ptTau0M4FGxgyQbI6GLgL8PF484Pco7RFm9mvg3DKV3ppFebiBoOc9Ux
NuMaMTVT5NhzoX8VpXK/nEk41hiFNeVY9iVzrSssUsg34OlA2u6gfb9p+47/rECCT4YwlT+KW8tW
Gj3IyS3kln6oqCJPp5eQQ++OSeEEFzA1TMcf+Dnt6/vcP8dyeh7m5OUYsROSP7+u7oy3SPedK1sk
8nOCGI7Dh5u7pjhIu0d/9chrHDz+hhoFwFGjK3uZSv6UGYxw4bjArPzJXZandzORcttwnLMQdtoP
alK3zFvvpTr5M/UJVC2P1PxTU+G/W0HQDTBsopG+hajjqv+/J99rDQv52RCCBF36n5NTdzF/RVLd
XWmx83ahFAP6Z6pS2RgTlKxHcVeMu67FQ1YvMjQ+ka3aAdle2n79nQCsrY8Z080xsIl9dj4mWa8k
+8knx6tPv3QmmdRWC+oZ/y/07CLzB+EBzL8sQgpGlI+X/59W09DKVE5KQeTL9wJtDe5xsDR/fcpV
05U7mNJiWtI3ahD0SG2vdv5xAFHT3QM7YydJI3c6pwGEpfdGTsah66cFED+C6umy09p/v1mi3N8D
B43w9w/h47ExUtxYDOQsSftg18FjVKuBiLFokglmyHsHMbo9muie2gQzrQO729eGpTfWdJTxYh/M
eo93VcX+7rQ7hECNtb2GynRr/HLmWwbarjBWrSv+bhwdrcx23O+chQUEnQO8xZ4fq02vE3kvlG4H
DUF+VF4FZJb8r6d9DWzk9RGOzzFoSnRqMG7wmt66aTmXhbKkH22MBmKPdh6V/o+iq/BwZdLto0oo
pUo/q4lqtM6Cd4Lsv2NZb0ujzPbKNfsmbX2OU8GCRLnvkPCJKyPb0v9Hq9PlxRM++05we1SGFyOH
DhFoiazRniSooqZ2fOLo9cqFoYphU2giU8FTYS5RIpHZnw8sncFzwdGr5+GpinT2FM59y3VuphLk
g5I6ueRXvLoeCNwEZEZwRf58J7sD/hKEQJCVqyjYp5k3lCF0cQ2fCiCxERtxNpW/kLfAZP5X1/Fb
l/6NH2sJTgt3di6FRTkjBvRVBMLn5+5UpR1iRg+OvzU0ygDZ5nPiz6emvz2sdzTmhYjIozbGt3nX
evjEr2jCt0DydHc8QkfmU/P6pYroD//w6duggRrloopYtskc5bmmOZr5fmQx9NuMmpvvJtdbcC3l
MticUjUl+cCUs3ouP0EaMXllEdjJde7bmCaw0lpiQdclvsIHr3BdCXIr9dOnxPmufK54necX8r3w
8wzSCgd94F6Ogjme27Ojcurth5wuTZCnuY6GSbD4pAhtu4FDP6E0WGmQTEtUNodonfr8SmhlQZRm
txgGhNixXKNtrkSbbHQ+VNFgj/PKD4MbrZkqdpZjY0b5op7CIU/SX56T5z/hnom3UXKKcsvLp56L
FacB/qVOtXkwq3WDNd8OqpjmoFsfmgt3fTMsrq3wwTHN2vKWTa1YvLIiTm2NZN5tkJkg3+qwY/CC
IMi4uIjPBBIvK6MusP6NdqnWDYFI4qoBvsWoNaW0C2stNo5dHR2EwNvR6xJso+oBezgCY9UNlbRu
Ha4N78UlbOj3hnlUPcOjxotI/flXeSNUgfErXiqBE32InAezNQ/D55sS8h1fi3jxonnvE1khFtGc
4dKrYv5yYwuTjP3/FWa7qf3N5/uw0GWIT/JaNNjWu7kBCePXuQKrvqOMfA5KDj5fznDd7tPcvHz8
rpUlKiuPitkhyoohNRWRgvpSWmGvATH5tk0lvF2B/0et0oWEEVvIh0yvK1fUrsnyr3Udq4Ce/4po
bn7ojbcXgcCnCswVwAiUqcgNGYqcakvFG88enaSDc1Tuno+VJ+vjQL73VhqAW1yOwGKNYPFWy6to
rSqiclHSsbIndsMt5vA2XzUlhYaoeLxTOs5T/TH1FS7su5sIpELwpQvrEUZsdcpmF01Lu6sq8NKM
IFxrzIGsBsSH08ER/49Gq8rFlfHaUQOZi0eWrIJ/Oumz553qeqbOY9nU/3h41UVpCZf6ITpmidA+
F9efcBNkWoscIdcOaheHLlD1yAAQaRc3GIRUCuxvpY56l+KAHGU3TswvXWhoPo9QZvEIyw37+b0x
CS2KJf5McCHibIqw7zMeA5OTY/7p8oM1MVAZSX/g/uuWyg8lvTB5PrcPBBjQJz9K+lftJfZq4Rc5
XiklzPDGy4o5u5oWHlqTK2dsCJmHiF+oOMxoZyrfv4bMV0bYwgiNEgUiZre+nqPMqISIxsf+2voY
xh1ijoEmeP8QBwrLYElvulQeFrRe5nW9OJRp9ctkUGHvgtt4gMA4NrL4kOX+03gkqIjHyhxR4ot6
Tt4wwxu1Gq671F4lW2HC7/FeRAs+a458ilAB7xqolFOVeDB17t6ZcnRvOEHUkV6XHVve0W56Ouu5
CjJsWSQRR2HvGzp44mRKGuRDVbt/uZ1Toeou2bWiJ4U9BMUFceWz+uMIYZvWqoCJ1ZSb1t3+mvCd
eLFl9/KAZDzzaAKNC2gIKWw9cCnfM2PJyzT2yobywA58HxT/LE4lSl6ZdlXOkIEJ5GAG/caMSCPw
4rhGHzxbnwu1b0HOqZ/L+zvMRAnLcscc99fwWKhgVsV7BTh2O7fDiQE33mvKAfjl39gIkgEu+3G8
A8lr6mffGnIw/C+i/bhlp+rk2yeRQGKkJAN6HmPS2XMzvWPEF+zLsixsumSgVm/83jplZjns30Qa
9pfEneNhRk3g4dBTmzVL4/dsBKNuj3+xpBzSLy/jLqx/rscCkouGABWVuv0aodDEn0Re/LGF/zCM
FivhDab/bA8rKHjcjnNzYNdcQ7539rsxAWQh/R8NZBDwpsRqopNWV0OiyLtJqSyuStthV2/cKGp1
rnRmfGr/NvCVUIydOtworeTQom/fwmQ2pvgTzE62Obur1igV+zc7um7pUO2Ttx63TiEE3CTXuT13
BAzQ1MqcOPWiw2I/0EWylqTFZpN76EYijjK3SR++CLhrAndRzO08B4Pqs2ni7g4NhH4vDIpvi5TT
YowLQjPz3vtD2BD/Bj7E4/zNyrjEwMGFPmrjZfD0akybMPHODQTu2p9Z8+9BtG4Nme9YleYMS/Zg
WAti8ZDgc9fgXxMYcY5Ng4ZbxuQSiPxx9r+xnDdso4MrzB6vHXbrLYS7oWeZHyrKYuPGR2cPqcUP
lj54nVbynV4pzrqrZ/+HYtYncqgTTaT71hHRKK+swVqUjdC8qLkUBS+bd0tT4cPet/eA9QRS0aSd
2hqQ6lInIJwGvzbPRkpNn7By14kI3sh4brEFXTOqk1WqgXIruw7Vg6LD5kL3k/syfs58NcMzHrpA
cIXe8I25rmh8Mj916BrSGYhbzFkSUgczs7+nbIbP4TOS9N7Z2ZmebTXw/woGKpi+/W6SLmZUefpS
qFJNX55Kh1ZJ4fU47vn0zKXc1FrGoDYBWTnT5iEYjncdWBt583SCouQFHbdlC2fPeizf85kMPwR3
24XkOtlCailgU5T3mKuxyrTWKcmsvn8oWIemHCUWJTKliIyWBu/1Bl8KETVZgc1Aa0ivVxmm5x8/
N3Zq1rnvWojqO72eGVjBu+iq8Gqw5sPeiWz8y8jKerKyFdZEABEaqwaY0BWo9Phn9bjJZDxw20gP
Wzz3iS3XjNRmgqeQDoxBwWQho/hOWcUI53gfxscFnP6doInakaKAYMmrEFt+ySdDjBRCvHUPMq1Z
tc9V6NGLe+G8gGUByQFC+noHHUpx4L9Zhpy7GDsxCh/+H6hciyjrgTSRuaSD6FBNCndxaP5d+5xT
FmzOgLtVvIs2X9vXABJcUWYew6NLePv3peONUayHuzSS0Dz1e0syCvh1eG2t4EpqXY2lyUBJ4UVn
UfWbXuyiExOLftRcU0v5y7VR07e6kMICxVpoB1na6KZ7VzQu3rEGw9YH+4ldf7Hh+ttqlDeiNg1s
tOE693BKpZX+Dl6IUgnb+NbT1M1+ksNX/0WJ+xlye4zdRvYcEjq64dnCtISsZHtDOVDwSTBImXCj
uMNXHw/AIOTrY90ncSjAR8dNSNgfHFHW+Dg3syc9IGfk9xahrbvfgI+CK16NkoyE67B2PseXcpwI
/MZVV3E9KP380r8OBxj0flFiuKSoiAiIrPHY0ZwJ+iDvfepy1br9KEm3XEQtLc3aS/7dwkEB3Jx4
CZaHbEbaXT+ziCEQHo4INFqL78edKjrh+OUr1DtOS6hBApLA9G3wBxMjQGUQO7Nq+3anxNCHKKp5
FVuloEyFcmzAKo7YJkKG8Id/l9EnIJZagvi2NHEyM6M5kzIMYbE8VDHoAhe8wjZERSjoVI6Phfsp
kap/Rbo+B3zpmHLZgGSfUxHsfJhgUMCAAUddy/0yXgaB3r/Cfs9ikJ0diwz7xwlW0Q5OTd0qKyh4
MbFhyDOGHukOyNdPUou+grIOGSHz72ULhvAIa5wgE6y2bw2eP9SWSrzU7PrIZ/hA/NXeLjefAgLf
NZs+gAaqnQ+bVoHxwZfE+ltZibNCExNwiShFbV7+jR/VD5X60VJClveUT05YSWwOh45cA7u5q0AU
+IxazyNRNPXgGHT7fcNm6AOW22nNENiYiLduFTsaNnKs+I5zUZQNVlIr/54/YLyb6eCIMjiQMinn
HZfuhUc9qHcsvwNqU3m030Vnl4pzvUW3lSEgUhMZCPBb5y1Fhd0PFta9jU2rbAkcUbj9amwSKR98
wzV/JYQUdW9CsfdO2Hf9kHPIAenOgj0DdEU9TEZMa9vMR/Rbng7KFgyT2U3TyEfCDBoY9xBwc9Vv
QoMq0P6C+H26BAffVVQlJMRgeH42sI4MBcIlxwQQsn+7CrX5ytuiiAd9J5IuT/Kpvh0wM1bfIw2o
deP5mX75qCTu8fv7w9vDzH7oQmK4mhltPWJlwQpD8YaVo6mF6sLvEj5itsixDEcXF/B2/juUo7zT
u1kM4VPdpHZVIA0B0qBFhozGRGU3oKpGfsJnnRuubLJvbNEQEjxB+ie+7eUzEZRQQ/+qwP3BVwgK
DcAv9f1xo32SczaWTH0cv5f1uLD3mw/1Xiz+0Y8LQQZQGD0TG5AFObswck4vaAn0JirfIySBfX1e
mcCkxIOk/a8uAyHgBpBSkorm61TDtlJpu1TUYOU+spRh7Q7r1Mizb5ijCKHs7DrY5vf8ymALMB/K
jP32MsIOTx7cS1OVIpq7e0cuwumDOubT+tQuA8+a16szTn7a7J5myF/P9uhqLjC1H3qwvdEc4wax
zKbk4hMAfYv1DobR8kMyMYxnrAt1oeZE5frQcKaKfKGoFAPFamQhVUkhRwpNtxFdo72KORZARQfA
G4nY5w1/qiMAX8GT+G0bDdbozF8olTgCuqK4MZ9CFYKKS47Vs7NSkviyzlN7n0prssPMlJj2G4c+
YJokxpEpI9l274Pfwepf6elcZkJB4nlR04Rdq+oef93uIOCXvfWZMgb2ldDn94VSGn2w2cbaA+PJ
p5dZxSfDaE3bBvkM96HoMKm/qydd7nFUukDxKe6pVsSNIEFoPrY0gp1pjgMe+Jgg64rJBwGLDt12
YQeIxItl3yynXUSD3yLABbyTiHJPJ4EGF2u6ykAsB2rlXBh0wvxXdlho49qieNuew+7poupGn3cT
MJX77jN0M09o7PHaLxx+I92b0weIuf7Uk4t2Q3QTvu6F2R7I4EQGcMw+VOgubV40/98/PM4YPfFP
xRtqH3s2w4876+R1wnpvO+6L5zbCkIFujWmwMjfnha1H8OyMVXIeSx2FxWykVcvATG22c122Z77M
KeMVIEdD5nBHXlHd4VOzOUTWsYe0SEPETAFkJhPzKnFPge9Ar4Z4bML4bk1as4GRT1Ogl27LM6se
klXjCdFSUgr4lAlf+RGNVIo7DRm5ZYvlmD0DJghooJuyvVVySzjNDuPrI4o3g9wAfKnA4ABe2VOs
qhNyTWBuj7uv9KrF3s3gMR5laianApovMHY6E6/XIJdk0q75+LVIa07eqGfFWsUGcG9AQbJVgpRB
BjjwjZ/ceDVANQpZD4YZ3ChEkVG7dIW/3Cn+fWRddt2QcW/iWDhdKP7LQoae+o4gopl0vXx48xQw
+Xwv0GA5+x+JonB17RS/1wZlj6uat1/SwETq1OPQNwA0a2WyKU7X43hvQDpWb8uQBovmwvpS0qZ+
77Jon39FLUSTD20MZqDqXcuEQJKr9cjtCRofVw94hkVLiu3mKE6iBBIYCBVSgg047i2N3Ye8xocV
gpb52b1jJjH1Hof/UgxMyMwZe5UGqGdUuIV36pP95CoYfDXeNW/5Q6M7XZaLLcw7Ar1CyckTfuAG
vs/oV4743YTXfgni6ZYca+KTAaDecBpLl2qE+Ed0Q7IrkthypYz/VOjevqpyXe+YQ0id+fvdujHN
r/UY7jtOW2Wav0LgSMljuezxsb3NtkxFUFNCXGlevFTFyI23m9SxosmliDVhGv7Vm1Hz78HGoOJt
JCP2WGutmV2KjzGXruiqxwnaT3/WR6BbBJtd4nTVqSLPIr3Omd1hpMZ2/mc9ESxdNDonBTxAT0IF
B9/WjElgXaCmP/BCZAjfsOusvJEErwXbVTkeS70brKVWcbREqz6CvuzBQ3FOe/ldUAg+W7C/lk/Z
vjBPG+AG9gmJzJ5jOPPVIvldCmtoH6uq/eXwiif1Mxos5cw5GISzU6my4GsIobWD6YWzcieAieGD
P9bphIXKgW2zBJhnAHWXEjmNCFzWaG6Aj3pjga0RQ9KcFV5cxOwlWAXaj+JwKFe7W15pm8PT6mpY
ha7+qmcxHnnqCWOyvbfSAxOfHcrRwTOYnGu77Jo3E2w9ulfpOxjyC4308PeAIsupBcqT0vgqHrO5
HA+42wNMQgr2XzuHd+nvdGgnM54HZ2xfqsMQzFIhLPbHn5Z1gIPof8F1S2OUYArMCZv2YtuNalUR
SqYN1YlnGlTQZo8h9vSG8S/+F9/KNJQ+gWCCD9ZDt9LFhDw5Jheh/D5arKOXj4wv9c36XjWndIn8
rH+Vis5EYuYi6/+TcaRRG9piQGuJba84SCMf3/wzR93GTea6YybHe5W3FxoQtf5vG/H6o7fbb9iI
opX3HjJqfchCfGTyK9W3sSHlsxd48Ms7PDKAigBAivD1dwdgfnHPnZgXLDNd3AksPHUUPzLCxeZM
VcN4jtO5O02Twbj6zp4dgDEjGX5QaH474t22fk0OXdLPu67CTT6aRJ8mAXOPnzklVCwGZXxsIcg2
NS1EA93GpALLIz0H3FcoXrqXuLsId0chI73TJIU6xvY3K0Y0CaeMAyJHbjZgfr0AceodaGHTYbSU
HOaDcrAzr2f1FCubPL28+sHHNC1pTviPbyKL5pAKesZPaxI86BfarGuZ3q7jUvjbbsF43fvsFhgu
r/A1WR2GJqO2VCD506Zbr8i9bTrSUtt4ojRZuqz9ByhGIGuSGQ4KsFeds7l2ASqhXh1ifVZf/MGD
+fx0SY4YRTgMrmKMpJ6l4XZe/Ol/zOs6+5Xd6AhWU49YPphcnRmuKxfj5M1rfcE+ntf2o4PLAMHH
AnTfdTjpqMp7VilOmJflmRE5+SpbI0UYKOk9aIxvYxLcjtoqhRynPNVvlRMKSEARx1+bAOcrLd0b
mJC7yfVHt3AkWCnjWfsJFhfPuO6sIGTp7jvVHKn69DCW/qJGhyh4MUh4YMkyEW0MFWeQbATBX92d
88c2BjhNxqorWdIsdI+/f6KQP94zgJCL5Csk5X82SURSLgMCiCWz9Ah5003V+iYrS1XNWzqKzXFS
Z5gKAii/7A1BBijdPVYFsItpwSbiC/LctiRRKnFbqGjuJzjLm/1LE1gQRcLtEG9+KsxWRR2LQV6S
aIEja8bwgYjorgKJfzJiDGwwvo4EgDfdQwRvLfXVGTxqrqZr+tf4tseV31PwmgpR67Vhiquggk9a
BXhiCcG/XTIYZ/T5ld+g1H9Hjrc6qevy6Oow3jnIZ5zjknQrQo/IdKvwvBTdkDcMdrHPNzUE+0Kp
GBSyi1yd7a5ayVccChCBbc2iszacp0iiKcvNMVQPZPhPaz9yodR6KJ6QWiFBWfCKjsDH4RH2bjLV
SUGRjCxadasYkpOVugwsTPcW1yrrdCUOEYtxGYKk984E0I570skjzRSiCQiBGyi2l66cv+fijHxw
y3lg5/vsM2RZeVihct6ropIClXV7pedXhezKMnqEaT8zEjORFcRJL75TSPrp96fwWoZOOWwKplDK
g+6kOeZ9+Of6HtBSEXWiCm4G2+KUFfHs70koFNqHq0XxwdCH5eRDYAr2MVraUO2VrK5PMDSwnURp
yG153NRTUzib2j/r3VOaUhqjOtFGLx3QHTkSpr4RpL7a/3rr8rK56tsxgbNvlME1MrvYO3u5jS2o
+ELGNRI2y2WZOTbZ1WNS0HAAoVpbIwVIK4d6RR1IlJ4xRHVVLWSWHrclMO9rkUC2KX8CobZxbvCk
VC7Oe/zCr63usGxmOuXiNSWiACcVdOJrLlMoOigMSQKOvqS5V/uiCdIrIkwX5XJgA2wyYLoMtg6I
TtB72dbBunhnJCjdoum8e1pmDtQ37AyafX3qUc3+JQJiZtC2/RSxymSNoZW+Wlt6cBQO/dEdhMCy
19SsDhYixa0AKpOcrWW0aEgEm/H9kuy1KwbgHacq0JK8TAIE8A+qbdmRWRvoWjSNI5ZT49dawELt
Wigltra5aXtkh28eqgcEYSGixVJWDUNztXIPKHp+d8gi3rh95tyXXx1VDWs2AktaepQnfM21mBsj
0w5Mf3grTy8pY8towR4L95jPK8jeQN5WWgvJBE7J/1PKwy/0imx4nHkduKHoUjcc/4Y3xvoEQkKo
9vFXqogEVu9CnWbitHvh+Wt+tTkT4eW6VCyK3oxfsp8Ud61CC0Ndk8RUCNkcUya3TLhev/H6T0J8
opstwOslAb0V2Mt3P/hrvI5Rzc+oNzeclZPHR/f0W5TncIV/xwz6tL1KGkBdQlwf5unmXbYB7hGU
jNqEHULdXl4+oHsJ0DS74d0Lvkvkm3GUj8cg6ROYuSU53DWCrZzusD5PBV6RHGqFW0g3cDbV9OBg
nRRPzj1M/zOkfXdI+bP+I2ql5MJX/kTJ9IERq7e1d0wIty2xS7JZRN9gdJ4u/pPgq4uaR0i+IFJ5
4H9+Vocs1nqi2twnqlbhIJoFf1CUUwVvjalbhjr86VH4rntQIRuTplc+W2/fkPRC45V6ekZ6qWoc
RJaIFK9aBqJtEXnvezHOkoo6785Fp5PhiBlSOxFdYzClce2N+1c3r3UVRkWJ9uvVJG9CQLGZRkkO
MT8cC6KpWTAVsCFKbbInAGbXLofo+IbABccMbpi2PYxiRcqb+KOILD8egeTy5BzLtOwXQX5Krzv6
HI6o0ic+ekWZw0LwGAIA7ugQr87h96Wawf2UpL7YveCrxjK4aRx/iwumMtr9kDYcLYx+DRHDCJek
qSh0DD8rGHK0zMahEd1swufSdlWh1SC6Wl9V4rexDwwKEA26KVW9FtrlSTIxWwcdS6Umag5Y+znL
N+eMj3GxxndbieVW1kro+qCuFj26OF3A/x0WnQBy1npIx+y4xrkQOPkhLd/Apz8J13vBp+lybm9I
Ei4G9/d2k2FIXnhNHKT0z367rBeMfn4rfxsEGmWDA4XmyyrXVlwhjwqcbFFA3ZAzdWQ3YX3JCxIJ
aaqfplQ8qZkuDcwmmWwj6BuDIDfCcaw/DGggA98f0Xcx6DGIRYjV1xTJAgD/T4AWkuZnxDg8aihy
wXK6J8CuV1jJwjP/WLcMj54PftX0W2iMltn5K7ajTRWlMYNuQ2EcXJiuQ3capeWi7wu21jviFxAF
8ZdIdTBxIaGsUAkBt6PMQLpcEVcc5Z0olxIgbAP2njmq/A8gDS+z/yrbjcBOHNeyO2AxpHhG2Kzy
p81wsSM+YJ/CTC+XSJegTnlb7rIC4dpb+MEu3NUDieRdvvm3rdWcg0K/fH7ocw9mq1G2u1uF5/Vo
MTiSytuR8J04Px2b3Z21t/QbumM/OQDxCDdmqNdMVYWME+c3L+eJ7BSVYHPUq2JtkzU1lvWHOHTB
QOLkgXKM7c8dpHG+Io6A0dTTxkwbT5ilQIsVjqjTQOzKhdEXCp7NJ/CKALzfCZQo39yNW/c0XaIF
LmflS9ggNdbPHP0VVkdq+qjHT+ybXK4BpCkMefPvrbM7QPwhZLHcZI+V11IvzjBkAl4U+Z2VmUex
JXH0p3SD/4o5B2nBBmcUGcWaCzvdUw4/N1c58wLQOlVsPA7QzpEMFGLhFojM3vhT0i1IH4Z9atNj
5fo3xDwAyGbSPkDR4cfA/Uj/InBs9ZZqUhys2yQ6riRFritk6JYoroFZNuEgm8X8D1DT1eLIutwA
/mrbm7wMEj9M2ekDCx2hLYf33ENKIDsrhpUL6G/iqMINfvBj5lpyDZdpWXJ2JF8FdGo9scqMbOff
3L1ceMkruiVDXVqrSFAKMHbhOn0KNBE5WJip7GUI6C9oblEUu+3biDEgi14y9KkuzzN78E7CwWuR
HuYRB0d399lE6B5+BE6NQte8GD1Qpk+4SL4ZRl5hcY3+u3M7CnCsbItjbdLdUZt3H6QM03RvBKm2
95lqxdVj9m1bTjRJcpbbDieKUFiscKSCO1kE1Ar95Ih2zUJZWj7Xp3OFmhLeJpTdgBdBtiq3PS0i
Bgn6Y0iMtwbjK/EViDS1cscPPU89XjkV2btgU8VHhSKMAoo2Zs+lS3Ld7sLoXvlRr4UKt6yM/2VZ
7XbF73pxSo16EO+h8WGop2qA4K5/8qul4cIGvAA044eS92LwyzTL7HQY+xPr0aSp7m7JkKHnsX+D
rvebBEQ0g9cJpRSLtIWqunnWbqt1zsPDfCqF7IGCdSz7ZZ2YtiNnthZANRRRF6AKlV6bSmqyhIX1
TLCHy31Kf95r2ysdfnHMvh8ED52hQwyYToFiJJgftjt9T801nhWYo7RU3XX+cULPOAguAHgOSg1A
fePqhoNtJ8sZMuS5bEtiPFfXUc6S/8vaa5LoMJoSK1RuMg72yzP+lLWEMKmNWY5lFhZrV0k5XIIM
IazFdxNau9ZJaXSZUJPxbdQApEFOcqytBIxEegArY5sgtnP66lAa7tfvP9/2bsGa9I1DIhap6lP5
FHP74xUpt7yyQvpWt1HRs1zK1gwCf9syLuoj2ek6eXD2FPQGtogZJ8Iz0k8+uWwylzD2WxkIr5NB
KxnQuBZU69lyZ3Ph1qVFstS8WT9YLpbl6najZ2HUgqYs4+m1Btqk++6v8P4FOFPDcb1HJFImGbn1
5Nq39sApBQItCKkWKztSbvX6BUS14/TDJLzrP4upK0efLCr72rU+KVRDgHwKxT/2DxIK9bqOZTru
7F8oUlbbWA7/g9xcFW5AuBJNkG9Hd1yui/KtBrAWljo3epeGZY2Jsq3PyhUUxNlPXghy0oZFwiRh
VEI1BK6Y40902F0bPAYb6LpoysgoivOXAhMmsX3bR2KMouK/pIUtCDSkCliNUQBuxNm07cjQKwS+
icp5K3ECMOeLE2/fULZnaJeqZ55cEvQAwZdRpj7SzcP21f1gJcyrJ7EyIdxkUEU4lATG/vcAsZj8
iaS6hbF2a1SkZNY4VyQeKo0PYNXzu17Xnxl8jGho2PjkUycLHesf4IocLrkhi3BUBuQbQXHPLQI/
abgze5sEnYLeDTWIubv+AWuCr3cgwiLCPGPk3n9ffORs1KTN+LE5dCgiBL6MRXto0l2C1o1Gx2mT
323Mj86t3Fn/rkPUORHU7+x3atNQrNPig5Y9pBQfAqhgI5XYpINbfshGLnTRPpTu5PyDemgZuGVK
li3DUeWGFo2eS4WWQ9ZM4mYs51HV7nyX5Xk+4BO7aoJqj/xrOj/wwN5KomzdewWmqL5ggaAzXh17
OBCcR9DGlysYlKAwkNr3i4ybZ7VhIYc1i7XhIiw4x3UwwUHLP5ONbWEL4xqyH1rQu5ncWsvYUcuf
Kj+ye958XhVU8y1AH6vVD+Iv5BoinLhK9NOlyYSX9WnRLjE5FLOIHy4FpZB9QDJmshMxiQvbcsyG
iG8yE+EB+BWpXtqX/r366zmjkFC8BpwShyJJnje8iuMNbgUHdsQ4XApuuo7mw8DimYP72ZtHRjQ2
BQAsKy2FNVqnR0gDM1cytUVoI0NB334vaR0ALmHvsylEeE/Fn4hOHM5Tp4nwkgQSbGqKsy4GUyBF
wQRp8pA/utCpM3gJoJLtJ6TUE6ltIvKcZD7EeHQ6YNk9vqWEC5Udm2GtqjB80u133LhvOhqayctD
JU8/8eHlwK0TOm3g551j4ffee+T52PESi5BXu2kABkgZW5dQvLtY8ElvoA+K1lT3lfZdLCCV/J+G
qxD5Z/l62c97LeHlQOC3BE2FYduC9hLP1qCVJI3zViUtzyvFCP6WMkInWHTTtAmUj5q9D1j21f7x
VA3UaNawVgGdV2CEQyBYLSIjgEl7Uxb6+baVrQtLMVlPUbheCdk2P+ODbtCrcj27IOnKn0oLHWP6
BAEb/96UDj9I2wpb3lJqYtadSEhlSMToCwQNR4fQhL3LssV1nq9cxsM1NgOU2dgseaFO+TJ/nMS8
sgpfPGqlQ3ywT6MFKe+IeSgWzJfHnamIdM9+HeeurGPbpjbABFL8avl5X6yeCFrhNOlZThAy/Ysg
bJ7Hd/gYKf5kmsLIE3sWTw0wT1sjAQM3i7jd1oHMEFD1Ogx18cFykEaNBVU4hVOUL3gIXGbyhqTK
4yaUCkwSmZQaeNiLIBuasF7hobv2bgX6gD8kIBLzHP1YEte2dikx0g1TkKND52yUEBmJMtweqKlg
Q7rQS4TDXKibBClUS+XcUYIfO4LTupMoCtbFrijQi/irWJha2c0U6li24zzyi2NI3ZAPyLgV1lN/
Gy1CrjhQPFnVwecCm7ayGCf/71c6CfrvpeF8ss6O0rDFRUl/MOs/OoANWmHB4SdMggKaIVp9GDbV
gQJtF/sGw6ij2r4Pxdo3Bz+H34+DekWx5SUVx3cJw2WOQOhKUkbho35nQzz5shbYGjpzmrMolaeQ
pii7PDuL+CwXu7+37ecAv9adJnUWrPOCu2NGU7sVQ2wjkRjw5A7Zupztb4HhD+/hdmcMa0+jhuQH
zeUbpOY1NRhtQB7hoiZ1yv7NZOtHJGaGehyFIqkFEXvcQzW9OtpL944YqRMKyUgfu016PMQtSGOb
rX+z8saclVlG6uSDvgsVejSgmEXmtdQnj/6oRtGy8jGiPxeDN7iy4R7tq1kFAIWGc6RsrUO+IStM
YZ36ztZ/1+0tisz6C36hdT91dl9AQ7K5XcjS5oWVudjnsRJtw31niMuJr8eIUyS3kSn39lrnVTLN
VdXaxsw8Jy0crHJI/x6wBvn0O+1kqyt7YwnfPYQUTqF0OkVbG+lKJxxC+nECPIaGms9mlPG/6kVX
vV84Hruf/QAOHpFdaIAzntbR+3yfDDZ1cLAfo/W9GpTiHeTCMSWMNRBcy4EO0p4sE9IbLTJE3CJC
BiX3qSCZdnvLZyrkhRNKehwYMqEkAoM2KT9QQMWpAU2hhm0NXGahRgrrX/a5xokBJCrmm8kk/uqJ
QQhcVxwsp/6wv9Aro7CrGmboShBISVsxgtGEuTT2vxg61qC0UwTGqbTFBfQbXDY5IdvnxL9gpaXV
A4PDizwCG8oOUZoA+khFgGijQbmAYTJw0iSFbfBaBgO8+gkK/ysZx1CpjNazR2bTTiWZ/QdIxru5
kec3WiTIOh26TNNkz4DI49bxMP6Euo7HfApWFkdliB3voEexyLdIOFLps68AHgE+dgrJRC+49Pi4
VKc1Uq5HTRuRPz3SKWEPK1XSQ+jyNgh+bykjmCYO5zQRkBbk0EqtdXzx4bTDmWUQAuQoTLTkzq78
hZKd2FRk/RBL3NQfI3rOD14XsWX6zhtyqH3uR15cdn6uirJSrFj+EywcN+XKVdXXXDcu7yDxFQDG
tF2EZ3nu7cluHlHK6hZ8nxCH0wSVSqvfhz0WQeMDqWSt4JDsFu21kTzHSw+0T3vkoZe9zejI5SiZ
qhaGXcZFcYgKlQfpT38XcmgFr/5zT1xpk6APDE8J0Y0YjAiCZ2lyqtgt0ol96VVYQGkxCAitTetX
TpL5mpheO02Ie4Y+soeAV8/HqLv5w/iyOXSmTNaP6VdMcwEGD7Rt4OSNwDRuWvqEUUryNoaBhf8i
cMeuTowvD++fMKIMlj0vRyL+E3XaZnksJ38dppescYprMLI19fPvUBxHC2r18KTffqHfquwG0a+v
nPC5KhVogY/fFU8qrE8YX+YwVRMr5d/rf3jjOMRF7kcQE7v2KPKLaC5m8fcyTjq5K9QM5N7bKeNU
inKiq61MH+u6psaoq0Cp1fXNgYyI45lZ85G/K8dflr1e2sJ2jVZ0L3AfM/x/XzuM3uPXMNEt2giM
HS1SLdp1zW5aLgF5GDbJNBl/1Yzv30wiwAZzLLpEnqvjUCUiHcieQtOQuQAh57xwdtvAxl7i9i9b
NT4AYxbR4f8CqDskHr3Jt+GO9jFxMtz/MbjJSxfyp9YtLWzSB6jAfHxnyUmyZ1m2cuVkpAYt+2j3
bK4YSUpwU29Q+lJjMRakzzQppbtfc93yY8cDFqPxs/SFqy5SXMz9182aLqHU7jnOXfx5gZ1o52W7
UEEym91gP7G43cW9g6x2ykRhgnHSV1CgV7CHPCRC+aN+9rwQBXCNePgcugr2SSJ65CqMb34Cij4K
YT4/8Ro3pc9sIpdQgGpg+cPSYLZp2oemfL0VJiYMlbZlTtNGVNBmWYJGMM84dtGRwG4F/qffbxVS
Yp2wXjj0y3F07hDrFIA8JYdx/wdsG7H8WiPAETUKTcCv7QX4amokL2NZPgnwjO16hEofiTLVIUay
GWigarP+CUVY+TOCq6Uj6Qkfz5ta9h7YQaLD7fYrfYbQTgREGrKh2R/LwpHwMJ0BAHDLjo2ktt4T
7OcThpv8diGtyAaZiq/cYSaQB4aWXaj6W4p42mc02IIhtQJZT+hlVGh1066gwNISNPRuTDx3L53r
S5reDZgdRN5y4BCUi0NxIf8CGea8oYYb1ukjzjzkfD18wMNXyS4WO3wccAwVjcFE83lf9WW5RZMl
WfBK1vCqnQhc1YWFJPSReGkkDvZg+e3sd05wUtW6GpCoGYioXb9VNHcfQm3It3L06UV1Ca7jeOKK
ycBx0qYSDKS57ikGg7wdDgUOTsUwKDVfsqEZAs0SuAnJ6MOv/HGFTpl3Lxqu7vTBzTGACc2FfxcA
TUpn7Xe5HVDRtwIHTqNHdZ/AMJL6Ot9h3W3Vtv7gYkfAGarfGXzCJeKa4yCfi5aGJPYHPW4/UTkU
b4b5p9eACYLK8xbx5R7sF4ebjhr33MtHwihwPwBoE5BkUukEv8O9KwLrP2CAF/aoXIM1J40TbA5f
5HOwtYhEmbCAUOBYxLoJoY7bQzI/K0q1bX4cLj0AqpkQKLPEr+T1hkZqgv9+JZ+hezRknuhICEP5
rNGXC3Sq/O9rJvFhasZo8sDRPWu7QHbCcgEVlqC4a4Sbo1XUEZ9UdZ/HFNMn2L5aabt96W7IkIOP
V7TEuOWgN939wPUrF7Vmrk4+B9raSjJw00w9wnZSj+NmSUwDZ0O7Db8to4tAb3CkQZc+9pCcutfd
qlazk8+WmiATH5nvhlKZm/qo9b8vcFCfj43mEIX32p9MBCS3XolVn3a2f/4uJIf+8KJq4SyLuqwO
jxe0SjUxMQVAir9t7fyMuXdE62QlNpEUP7Eec2ASWLT3R8ernXEg6HIAMiLSDyBpHI1QtVRGFyXO
C6rXuHuIzeMpUntcGYNfajmseaJwfYf+gvYxTlfDwtLCN1LGy+QAJ0rejkt+ars2daWr7UkffnTy
INhlfTfu1iS/67HmmNsuJ/bPd3wK9rvl9bM4kzA4+WN2IbfgRWyMyBszpwFetsbqHKKPU1sL+wik
IuuBU8kmxmpvIvRH6aRiDFKZ9kSZ/PFxJM+wTHnRS6PBuDanUi4Z34R2e5dprftW+wK6v2IM3a+2
N4Z9Jou7C44oJcaND2s2yfpReix1w4Vv/M9hJ/IIsa2oUUwytzAkIYbt2CgPkTwhd6Dg8/noKSHA
LeBNH7eLDiPbAVDMqm6Itc8gtGbzCm67Ctx8Lfwta+XflsBodpj01qLCPEpPOM34lWhF3/eAdtZu
8ZF47eVKwn7EHIQLi6Yav4zKZyj3vmZrhTPjgHW0vRCqBL3V3koQCcqfUaJvK7gS4KLEcuY2eY7M
RLjfMK+qxZsiS4Vwuxl+5yvzdWgEEIq0cMK9ca9kwEfI2O4HyDfZu9BuNkrH6JIVYScsCCbS0+2e
YE0NTSVul5VXQ4BTZyeQmhCi04MPkn/L3oxznl1EV3JSGv1XbipQfNVd/k1FngPeJxgx+2hu4Zsg
LyfXDrLLYQL4PmSBJcz8uKlEomXGgfrbgMGP0/RK/2KQKF8zr8k1+gNaF+mADj/8nAEb29eGmccN
Etyt2YegHqIT8aqWwbD7HSCVopBZCOqZShMKZQBxg3AFZewpX3aDVC+g6oG9MjARXBIc8uZ3lrUI
meCCDoT9eAaQWbqa1ElsROOtM1BTLdbBywZTjb0T3bQWJeXlBVM8gFVdAi6D4vdpt/jW5UKov+Hc
c2FaHkvhqkVBZLnOm7exwE+cHdVeeMpRwmZ8gVwx/lXOU9SPARN2tWT1vZUCVDpY2yHnckOViCJu
DEJNBujsjC6PxQbj+7WqtUP8zsYAwBZa9xHe9iK+PnietRILayElXrnHJVJuBp7IhPCrRKrMCw3w
evXGg65EBjM9ZOdUehxyNVvCOUTgKv4ncdcmbIwhCd/kRe1tRL34M3gIcFFfG4drNhhGwxw5lJj/
zs8IxpdfCidkrDXMM4V6kiXvnWMe9Oe10Cq34z0UgOJ6OFEZRXegT30A20Effp7eV476FDHVBPVx
FxqchrdtkT5L0082FYpn/ezQgughhvCjugEOCwxgAXZbCh70lGpSIAEinEikVAY0/zoMsEj448vo
G4g85QxidTWB7DFkqNl5E8WsbYT0e316dfPAFCUhcxxvMCXa76UUtQscIsGd3SJ1xjV98j4Uxppt
6fPPQ+wi+JT3RpmQz2K69f04yQjzoZ8vKuuNyo4JFKKygpwSbK3Ou9kVyimFWU75bztf62eZz8n4
zzchumOJHKSogEA+42J4xN+TKR+kmuWHJCOkjUrhqtIyd+eLDyIQorRje4BQL0BIF+5yLg4z/vMj
SR9Ur3QkK6AbPWXIkqBQqX0HjUd5OhcbnZ7LIaUfRxD164i3tQwIyYVprYd6zF7e+F48sBKfUwwS
SiL0lWuK76qriEYWzvdkTB/35M7hmaKxtXvY2ftUEyuIP2qdqfGK7ZEbAbkOuKaJ7MWe4Rh6Kkiq
t2i/PmdqGHt2hYThDn0Dw6IcuGgEeQF4+YH/Q85YWrKGLujJiM07qe4mv1vRtvbatwOhiTbrPWlC
2u7ZqLJdiPR64KKDo0jtOKrkvD7hd8n7+QXAR0C3d/iXrlqpXij4vmM+SQl/skSej6j8yZ/5hTz5
uZXNxVAVIL9+6laM2z7fh4QGDMn6cQ0OK1oXHtqZsiDkkpfkr/WE1vPMCOX/wNDWbypkhasaLvYn
TbafsENRDD7j98etdLX5HYCpzoSorfQme7bkafjCPDI/PNAu8VK6rr+ci+D1OSM1bJ0fNpOztPiV
ZcZEXH8sOq+qlkJw2Q8y2UYiUdvYI03uvFTIULQczE+0qLm8g1z/k5OcPQ8Nb3XIUHiX7Ju8RVU2
CmYD64KA/jKQavbKh2sH6edmm5EwOFU93k4MxAzktEaomxe78bWSOK560XZ+98vIH7d6sDMfUXge
glnmF/y07CNWo6mu+PLVJFYpV0heToLkOta7yF7wVp062SQE7EvEveITsHp/VhuseaV0cHO9h8U0
Dw8W4GiZt25zdTovLmTj33mvdMNpqMlIIqTko8h2l2n0GNYxF2NULbzlZXua1xvs1BmwqTcqH88B
i0b04vFJ6WgoITqfEvv7rDpIKS77dqOTHwt7RTut7aWrwFvJ4vB+6lxnLBKfRWyYArVICfOpvlS7
Fq03VgjybKK79KYKqOcF2FIcHMVkCsnfYAhabNz2HCg2BlnBXMRKp/e9v/KKMWab8DLNGwHK10D5
xpsyc5/mkKIYdDBAnXqdGPTaPYT2ntAF6c8It6OeYcbO72sZymcfXhXky0t+knKgq/IcpNAho0PP
rczaXRDdydE5pylBk4CTc+wN9prByrtrw2apcdvOJhRFRtydyGo+cWy3wyzyvDZ3xsaLSoOOvVRv
0RruMDrkjhJyAhK7dif02/s4+uojctwpOxz/ZiBv0+fHXDQ+hDz6U1V+pxjY1Y371U/88/qRx0KS
qcUMwgh9e0nI9O4jTL2YxK1OvNb/JyCZftcAvKkkhul9sgqFPtNs7s6ZGDxjhDODVeche+F2AbRj
dB+2/kLwXrJY7k4i2qum43sA9TlFfFivn8JbjR0HeZKEmJmLF3+v/s3dNqRy/Cmfbzu2CUgexUds
ooDmpQ8OiqlmgEFTqiUpFwtNv6wF03zs84f9hHC1UTYcma8jTNa61DXtiMRLOE1FicXKE1uNqJh0
keKxfGvENt714dPI7lsW8dWJn61xXk8tsb+loRK3xS2NQYrAgea77OZYCfnVr1L56GWSlNnUGz+g
T4Gw3fJkg50H7exqgWprXCUsYaMUhBvZTaKQKSx7fL7tZqRSKT7R25GQiiMHB0aDBi3zEQEb7kKe
9vnvaU4y2/qjh4SU3xF9yPVXGYDOY2/oWrpCibeWyyNV+7p5EEiqW+w1c41CCDQFFbG24QfHLI96
4fkTvUWqq/Mg1LaV7CpObLOsY/9MdSyjXiduREkbtUr2LL8nWT3XEJZd+aVAC0DBD9ZVEwThtLcE
o65qA+UdpSC7PPIos7+EnO9WfVvsCEdATcy7L8g5p/YyNxy7wRxJ6DQiJ0WIby9tSNzk0G3IYZXQ
dvHWVH4kFJa3RizVCd2FDwxcpq7peE125LNJ9DuhIZ9wlWyj89cjnK1t167GFKebtYoZxlPxicX7
kwXOfpKxDji8nh9g76MMTsH6xz9uvoN++CV2Y+qBKdu3AjkmB6GkaeCNkcq5HeD9PAM4hBoq59bY
/3BrGyj5WNTnlfosirNNmEYTTBARdsDFy41HGoJgmRinB/EDnLtzVKUwp1omzoAQalymKzGGIP0+
jZFtecqZI+C4Jp2yD/Byvi6/v9u6Z77Ne8FE32v44JwXwKRUY9aYYkPBdskgO+S0+LULbprbyiJf
mYyfGFYlLhTwr8l51GmOWlNMKtcWSTW7BzfJ2udd9smO0SFU96oM3lmqlo8uf5bMxL0twKEe64Kh
xZ7n/KV4CNxgVd5Cvc1Th8UCB+9aBFC2m4VvU8S+tz8j3HAD0461HLTDZhyYGxDd1gcQgMOeFgt0
p+UmMhETj3aUIqRMb+UuGh+73O9agNuPA9/mNzjFrILkmkGEoicBQ9gMcFI816Xjsn57tDOTfXG1
0gSrswZzJglnFFYb0oGMtBWBGQspl4N1dIEEPn13bywQ8SuPAM0221Tb8ypwApsHkevO8sB/nEB8
zeozKH7nPGdGOT+A5ajCPxbqRv420dMjilJLjSBvj0KPZcPEvPp0PrfJRH4sE737MLheytuCcLhk
jckRzYvSQp10w6GE2CkW+ZhBUa6rPhGS6crAxiU2+aFQIg05LXH0w+uYDiqK8jH6RsKhrbRKnWJm
0nOTxAHNvwJJBRgy4cCl1PD9XjYWhyA92PqzMuemhbVWdnVmA/7rN7V3gZdBk7+Js6Qgl4ka5/Uc
OG3q+l1Hl+09fl+DQboiSNDOFSh2S1TOjOQYatcGRa1tnsixgZJvxl71DdSdCkJ1VzzxIsio85rj
9KssV2NXYbMNC01M5Bx7jtdKFLul7y/4D7b27r/XN504owpPuemownekjOSALCPVrcICbg3FwSCw
dgVlBEIpIB0Xwp6AJ018rpCwQpl3C/a5VVlALmSappJfLYgfHBYO5jSW3TpqclySvSv1+IPYaM16
vXKBtdgpVpUPQ+/cokbwrvp5YZmYM+XWhn8fOvsvVZQGQVUE9NlyZ+x175bPSE/LtxKMGUQB16rS
ZVKhiXByN/5Ojaso/J5i/ns1nTER6nvOQ4hLU/PwYdh/0i/e7fU2TPHH3s9Z03jRVglxboc6+ro8
a8QbjQebv4OmmzTtGHA0NrGxkTRs/x+0A/sANj+lxtRX384a86CSEEm7P4QkxdJH+cjRL8M/G/f4
bG/LOYdVtdNMko03aRBB0QokDCby1/oeh6Xiu0uPpzztlybsHnAs6kxCytrFS9OJCfO+NfgxknlR
uxL3gEgrAWUrk+Qhe7AltbAA13QNtd2cUVhRNMp4BhjxdNm8CFDnYpnYa8/AQulg6PGc1kQhlJLH
yDXQpMnynhf3izntfy2Nld4nwpZCj6KXuek5AKNQJbJT73wbrR8BbJ+iIYkVfhw/pT4GA6cYKIkI
cbCF6VMYfBI1oc7NWVJbtWkhwZnhHwVnk7D32/euq3ffSTpA78Yjud724Qpg56fXizwPxtS/PCv6
NqH18gS5PqBhZWgnj/SIE8y8fh2w8pOJM/jwt8qc+mrzBWkrNHkGak4N7FW+GzKkNZndvOjO2LhW
LTSs0otEk11xF9jo1lfBSBINcvyaLeZA5G3AswjP2KGCayPbjMlyi7lX5a7+5Q34Swjsa8WVNTpv
Ojo8T4GjE/qSBFJZYPnawLcUx/RD4Uyn9zuIZ1JzYF4Xj9hEbOrEKaARA2Qc+56ZQCsEGvN9F441
8OhkW7FB4oGFQqIslIsLmIyPEpf1d9KM93we0bw5Rxlk2RRyqdaGWjU2Wm2CwLq7kGLXGsWslA/x
g+qbcAuN+9rSpazij25r5XSchn0xh1Ympz4kJMMt8Z4woyTaDhclOsR6v4MOE/4Tw/dtNBMQhFWA
74XdOwOn0MnadqQp4HwzLt9567E6zedKghxYfiOG0Xr+TxtmjBcShLW4c6hBpjrCVykP3an/jmlG
CsR/Xnl9qLfYVHeFYUQdT+NYWzNaD/MrHhbJwj6i/Qv54nHDEZLLjX5ibSNhTuWQ/uktLfC/3hkV
UlbPmIeuxvTkcarhdpgnOWXJMi1Gqzklrc+54Jswyr0+zLdI3K8+/PgA6xwDiG3BQkTzTmbttXTe
1nHfMvMkIlusSebKTV3x1cdoN44zl36Siho3O4QXspZYP7N/4k89QOCoG5kjA686usLsieFoKemo
JQGdAXvbTXuwp91h1AIKa+4maShTNgEoV7VNgkkscQ7YX8DqyE8JP5SYNA3FOw0QhM/ARgiBFDag
QYVLwGeU7FU8FNmd1/qen0HlUU4rKSy6FsVO4qjfPDsKOOCGKzetZkqm3U1HknU5ZsF3pcJb8XF3
3kpGi6r1+8M2lie9ZZYvVH0D96c2YaRwOBqRuPdJQvJ/w83zvjxj6MJ/6KFDcvEL8vIqze56lfuR
gpODio68D06m/QrJ3XjkULVED6MuvnzsQHq8Sg+IoLu/g+d14YkVvjn4Aej08DVWzREGOw8nzRhu
VbgZU/Z7ZstxjsIbGFuURueUmH6ahGwalirntj/731f6Y+4Pdh8p7c8Uq9OC9H1VfjmKSSe3Qhfo
x3pMuIohXFug6BYKGRHoQxzjeWwOz+HaA0C3jkpEPSohcMkNZWGjjNEiIYYamDbfRGRv92scXJhc
Vk/pmbCYLS00Fq1jIfRa1LaVeCpPS0QqDIJ/UumuyWZECegmTgFsCrIOGh0BkcUwu3jgg89wOfcJ
xwISAzgbai9b2/xX+Bl+4fkWij0ytNVN3zGPqw3ufwZ09MkAZx06v/KgXvcbBlg+SUI925SRY7C+
hZE0FJuNgC+RXgaw9M/jepX2L9LdlazCjrYPFTfk20yQSzH39kE4PoqOgRvuAOgi+3Ae6RL3/LiE
I/QU/+x4CzCtX03wU5xf58CAMe30qO17xX36EH9hE7DuflgiBF44OoZM2aUu0tCMcGOQ3/WXvWJF
2iWYEMIG7msEVozJ5zacWS2A1gmNz/OktKJ/n6gIdtMrxxW7Hj/v8qn13fyyCX60Q4ZaGDoJVNkw
BfyQRtVxrLMrNHqIR4SHqaTy8tAeXYLek4ZS1nOf75T8LDiPEfDviUvqUE1AuFoMBqWXLXODzt3X
wMVC58b9Nf3vemf560pVRdA7TO1EfJQG8d/Vuptb8kmRoN+FQ5l6NyzKkXtKcyBaz+GJgxv6UaXI
+UqKFKfkhc+CnaZKQM6wz6gJO7ye0snbDjNsfc2E88nemQYpYp4ndLF/hy+vYgWAugjOQ4drff4s
tpt/p+MMjcxp/w31j6BDPJ2EsRcsIHnqMQpLfUUYzjOOzxcHJ6Ekp6avQl2ksmc84PVe2c+iPtkc
pJyHPiiRlicakLmNsNk8mmQzQa2kjkzHR+jPt5AF4P5/K7eSOnh+dICTtBpNlzDsmmxIHervMT+Q
sj+al8ZKpskS3WCjx7SAWDuCOb1KFbuQzVGWUfZYOWnu9/D2T2SZzWh2pyt/6HWbKRub4pwOl29P
2mgxTyBS6rRRocZ0A77wWH0xDs2eGO5RhSzqAzENUcffKxPThBSLdttOyUqc6o0sVffBGei8XjHV
tuR7vQVquGTsBdL9yZxW3Tm6cAqesR9sEPn+P9FZwasCUVBLhlTvsWYvK6SDBsVSzxztWEq/NwKz
skGDxqgh6lMt6jCLs4WlhzSldzJULo253FsXHwA2gL4Ub6MeWXQqXmGQCwymFaiSbld4w1bPiq+T
MJxJoVVK+/k0O6N3smxr316f8tnQed0azmrlghczWTnCq+HBy4cvLWChvJ8K78M/lLRQCiZzF0N3
kdHXzVszxN2uaW1CxqDfooosENBzGYUfzyTjhqiXwTtcuty7LCXZNqWt/EgIFpu517iBTC0J5+ze
f/RF1J9SxLWCDl05uuGt0Pw8CV6EpHmF+Iufeye23n++iSB0XZKz8C6sv8RhTPhiQifDbz11S5bk
3SaZqH6MWnmA1ZH7Qrqh/nbJlA53rQN8B7+R/nt2JlzMJbuvZdwopyeQuLhnSFY189sGxG47szog
gbjm46s/zVnrwnbuYy/8xIsnJAnfHiNjmvfrCqTbtNxRbVajVd0152kCDKlcdvwEWiv9O2hpF+6d
bmbB227pI7k445+0Tw+XYVBC3JJReCFkb6zj94R/mmAUlxCVAOlshR+CRq9/gfsJFGE8/CH1UXXm
bfegp5im0CqXiabHZJC+3Z1heLvq34ouSL1YLbemG/4UFh/bTyWiTn9jPceqJHdCi8rcZuxaBQGZ
bfAqJ86CNl/VuLJXgTGSzyjxa45b6g746qfmb4o3PWGX1Jq0ilufOq/Uy0jtHbfG9ESZBcbdGRJb
Tn3xU/UYzCV1MD305rLli+E/2+QmIHPxpO1GvJCDOvvyPA7QI/MRJnlendCaIcEEd5iLInAuRv6A
O+LKu8SJN/MvkQXkIg/k0aw0Wdqw6JF/1VqVGoAbU9xy6ekaw6iws/ho/xCCL0Rd1jXyAbo3rntI
YHzurEulj0FG+RFAuJRmwWJk6eiR1rHxZ8O+o3s/816o6jjV80OUIS0n1JJMEaG7JpbOsCTe13BM
4EQzXdSSgqVdjqhZoh5UH0ARKliPkZsKqlDmRxu7GErZ5oOZSh43JyykXiKPcW9yTTw0A7V8L8MZ
Gr9DvQ0cKpmRG6FoAxy1rl2vdiMELRQ2OYayk4c5ohsjS9pnKp1Re/Df3yVLauz0mvqQFXQduyMw
wuZlqInZzZPs+Qz2YHJjniS50CoiXj34GMhYz/Glo9TC23ehxx1AH2ej/sZe4F7+cNnRbWrh1N/F
xEjJk3pZgvSKenlwrEAa/+fgpwLZhAJe0PHOAwh/VMdxpbdNnG7wC4o3MR0TF9n441EI452GWt9s
k2PWsB2nEymKvTRTVfryrr0KwxsieFt9KP6vBkvQgyT4+AR+dBVD7X8CSIsdf75KuVThdojk77c7
Ai6hePbSEQUHUpra32AxoH06reYaxSGT8jdly6gjaQwCSkJ2RLcTNSS97zPkGsiQPd/TgaP3imwz
b+k+63cLAODq+brmNKlNs1/qGQRAUAB+QVdNeXFYnuddOr1Wg9QFi0lk5iHWSdA4ahlcemF/dkWY
UrfYX2Avv2yHsFWU3xy+foSt7rPS2EifvEPxgkEC9Q/xu9KcLmbtwqPunEQDjkfm2d4F6FGcHvew
aVdO7wWAlhIINORYZdZV09EIOdDjihkaqkwPyyJkyhWLMNqSWJa84Hk0F/QmRW4gEaZ3+6xbXFDR
LDKAAwvzN7QVQJKPy1NS9T3lNTzvCtht2SzYo9tVwrr4BiaJRrwK8W9RsN7GxJw7VqwpAbJShavR
GAP2N+R0VWtkq3eOjcWJorkqKjConcaUm4WemHKgdwIO8Ux7/11o3DBe9JAyZsv5gmQ05V4yVPl4
+2A2TOUe+qxpS9rf/gIe46dvyBVO5jJ8XmBoAvzOZ9lu71yqFVmXLyMNt06wv8Ho24oDHkM9kLds
9uSuivo6bPJF1etpxn2oeNjCB1eJ6qjT+Y5qyexCKqEXndVySo/zjZeXX9hlJX+E+FG7mkKeuZkW
mTgjg+ardsBsTEybEUYThFlCuB5One0lq38F8Wb9rudyhNJSy98HdnDC6YtrmXS0BSe2AuB13Wv7
RabfA5+WGdpYxOI5msf5WL1EgmNcdU0TrTT0eEkksIPr3jX7vMiWEIoafIMzgVZEk/bbHyxUuQ1b
1cc/7fyyRiarl4phc0YwjdedLhEZDWAndqspufhpqak3TwS3Mkq29XQqxg+mkT7D6tx0ZkwaSmLw
OY3kbh6xiBpOh4vp2tpjLztdtEsN7xG8wOGfxDR/iTnGLG5aGT0q93kUdbk3o90O+2uj53WZibrV
wH4YL/OmezAg2neBfkEfKEWVh+wOhVM48HVJgLmrbUkuyBI/LUX4nszuQ8volKpZCLAX6Jfrvq3X
EAc1VvbIxJ+kR7R2a3PHJsUo8JRlPpRpO+xCEQZXut2nppF2TzARoEl48XqhlyTCBXyZLh2/z3+o
d+oxKrxiPaKTYv/Hhy1AOOBo8qfEbDyiAZ0WA3uJaQsQgDZhenruEb0iWYpK+xAcU3sGZxpbL8Id
RuidE7SCxSkRTmJWAUCtvG1kfuiboBsUhaxWggP5Bn607IHIihIvoD/2KuSq8IENit2DnJlQKIF4
jqk56iSJZ94BrgCrp2HeYhTZqJtmx+QAWMJv+fBaUKNqbLPSBSz1injjht06aSKvPdeRcu1sz4uO
1sDiHSz/GQCxaf6RM6l2EuR4pvaX4us1Ngb273QhBHs28iDQmwjwy7grIUYRSuPrRyEoGP/drIDW
//7kiHYUHMMqO8CqOkKZWdguB2VkI2WbIwO/BykppB0gIcO4k7fPH+2hJtDQcP0s8vY8t3BsgGiR
RuhVVH89UF392RU8zuj/j0XpoxTF865yxu9kJir4oDfomYJ4/ynacDyXe+FhuN1B0g9OuDvfU7nx
z1oXPASCplbRX4LJ+UaVqxSZtBwblE7eakuIN6eeA5cgmwP6D719VSHyUAMo65J4c963Wskly4EX
PB3QiLy13FuCgw+rOlFFKCtyNKoHoa29iO2lg1oiI9e0CfTa3JIx1XvR1pxpnvx9EaVA0hTJwzYw
QHUhLvaWZjXJx7HcX9LsGGAczqvAhs5OXrm/xd9+zgyb1lXxE+6TNjnoXmoLrfNvmzxAlxA8sT3g
7oqOn59euSdG2nQBITFj697cB++wxPhP9wo5FfN/UuJy7ps7W/eShFkMTs8Cl/U0OTXyH4996sHF
gxCInFPcek6V+bp81RSgnCP83xBZNJlQHKSpn2AG73QizHSElZOIOPm+qn9KEo0EabUAjeTrKBvJ
pXlKnBEnMKm7/H5GTifVg9ShXzvOv45De7I2BDADeVaQvz01StxIPCQy40D71tHguKh+b8sUEQdt
bOa+XCV8Oi0UuOScmKhK2zGBmJxtrCD1tCAfXXJDMprfWk9eu/3LkJ2zFhsJPIkTJpl/phQCw8am
Q0gXDMcabBTLxMyHMD/Mb1p8dSNGZu9HhnIwYFsUzzIm6WL2Sdy8I08/dPWFRhZ7xrA9TUpAIb9d
nbIf9z3yO8pjDYgcCnDm7k1EIZDuoIEjy8LIrnOMBKVfWz6DiwnyDCWTtTzy2lKVLNRjOjYyADKd
Rt8sweM28EvvtrGwCftY3YbGpnF279QcFkJyHWTBXEtY7YN8PsKdxgozaZgPxVwUYGkSEP9FGXTW
AnF/TG9M4hGoD8u9OwnRASNA773WcxvDvoYQ+A+NCF9g8KXqkS0611FZOA/2op7c9neg3cOgAXJ2
gOS7CrHCef69X2C/fu0v4t5s2Wc9naaK7ArkUE3TPvkJgcv4VSV87lCpKqN2VbzfZHJjwwktWqYZ
cAzf68z+2dS62cRHjL/FGkgjrYlF4wCmy9cisuQTOfMt0izoRjKU6sfoXLFal7Wa9G5rrkQ/3adg
Sb/9jkllBnzuUnN71VlYfJOIl5pfu2LqFYdWPCQvGWs2xSBVHLrUnYdI5oxOPU9bHLn3rQ6HaKjO
fSGpFF8C1I44fPGKOLTqZzUm6oOvysuYvPSg6UKKD8NfK6YjqOr3ZruA+uq1FESG+6ynYAj/HJJL
A1Jv/odGwmfT24Ek+PCCLcMF7B2Humwcem75XeKMzCEs4hVuMRxNm2IOVE6TEskH/kLnIxSVxUKM
GslcEbNXX0hClUXqAL/78X4RRqIuvk3KVpSIxQVoFqlKDuUl1mi5jRaCZDVzeTz6UM/VBnJ5L01a
92dcO2ahWUM7mk9Pcl/nQ4jhn8riIyAPp9IP2kdlIzdbmvLyJWk8DQZYxbJm7WjFFOpdNGJJQboY
MSmbhZQdYw+Pcg7l9Vy2MZBcFtR34WzMUrFTyAJAbn98ONwNb/cu6gasvK1LKBI8XbjTF21GPeLT
JnPGp5+F9reKl1qUqoSCR3/TgGDUyQ3Hnb5ahUTDKTRCp12pMJrVDlQvfLQIHWSO4TGgGlNzXyJY
LrgGoa2hUJrPR7j94BsuVFbHX7pujvEtRdM/g3zjYhLdT+vWRJ2b+7mjAbpALrwCibOVHCkf1qJv
3JC8B90MFDuOhpQspgWl1b1ijt6ZvVwaAVyHxf9mdh0h8LxmKVtMH/rwntSHRK+KQG9TZBN8x8EL
gCSN+6Qb2VDhNAlg0OJtmhzhpIgnCpRwvlS4AApJk1vRGXib8+p38igXoHJvRzNupHHIFQParGjb
Zg7uYPMVCwkE72aDOIDent6Bi8Zf9XMeD7Q1KqDHxVfPTKjo29Uo6IMC+OeKCbQs6plSVDVmcnaZ
dT0K4GD3zd30AbOdlzeIntlg8d9BPhy+urt5ao3RjGmOGVLn5NqAZNkcOI42a/tr8WnO54u77dCM
+BSnS+mRTSOU6oZUS0GEMXIcaYfVDnlMvfaCX8rOlmOkV7g44wfwLp2ys4IoFNb7Vi92/tfs0/3A
SO/2QxnbRqNJ1ZvMRF5kJIHuesYu5umsN2UJyKIA7eeW5pAImDvcTOm6JZYjAslPbpWCCL8kfLGP
vUGySkGROCR8LJUJdg9vQzNBDQC0l6fTk2PnFSz7M505AG1RDlfgS+zSPsH8q58qjGlCVyt9Sd2D
YYYOOUmqPt8oIIXh0fhmlrAnPOJVSl2wu8K3FsjCONer8aaFe4i+4NgqlqkpdvXh7OSiiDidjR8D
H5JKqJzSiBjcLFVPLu578xjf0gchU941RsPJloNOGrv514KXYUsSN3m5dvMOAPelM0/Mlim01Lcp
BRuu2tmALzjyhnoZ+iKMX72XbukbO7wiAux0ldVOmvnJ9Mm4LXtbXgju24Ms5GnWPT/XUxRufmHV
Nx6YOPWByiCnmDIFHM8hwAd7nnkgox5aNrKim5pJEEERTyaGEvRPOyTE76zpw9hDRQwSLogB2rrM
kBKV9RUMjAM+AcqTtIBp0Muv7R4QxejjegObvnpBLrMmxTsKumxDD1qdOelXpmGTDUXZp0CUc4tj
xpxizqzmyK3JMCf/+Cz60dlDMoSWZcAG+to8oHZhFH86jcOeiY/MAPPpRcEyTx6ofx6nqHJI1qLs
Qx1pL3pmU1hntwH0JYBYBlaTFmWTnPF8s/w1eAbcfDmm1/VyYdTi+/AxHZhOWVfAARmIyuUNXgi9
RR4BS+F/0lW/qdoGb9kYIBuFL8JLcwcyANV0eENFIcdynSTgjWxBDBioVjlNMJMoLP9L5uvEMEYc
adgJnPiyLbx1UVohuFh9pZEQB5QI1BLt0D7HTpyR6hSoI3UOe3J8m5szapqV21EJ+ySjlT+n4+T6
SldDAAvwRj9nKtQXsHlkgGThfY3AhaHKJPUk6IC81vnxW4UJ9F8CAunqHKPfigwWY6MZJx7DF+Jn
B3n2229pwlXxicQWfi0bV29jlBIkGmjH1VAExNKwRCA7ZmU5XJRYO1Y0yS+L1I4aZJiICPPeudVO
iSCxziNoRlm15gpmZYkx2RfJPfZaQBPLZmqsqkz9McOAQcJZ/TUlIEEKcXsPsrU/Evz6grtX2tig
b1vLdjt52FaaVJdaCX7vIcMGH75IQgdDLrA4yd1qVxXNZR82pUthXbviT7NbFZ0M4hrLbhHcPVI9
q3h1M1SVw2m3vlaPo4woX8/eYKoXGugjT1jIXEWMcz6mcLyhiVOjLY31EPFMfs9KPD6MtqxQm0dD
owL/D8GEUnniK3bc9Y4z1TNxmdtNE3FzXHWnuYqR0KoFddbd2tQSffLrWW2fm3Idw2M9Jun8HRUF
YLEJCSvYuMm5i3onLREqVH045CY7f5ZAcgcwpUZnEOxidZFmvrff1B2G2thR4ehBsV6FL7Zb9CGk
PH9+3+xLCViINGACOwu5fCJunYSvdJWx3RfxqS1+kXJOPTtU4AAVuNJ52xE8WX55qTmEkEAPh50Q
E5ftv7Dpl2GlrVE/fumFt+iUHy373cRzd4w/rRcEqhsGq243+OKn3TJ2pVNyfMyUFtksjgYDqARX
FIvVmGSQV5tqXZIRYoWuGyH78u4DKCu2Fc/BGuK17oqnv262wMWoTYnNuN80JXL/SzaMqIk0+DT1
mJjUBZbAQ+y9wKCCRxTPswtS1YipIB6lHYTPFFuM6gjI29Jx+4elnxLULtg0dRkW4dIjQ3OAUNzx
cncXs1S3XCbXqpsyFNZC85aj2u/Hf2bCvDWUIE9203qyAObmd+1OspZslq2Wkf2JnnLLfjHfL0Q3
beuS+jZavTgqvcAujoPx0+hPMeq6Vi+c+nZSpkSmVkXmG0Lq+QZWM+SxhrglQw5sVGJ7mRP20wxl
AuyEctJ8Z/x/eaUgduNIG/YWVHdtRFEQuNlc+bkei69zvd5dJJcRMpsJ1LEixixaLHX3gP7mp7ow
ZfoJPW1CdU0ErHGhpU9Y89gESO+X1XbiiQi0rrXzrsi/xtE9TUaAb98sfwr9kqjY/Inrg31GCZl2
4qFat5ITq1X2AjODFma0AIWBaxl6poqNMVICvTy4KzWCjfxtGI/NWANwgFVSESzx5N9R9Tcqnoiv
ukD+KJe//Uce+4YSNMSFy7n1o1s22EcR/s2Hgg54joIZrqP5xLQ2dXeD1aa6FAcfHBfCoY9FqA7e
fYAp/nTJtcBaW8Tgyec7vEWHmY0pRXEY/BBJl/Xb/XjCFZBkhxBbuhgfe7xCWnjU2d+AfwFO3ZiB
wLylW/jdZDLii9kuKQ9GwWsPGGpVmyYSMIHDJkte0d0FDhqO+O6+2gPXNsuYbGlKSPZWW/cMkM4p
uDMZJqfMrPbkbWjqHahJMRS/xkLRqRWeI2eKIzWDHK7JdUnqAn/T9kkXmZ5L4i1M2WhZ2ps3xPyQ
CKxJ6rEKlOD94UynekGAgo4wO4u7yr8XS4c3gDsgMEqQn91iuqVwuU2AyIRDBjLNO8r6HF/dP8bA
icF9cR5McLRfZ0F+U9rOEF3J6jRfzgjkGG/z9fK7WIVRpM0NXl6utOfm8/oF//4O2AJnW7kv3YGM
t5VCpDHxh3KEMeZxrSG/mfOlICh8SVjJosd7iYGz749ROrUp6g7ssZ1ynN8gSpmCJwK+KCfje0B4
874HCpq097WZ/BkIAuiLD/iWmWLPwgtl8lxem8jPLbJqCJnbjTd1q4Md7D1+aqCPuMuO8btGiuAJ
q5Y2grf+LgCzLbpK8qV6KWjD/wI7BMNj2kR8ay2qmP/DgSzoxoAamOBJbZGGfoAqNfqeen50KKNk
pC9APvLSLfMD1KpenS1yJRNRk9WSGo5pJGaUbsl5Pl9Hv200cYliM1dqlK0sNZStovLod/JtzkI3
Bx9nO68IczxYBHLIYgNUk6Aod3Or0JzNJAH870S08wGAAomL5CG0Jtgz2Jj+gewgune9/U54IO6H
c0YKWYcZcxJjyQMHrImN91B6zkHFfGdA0sFxB+ZOfhiOV5pxSnu2qpKyR9+xdZkEUpXJU1AkAMY/
SclAbA8w5ol2CJt5iiQTdW3+PiiZITupZ1vYKcGhfe2zvExyc9kVsaOG9ypAV7+WhRdG1nMeHbwd
vcD5V0xC2RNUHaCsbalnQdp4GmNkNYZ4flcmstrOc6qZd65itn2k4XtJmUU8+AeNEc5ydmFM8BCa
yulVaRlifxwOTu03qINkBXrHgX9dmVg3CZVRmrZSKZ7f70eVnKtCNfZmZ5UF8REzDUSVgsChORmN
emTbuEYXBYRFaLOMGIU06t4VNPK5YoXSOAljdwNilouRSKTTGkfb51287LJVun67Vs6NZ952buSu
WgcBCbql8Da9FX/HNimLp6+6q3ilY1luF4SRGBNAjUoT8Tys1RZ5cySvcvuvs7Bf3Ty0dhEwM3wn
BbCP+twgoLS+jq+JKBghzUHXSVWJULDDrfKJfFetyWiC3Fv90cLJ0O23UZ0hA2Sf3cHa6GvEgE20
6jKUaUll1QfgDCeQhX6N9xUHM9/mscFiQDxid6/2EvxP4eoo2xc6I1oVb5ZkXEEWKEC9IHRKf+ia
AI6KIdD4CMrpiFmRbFkxsqkt89LyGVfiY6qQVZlw1bsTWCan06DkH8NkcMa7nSu8Yfk0MV+TD9o9
DRdu3Vcu7ITTTNUkrjzfI2+ddhyq6l/rdHH2Bp34fzId78Zjp1ZNIS4to0rcSROD8ycgGu4czVId
vPwgg0+79gKRDxi8K9CpGZraoQrkXN5tqU6o2bQKk/VBKYXZpdOLWOFCj1MkmY/q4J6VY+xZYhls
GV9lXFejet/ElpD/CHeq6Q4aRhFQn2MDnkuTy3D+16CrOoFr1QYldF6jbQcRsvau+eu4XZlQmqbl
q0kIf88bO8K43kZ1NQ7/0rs+vlQKASEE8qPPfBlu5nL57P0Ga+HSdo8H3pPEmPUlWIyKm7U8RIE7
8qIygxAIB0/6DYl0s12RKYQ2zpoxVXg8WlzREpOuL7+McgytsrGV663t2+NlnvImWDCTlDmCRSf9
WZ6gIWvTG5CA59+1+CEeamjNTVHsoF/Kt7dMm39gEO4PTI2y8kXYUhWodGidpYq2yl1rqbrenRZ6
t6Cd9mQF/O3e8Ta2a1WQVo4o/+OPmj0UKVKITfYJkjA69JAQw5e3p67V5GRjgppAMPUpO6ncMoKM
UogvnpVV6aUPFMZvu3zhk5vQPMOi22EMzxUm2XI9h9vESoYsL+mb+2iVk+Kl3UTgSH27x4077vYp
jo9Dx+jJNzcc2WmNqxH7KU/RbFCOZ1ykhuyoPmcQSfvnUNFX+x7/xVOSmPCeGmaeGm2OOAPYJRI/
n739mZOxSOb4Ims3gc4D69X3FXSzmmUG7jfvWd/9Fd0dj9GBTc8+TB3TFiPQLNKSZxsZi/nIz1pO
UeZJt24iLS5TzuRleO1dtfkYpMsQoI+Rry3di8LD0bfLQWVGoZ4heVGSh3wDEdsjesuv8wH0fbev
gcpuEWs8ghFC1sku9sqfKq5NBMTOFdy5DW9B9gheZ55iJne3+Dt/iBmWsRoXujBifsvvhAOjsxi8
BrVNWPzvtZD7cDrAb3+V6Qtz0IRLRzuKqG/Xl5+Lvuhkr7WtcLwhzoJJAVMhiPM8CkfU32J7badq
iR/Vdg3DAeYgf8ipWucwlWN59Gt4bBqeGIGUf8aLTBTsQsyhr+i12WNJyQVOdpHlrvgdcI7EsOBy
MdN8U2ktTLss6bhszeP05M06apyxKX0wZmfK4PU2pqhPuPhy1+tlYyzVBwPZ7etAfwwIsrrpk4lF
vwEzfcECtxUMsBdpAahVC3UMWqZSQtTiEjt4fObwJmBTBi4H6qGYbtAd1A+6THaUX4j9S1CZ1o1f
zPfm7h47gg54tBTOIMutDrHNWl383SaTTLPmFnX2avYnoJeX8IjDjLO9uflzFjs8iz6PdCfjW/oq
/W7ghgpsIQebxaAnLDO7GlI5HDFv6oI8SIxbZQVuR+ujBijDQHlc4TBsKpaAcVq+aRZkXCOvL8o9
TprtQ9shq8H83iT0/FCaBmVO6Re6kXuqo73bxz2RisQrg34achCoYGXHbwbE93OI72FvWEkRYNCO
gosbD/Oy1bZCJIwj/Xm3doTw2IPUjbrhW5VOJ5Q5+Rw1WT7wrjPBlWci1DF3NaP+D6bcpA71HWeH
hmVmRMnKWPpFPXrYQmh9lwrlWQT2/niYeuq+MCCmxDYiLSXfpIAm4Ya6fZ6k9jj6c8g6GHLaxIzM
bN/LhGkalwjGC7HeBOWh8kyaeqH1ucl8flOxGqoBRCa3k0jeDE90XMxi0bHeFetYBI4lCsSWZOvB
PidrnC99XvMdvnnqCl83iLLvAqm0eNufNpzn6rXvS2O6ML4fc4TDgCC+FJvf9mnfwySJzDt7j9ps
Q9u4XKFbjbjrZDnSIBal2kmJJxIphxj2ZNoT5Rar2KPMAliWLnQtShUCuJ9tc7vMiItmg1LoyMQJ
JRF222V3+rjZM/NX2FceKRwkHCTC6+EkomGilf0yPRabjldmEi/NamOZOvp/kZrmwltGaQad1mUy
lvCqunsDw/h9JuDDcjiewYE6jdKV4eNDLeAZxr3aMuyrrbN6Z+qJk1gC8G8r0TfI260QykN6m1bl
bg2zvVpjNDfzHkKPvAxOo7P93bGt6hzRK92pHVIdYf9Zm9GSXtCspYJNtwXk8vvLFO6F7uzqyDcB
RZCFGC17MVeph3CqrbNXaX0FbWg+qDsRiwGBRDh4y+LM1T9dMluMzZFSCl6Y5sJgFylE6zZHSddH
1J3kDIkYiBxkEWw9Mkcd0WBaosCqVJJiJ3Nnoh1RtxW83AniWVUkhYKy65ULm7h2zPyTxVR2LsEN
rxYmMFCr9ZgQ457XNAu81F8owPFPNxHzeJeEOlZi2dhJD8OB6rfLtUokBNmXAVUWyTUSuhVw2hfi
wi1C50wmu320B7jkCBtpxGQKbKr0seWc3djN+ql0AzsWLqG5d0lcnGGonTb/SPUhn/AChZiwojPy
XNA6Sp65pL4iw13S0ClTuMykoituMMt80Uw784TfKG2iqCGOaZk/waoARyf3U8VlFJufSz17QHe0
W5oSSEXbsccYpAIfalRq3oDacuBnB/LpKUxoLEhx7a6wJvCC8aGRNk6r+Zs7zgw30QUiT9QMQfbI
WWZ4tAEmehB4OD3es1rml2BEEbmq6NEM4qxpPrHxL+43zwOLQRjttNPV6TCn4IapYorxm/HutQly
0RrhJuOe5XXini7bpj2D0ZT4wVsx3lOIsbOuhor3Mdr668BX2YhNTDLXyYymrxkKxAo+SsfDLVtW
OhkDwHMnfY+RM+bAxuCiaYPxteYqF6+teu6wTVRgT3jsy20a2Da7QJO65tbcUrdlvf/u35muXK0C
NVk1lINwLY9l2R55+oss7Jrnyzjyz1Jn5OlBER0IXUUTGZ6TLawrT4iz7EmN+3grvObys4dju5FS
Iip9/kf44a3ZWYaTZ9AIhyZ9E6W6khL/90JuHOqiGVx1frjfBkS8Z0+eEqIiEGtqmJAKaO9yYcnn
wgMc4POlpPfzajh85T1uZ47IUZJZWEbpeIGwmtJVPvCusG/XGFiv8Zqk7//s8p96emgsbe2JuvQN
rPgRcXFFT4AcuZGnHqOehsD5W6kiiL9XAo+7MVX2DcnSDDEGtqLuyEYhpDTJc9IJv4IZ2v+lel7Q
0byBE+rAHY3hxAgWGBj2Q5uyEAH2ViXyVj6A8uaZtUxYxutP5ehjXBDm7nOMdlrB+H/W5Af+KNoz
2iqOPe8xtGGSv8tLfsN1cOmI4erm6IJYmaTa7K4tUm6+goT7fgm/XUajTUbVri3NlPGTFHlkNdJu
gcDz/UM6r0IM33FQrwRR1595sZWkKMwTnHCBu3d7jsf38CyU3E3RtJi7+wgaf4lAuZxc3mdZmAgl
NtJvBTVlk+DdCxT9uXs6+xZi+Zu8o82vpe9wtJhJCOP3qFOtb6G5PxnilcBvQubCRXkXaX0IuPy7
5fE1JZSYeaSx8iuAhRhTFpDPOJ7C0AifFk8J8odqUtNc4iSwc8cGqmKmAZr9icc04aSnV957NVZr
S2tOySPBXe7CbTJyJ3DNUVYzKk2XQnUvzG07yWHHGyHq4RnMCiDUtFpJYoLMw0MX00AhowDDz1Pz
fSijz29Ln6Az3KqQP1QUQwV9R/sfmPWyXtd/lHetvAyuMaRnutAa6BLcwVTcHW2zBsdQpiN/eWrj
QPH5T08fIzHnsLpYhGLvNoeyXT5oOxa72nXZN1D6TKcLy0CBgaKtrTWamPU+SNY4hR0DcNmECVih
A1dyuQZ97RxfpsK6EyPzlkYxHKJMCCPzMO5G5OcRI+cOuNmWujvZQVnCp53zK1kA5KhX7Pok0jZM
y+3mBCOfhFfJBtZ93pdAi9IIPsO/4OQ3foVtmF6BXyMFJoM4Uo1mgGoAbg6EGWjNcGvjbFfvr5Ou
936vB//oMrMEd2tw8IvDIF+rp8o3L1cflGIYb9LBQrWlYmnTbL3iDvcE8NracJ9H9JyZq1JaP3A5
siioJx2eMu5fISX8TIPxoxUQalfrInSEH2LZlyEW3UOOIUIvQLEmdkcvPDtNjkze2ANz19Lajzna
1sGITGxJjdXBuEZzBQ3/qHIZoBnsARr4apqibLkeHx/tA+CqKqI6nAmtTW29hBMOWdyLr+RMC5Q5
acAf71LMTkasPSdI8jo/A07bvmkhExFfnK32OWw/u41bZfdWKtQ+ksNR860UG1doTYL317vEsEnW
HSCQoXZ9gXab34nOrKdWnkaxBdnx3tZiQdJXtkt9t3UUXij1Np7YCRUmHFaFsG0EHVDJ4ZS9f28D
yxqZR0cU8v2lwi4egceJpe8AiyLQD7G40RmJJzAo4sWynX58ks20dK1omqlaIxfMXUZeelA4Q6o5
/pVfqUCE6gCNnqhLwN5xv8CQd1jF20RaeTj/M2QNg5941vAELdBooAj8mFUmGYC/EbmJLaup6mBX
bQD578V6ivl4saKc86vIVnE3LlVY7Phjn9W2HtdjbdcSKORRD0hPMwpezkw5kQbnN3w2AyTx0lFl
TrnAvcH+qiVl5LFC13+dQEfAxTqWKfc9Yw0GsB768J+uWk/OyWnrn0UYzOqdzrSV31PbkjWcdsD+
IFHFyDV2CM68x5g1bDoAcedIZMWFksNLaprxHW5Y2BjPDLXm5RggBDpxeJwIMK5mv7pwzgzFJdo3
FyRn+B/I8J398FQl7iE18nIa5apqFUXa77C/UvKBNmGlLXvN03qk+8LniULaQ/HxU4whPKd1t8xk
E5zq16tDUduTvLP9YR4y9h4Ssbokv3+oDCWel+SR7Bf1A/aqWHxeA/9KyiQcjQdAcekYLw4mXLRv
zFTilamqL7/X6tcUPOm5dR0QPau8G50oxeB1oFgDINczqqCLws4CbedhdFwMqh07TdTtymDs223V
B5KkqYmsXIygY9x41Y9USs64qzaE7Il7PQxTgRscG2nBYHUu1nlsRrH3U/zY5w64UAT76tFXFeqq
VtTWqo5R41uDqk3ZlkEsISeqMPg5kP9htIm8HqWYebzUAg2Zt4dHanakH5bLpbfkuRTWUsbjhB1+
p+KrrRKlsmKlbY5ggxJ3QZgiqAiAg5QujZ0ITm2zZo/hSj/7N6fkkH/u/E92K+ez5mJns1oKHkx4
iurG5WVKD7YjwuksyUBBeit7ljbX1HqzCyBQcAGcvoyWqCx1quMUzs5qJVQL88a59Nd6ohkpbM1o
krDZsGff2q2vxe10Rpe7TNWOVr7HX9cG9+Ok9JTGDo2sQzqTQd1qqHm7/A1e+20oN2upFf3j3I65
tQIBmazkg3LKHmKggu8tdY4MOeb1Zs+bUFXsd5lBtaQ5A4R+lPHrOkEMBhHXWawFxHqiG3qED8dP
AfC2jc1amOz1UyY+efjOSwTJJwid8e/9ss1lYWJF60g4oUGQacWsITQ70UxmE4c3qDSJ/mp06jYC
OTM0I2sxLVTl3luThrVgb4WZhHaVAi9vAVp2E3UzwIsZFJNRAxLh9TFEeiU/l3Qsee2TJ1ouCYOG
Y+q3oHhA+GoWV24achDQVJBX1U98vvrQMXvlgJPtSvxzD/kpoBL9dPUy6jbxhGeVkJiLJ+2mTCs/
RQ8zgE1uj0llAtn/sNYmK2bhdDwfVvQ+xzcawEk9//8XTkZrNcPGs1VgOAhMg1leuG9jXkrEXGex
GAdHQkn9vGZkk9GBqSllXVhAnE0MJZJdYtyCCm/9BHGUPwymKBiRCUDgcu6W78lMblKxLVfa1O/h
4/MnG0lPzpEF8TZBwO3UUUzCclPC/XkSXZAhRAAY5dzCbeYaaaWSBNyOq72joU1DqRVokGZg4VDL
d2KI13SRj6A/R71+1J18em3duojnmaIYK3bq+4B6nyta39MJROMM8BGBlr+q0XY6lbhWjscdtJ4j
eKHQQ/xu3EhtARy52H9REjeg5fygQE5o/ijBREDjYf9Lyo4R4u5tE4DUax+gQtTUKMWkwz3ji5TO
TmrRLq39jbsARVehcxsMQAKOgy9k3u2zIYBoK95j53eTNSddFPt6xANUEci9VC9vY7+DXD09lugO
zLP/0qUkPEQcNVlQGJtCPXEoKpM77rc5H7nbsLSdodbrtO+iv1V5z9PgWGIRbjr/8720ISC9tHJo
0UNITXEl5RW+m2VawURimQyvKj/mKq3R/r59t1t9ebMetY8h51th2aJ3Ii0Fk4C0fMSAXEuXc/Ys
mA/15++MzX42pHlTPZG8LxxNOj1Qgfpu/lZ7uleEuCxPyb5k6PPdGef7hYKHc5QY/t1kBoMkBEB+
BE2HUMCYrJax65AxAHfmVSiJ8zjkvHUtuBGelXvD59T+2QPu8kwGv17IGi5ioLJOv/O68GLjyfT8
Dt73g1SNOcKLgCRVifHHq9mvLSw3hIuD9hfFNGrxN/eOFhOuNwjbUDhiLYzwKGDw0eCiUSATt2CQ
naOkMwguWWiyv7ogyXrfTcWx19XB04FHYuT/WPNEiqYcMBiAjma7ZRBN9m/QErfN6CpsGpIe+j1B
+Xxlkiu+cVlgbW7nbiPgv8CN9PNbgUTFHHmqcfFQEIROURN2Qb3pxoRehgXE1PQwVnY+dUR/fDRY
8hBbFQqmjkDLun6jRCMLY3UsHpU/2HYQna36lKq7Yf8dQARRYjHYd6Y3LS47qSlJGy1gOhdW35eQ
JK35pi7TCDFUE6xV5h8yeH0EHUJGXtwtQ8qI83ngxnBb5kyolZ3yDTv0uTxwuQ1IRvHVmov6Lc3K
k8kCH6SSIG8BNUO0oLNMX3v0CPQLks+MYy7AMT0acpx9nhcY8BRiNks3uLXRVEPaB2QUq/sLDNOZ
xo51gmRXq9kkfv/yENQLt4ELGERHmIGfjH9kKLYF2Ao7/AazRYdGzQ8J5CYJ3UssUZVBPkXY8GPQ
thXl1bEqh25obx+RCmnZttqIDniJOO8BH5ZHIA8Jh4YOUR/EjgNDtezzEAqN1psde9XXMvdShAjG
Q70bLF5gGz4YCqGniKMMo1PtnjrQluOmHCm0aRWM4m+IQYxd24hezyEoAzdyT0m/whj3g3aP3Ac0
Y/BH/GaEfZPLAXabfn6HEehQo60qJzK7AWqO+R7tYGhjBD63EtJZLIIO/uryIlPBwUWFdkd2Yc4D
voedJIFLZCL5iPkOrZQpXa/OtwHHS1Wb7W5AFvdF7zPvmSkaGxtFIZl6nLEfWyVUFyXEzoJKDPZr
4cD/Q/JiybjDd7qLJGd1jJxGWYXHI8BteOIUqvO+SRwFzUP6kH/WZwVV/Hqa3SO6/MQTdcy5c/vC
tWDWjUWgqNLWVpx/ZejMMrT5g7ZbWS3ON8StWRwHC6xa0sWDrFcDSKuv9rjR+d4BJy9ue4eS7AU0
Wkqv2WTHC+ZJkzOv4iD+WJnBb0OHse08SBry+VWmLWcbHYJn9xbDZl9VA+e6XhfgdXsjbfyfm2p/
9/whPuBwkr2W+sXZETuEaOxBlT4zT0vj6HhT+R5bdBn2v80JHgPiXEg6pYlHu1maDzkR54I5xD2d
YjbFxZhDhE5+7rdY1oki76eL1x5Uv4Utcg4WDrySRiFAJorEnC3/llPNpEnXy1mBzYHpTqzQUX6O
1YRRk/cJOMjJAmH/RU9s8Haz9INJLfZqX0YhIgNv3932HsdaUPFG3zrPHCwP9gjmIR8MW5SUBtxY
aPO0j5R+oGncJYdK+rCOr0Xcejg5U+M2mW3V0tQ4rI/s4VxLCddslxYTa/WXljmeqSu2o+oXVQNN
2CdgiZ3LDpImpB7ELUtOnxNeeiQb0XudiVPTSa7g4kd1NE4lSCPWDM3GBA/UX2aY2cnuvWwv97Dw
EjCGCtmEIXsL7a8cxcbEjMeP1KkccyXii/7mIf+g6rneKI/FznBtTdXbZ4a0j9W8QY6a/OAvXyHA
6Zj0ScIMP8BFRq8zRWEdnRpXRkBzjox0HsIXZi3Y/LLR7LQEtPkLijtd1ZMAk8xIfyO+DBDFneml
b15jdmaSk+HbHRq6ng4xnCTR6leAElV+qVr92F1C1gfNuIXGHFQoB7LYq5iI9ffTKwpdeyej3G12
ijQZI9hLF1FajQNGUZvFoal/xqtsxWYf3mqmOwC+4zdJ6uIF/0fNR1ZDEZM1rqEZToP016HKZayo
t1T1X+UKZFyitO3YCBSfc5IQHU6rGrg+7equqDQNGSnLVxTtj4uanmUhuHHbkZGV0UjNEAgBfYUQ
IKq3RX2kSaDi6/DyiXlJvFk1gQ7X7erh+TUByIfR0rY8iGGCXr325juBTcHguau6tO673yAZ8KJU
blL5wTRbe61fSqN7oSwCOK967kiYCTemFNUjq20uDzfxw+A6QrvNYD2m7NpOcAkRgOuAIq+9H8sK
WPh49qH+99n+oh09MPoehcB2tdbTYmNU47GMhPNP4Hst3KLHO3UVK9IpodTMsFqnDjXYNKPwJbEk
IGt/ySFB9p0ykH0RYZKwrkX0LQAb44MywCoN0OqbCDeVFQVgm7uiPm16HBznTVEy6/YcZgAHogau
rIgzjoYZDbZ+wkBKFLsL/fwBB8aALsFaaf4FJc6LW9ygt4bBgRBCrp/MGBMnxueePcK9JnR9hXkQ
A775czcxW4TKpjV/DnBkuMiO1Ru2iPIY0AK7BEe18oYFzVB/YhrIZecPsmXa6BQjOpXrNvqWqbwh
QyONXh3OLtN8K9+IBl0Z4lxqDQuu43SGC2tFKz4T61ZbGTzwcFQ2VKTvitpp+weS847k1uB38Am8
KQNeLU8yQqrm5IadVf0gGx0niPu6HLWjeyKtx7CHft8mBWayaYGf60255gc+6ALYCayccryWWGnQ
zi9pZzGmDlDmHWUEn4CIUG0lyDU96rW8XxXlB1FutxZ8GZOaQOdy+0azo+B+nqa4oNInkYHO6dTC
sarD399Y6F1UlcGFMdeG7rI0QN2pxni/I7ocJgk620hK1yoJX532rSERLwXhMbwaXlcMGij3sAhC
EQZp9fNuGA1xeTwwgtA6hvczGMP+wShIX8DbVgKAk1zIaEONKQ0a1Fka2D52bv/v8zpX5B7pwlKo
ZPcir7NvYNI1OBL1mFpRqO3HXzKnzRcxzW+pdAjJpQ//RWS1aoBtTGoqJC4qGbgeoAD1tqbUA3P7
NEBJ5HWYXfgp63JPfeUpCNp1UOQ7Ut6A9lJBRe69Z01tie2Yu0FnV9c+wkR/d0vUOKU+rSkn+MFr
4nfahZuwTydUbRNOBDFPEi211wQuURE/786on2GoqohE+Z2tCAhhHgRQ5DnFMZekkmjRTHeaJDPW
8ijt+gWyk3LzWRtgE0rG5UuX4jqDw3OCti19gNV8JpI1atS1CQrp1VOmdUurRvspRm1xLzZb7/PW
DQfyLOlfHfqLAQwQoFP1qvPVQWXr0hCmbRrfAWWqaszSXntWUraxKf30VgDakYPI+ym0T7Mrv7Ge
MxFjG2O/fz+70NMStVVv73oSlTeHL27X6qHmvjMWCBHqblQg61y+7gDB4VKFBs1DpjM8MOAqtCAq
BFBhBKud2mtk3vSw535qAkVuKN8Jjh2aeQXqLTJj8+ywt7MR3NqPXsvXBT8ZIKj4/f70I6fqDiyB
9m49qDDj6YdR1Rt5JJc8sTuy2HYY9ulhDW+eWhFqiykbM4ibqKrvFGHsmxgs07KMpQcuIv/2UM9M
/CsQxI1OEyLk5FfFqCW/5o0nVv64pDdn44wi1XquLs/Xo/pkBAz/LzOFRUSzLIuLiGrRVQ39ZyZF
KP8IfUZO3M3Rc5cNS/81yFfE3qfaSyNBFU9qZBjtI9oO86/ZgrroYZ1yyn9vmB4M9xcVMtDnULdL
csPGRTWEpxH0cVx6/4xN1GsyE9HJcGFOo8a3bVN/vYO4599Y+xt43fZWKXuSmUbidhbbH0rbzWv6
AbPtay2SFLqLcqgpGq5Xur7kVcDsLDZhOkVGDcWjfDzObaG56nKGml2Is7tDMEpv+D/Uu0cLIvVR
AYP5GWcgZO4qBX3K1NH/RCpVfGAoP9AYoqVKEaz+0M8861iLxm3OMplS2tGfAlhVpyQ8Q4FIQHeq
HHCGT6tF+2qQEXJhUHFwljWXptysHdjuGd3/nBOYJDpFmqQppKLgWaiq16hk5WNxIdQF28v25/Jl
yow/wytDU4+UtWGxhDwBSja1oMK7Rr5lh6z//UFVPkNK8SwtHWilRs/4pJp6PoQHinNhBHn5ZQcN
39g368CJN/LL59nygvORC0GBWdeO0GtDvzS7TIk6AhYaCkcJDduiUIxRPOp7p/UMThoL+9AOX2iF
r/7MY9m4a0ezlPEzwxJOtPEFBWbVyhPvtJX2Uf1zLCLjbMiWssTSc2nUxlxTUU1UWaMXXo1FSovl
H1AFvwXB/lYhHg7FcfnYP7jtgLwF3zW1q79WesMegXq2q8BPujEdn2LEomBi9/YgQ9eWtg7h7+53
uBs+omkzyGwXH2v4Ei7x2nbexMy0Rop+7oc+7pOr/yaHkqouqq8e9PirffLrZgVwHf5HeAo8FByQ
3LSxmpND9aOq7syMkM5ZzVgwmXPhh0cK8vMM+F/YFUSi2z0N11CW8zX+W2NGnguepi6z8Ixot/Qh
lLiwgS/PZov4uZ23ylxz8hEzbiIT0hGcJ94JnCuCTDWA+4sJm2jmThuJdw6/Xa0heGiNsbHFtF/S
v7NEaDRu6hNUAusoFC71bY/GXQmk874hQPXUVVMXH1WVaz3S6gU2c4v3+5YayUUVAsyaUx0aiLLd
HZlFUlA07CSPMqaN7wDQclXUBAfvv7IFEKAVHIr7r19VyAthj5D0edlBFAtGUTlkjcw8DvfW0Sgy
hfaOisATzx7QbEnCSR/x//8ovf788pSeNfvA+E1IEehWVrSE4iwNNoBx0HlGO494aLFmnUUXx1Lf
l0SYDtrfmpv1HpS3TT/hvNaymT1u9ecwnjN1++of+QF43Ko/hOukUbhvgaXokrVSqPE2l2SlmnZY
vrQRY6iGUjEf442MObEv/myBYVi6cAzfbBh4bRzCzfKotOKkopQOGEfvD2klqDIDLmR4o+la8Zxd
5AusUtKHFAoxZZHRyYN+Ihcm9pdGM0JzcAbbZnAocYKVvQt/zPkHWoukzHUO+Kx3bGgRJJgWwA7B
IGu9oTKIgo8Fsq9xmgu+xp+9IRBSIgPLl+JRVE/FC8+qhf2hsJcxSywTsd15bwJd9iE38T5atmDL
SwfYKBtrqFHbkD9JFkcgLsevIQlYMS7f5Tu7PN8E/CBxk4YRBKPVHmJypxk/E5KKA7OMW02xFg/Y
jZCNXnjuVcbmssZrrC8k/liPvL7HgPrdKWD5E1tGK1hlXTQOPvo+/lPuQ9Lj6xP1hHLqfzO1xB5p
LMmsIe189mjKwr9djUMLKoYUot+kdRZu4uyIFZDevRXBKOA5oWiZUwG/qZFNZordf1pVP7G+sMSe
wrKkUAdtJ30N2wfjywCYPUfZujk17GNb6acrv/a7vRL8F3s/pr1VrjuyLvGKizN0/1J5bcoFDaqv
+7LdqemeMi0Cjs/yvtz7cHrEyaG47kIfruypfq2uEGr8mMZjrS4Ajco7WTARWOyxcrsgTY6Woks5
UUykfpqetcdEEYhjNv8FNoFbxkrUj95LejHICb+LinNWRgIRXqPvzKE2Mr/aMOU221s7OsFJoK/F
RnajQRuPoIynLYDv7aeNdYz2K2/LT+j+bVd6RyMe0U9DeamMWE+tBqQLcCrhJ2DFIIE6iuuY/5bK
GO8sl+0CszVC2BhQqoEAfcAzqPXkTChZJEk7WaDuQGBCTFHoKrFyJgNWgl1hYJ6SRxv5o7t8UKln
akQLhcVtLxDtKuRkpi/ZlvBTIj4ef9nk3l3pbedMd2zYDoxm2lZwLu4aa8CwcU1k5OHp3BPQZ9NF
ccOAllurfD+puSUF4L+PqFRIFdROUIsEsfPWHfjlRn0w/L6QnkHSvxYir3JQYDuqUZIoqzud0gYr
YvFSGfhr6YSp9u8zKbUspOJPLR0tavAnTfw0cbHVs1N2QFXl4NMb9iX6lq7I+FLjDnG1lbThd7qA
Sg0atB/qAXL/P5CkVR3zpyzInfacL1PGSFGVb3kIRdW2m9axgZby69iEZMPzVpn8vZ2nhgHeG6ET
IPqTPC2ur+y3Cu43D6CAABRmYqxTnFmRkQ0HWZj+DruYIMXVPNGpOoKTjNbdAhoGqbim7T/8GbQD
YBekIkfDIWFtvdmfHt8Wr9TzWPn5EMV9ZQM8mPW46bzVNPtZmIKE1A3HEsM/tp8rwoVRAum6Tub2
ii/v8e2lHBkbedwfHq4QmzXuY6h9ZRZiM4Lngmd/gRm6PmibvwgHboByFNAOgvSp9n8aMUrzPqom
xv24CCZh0DSKie7TEUZLjX2D4utpxAALvC3s1PwENIczIo2uleQ1Xc2ZKe3Nebp8PPYybEHc+UVD
88GGBYSEWKXiKbkRdnvxUhrX4PypioNnFGbrRokl9v7XN9TXPoso8BaI/r3Hb4X5Ah4JX5kaH+pB
ER29DbInf0t6RPjEkg1pQ3+LucRg+3B/vCx0k+8teHIDpJX7/E5lLgelCCn5i5hSJHdA1Iu9iGur
nR1pSorvzlG01v1qmCgyzRGHGF/lD3lIFRQIYMTcpXesskOEUU7g4mYbh/HRZICAWVwqIlXs6Hpr
pAsJX8Ne9edZNR4r9ArPsT1LT/HySkikrokrgzpLyvtNrVxCbhci7o2NtDDgFr4uXShIMPU=
`protect end_protected

