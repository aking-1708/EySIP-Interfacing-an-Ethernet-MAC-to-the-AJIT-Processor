

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AbrLtZEWaMZ9QRIEqn+KbGJaY9tnAHwhbFbsPC7WH49ehpa1EbqXv+qkeNRGupFwZ63XKanLVUyO
My0fDcdlyQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jBjvZpZ5ZMxrEO8+CEfz6CEl8aMhkYM5vXXCdl+QFohneB/4ao6UdzksCSxNPxkQX54YmGSOciXP
wgiPEkvihckzTQ7V+IwmdcU3758CZsJi1jYV4WKld6YxfbWBrziJy4pEooel9pwm0aG1jMx1yNUM
erFXjNZfwKELIgXdp9g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bNlKYiiGIQP+R/ChMF9YxWObkJMdPWBzZKUDypAuNCvFSKj2ODeFkzLXYHokfw+rz7RZe5YojYmq
4UkICxShbV1k/N1YYli9QKFi7npsW0xHaRa8L0tSoNNqAKETg1msjVmjBV5kKgQ78l19v/4te7qL
zUqdthBriU3NcZYre5k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0gJe90X6qrVRqoGU7iK/i5s05zq/0GlJ22Kt2H/04aXbES5oZ4I0aGRfiLSYUCL8istn1JleJ/n3
1/LRSIHwjesRoSy/6j9iedPDLLSSnKq+N+ZcvCJl8gg/L6B9ChU+h5YNE7HqJVfqJzqKWKPqsHB4
WVtjQ/Uh+QwxJp4Q/GXnPw1qlnDs2s6lJ8EK8000R7Any16QZ06T5S1IW5s5v9bKhWJj2Oj7lmWo
6QSr9mTUFxCIV/m+pXzsIOsSgFWqsBmD8jksQw5AorgxI1HaqEa3+sl/imtv2p//6lwEVtz8coiR
PUlfIUpZ3ecBYh1Zuc/GrakwiRgEs/Yjfe+jCA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ux0aTH3zrSOSGrjxNBhNJ8nXWhxNzkLj/DcKiIgChJ1nxm8i4YMzp0L+VdbHtn6L3ZPNF7NTEh1P
v7Gcx16JuF2FM4sw/t6m+FCjX3oHl0zUFDs/HfDB1IEXz+2hsgoR9SYF+bXbSth9Ql5SVw6WlbpS
yFwlhS2eW7RGdfH7yFg8yRwWXcYySMv+L+udV6VzSwe0SODgbmC4o26VRMdm0RBQjLnYxl3eT+4N
Qf9DbWnbFLLU2LtQWORMV3hNidJEmt4J99c08slF3izsh110Cv87/wiU6Xuvi2AB6jI3wVkno8/h
1xSxQBnRHm/fJHMh/8PrydoVk8qMhMXs9UM3dA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A3eq7CQ1ZEC2Oz4Co0wE9eavdVVL5N2w7vnxu/t08WjNVvgkDcorbVB3GWcUKigHFQo0FHxElw0D
PA15/K+npi+dagAdVUmv5cfV+KYrdhCLG+Kvl0Tcm6fhXM4RH49frRlov9a41BctZWlMEXzlO2Ei
69nxF8+cDN/RPLjSUoKp8oVTX2g6+udi83fdCBYaBZQYCaaDSNeGqephcoL2zlXyK7vU9KpsDUWJ
oZshHV12Yw5hL+4YuSmKv1aODQadN1UJ8qyFc0vRYTAqwP+hcDUwxiR48olGBo7U7czJnFk4AkkD
qULDB9rPKRIK3YJacz6Pp3GAHUDGm2JO78Eg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
MjERPvk1zdyyB5fHD8yJTuPsAMmMzBjc8n0yFOt0SQTgcE318TqzBZXmd9cg1lUsH/I7zKhUA+xA
HIPQQ3vE89HFdr+qfxvQ8XBeYN29Inr4Y5BmigUKQZyhMQCxxkxojlf6yNnlXCbO+cSqS/6hJUF1
kcb1rAongMJWAdHDmNCkNV1t0+g0bdPLAqyDr28V+MUJD+gJZCIVC+4pqz9dGJX+DlZL3m7TxS9N
ojYyejzwygAGmFcfQRNJO+XHFugxNlZbzC70xFs2WLHUCuz5r68PhTpys6k+DkOEaX5TdLv5MqYt
VEcaOK0sOGjI2NTo0d2m/+SM7Nr/sSelChIeKNrocbEBXsVClulTYlglKnDG7hVeaYPJ91LUiR0B
rc2amzCRg2Ot+ECDP6vCs9VkNHZYXAFeCAdmGXJ4pR9t/tOu3hEUzfHeG2rgzAT8yrt/0kM2DbFT
tzhyCIRi/LpEsITnbDAdAQMNwrMWBLeSf3NAXEhgKORUJTj8QdYUnRdMQXJMJQD7iVMliz2OQETw
MHnfMNNK1OltNKYpgkRFXW8DQwIWvwbJ4dsqvXGn/ZUCS5AcuK9re5rNrTTc1KmwzPSu57Qk82ID
Az4FhtLdGUuJ2sj/3H4M18k+LwwUSjnG87xTlusgxwyMmga6hQpEMpyR647kFhlUtebRE0/Lgonb
IEuZ/o2dEw8k/h1DmNbQOOPBFyePQfWQcbvOypUop2M1n3IdqklauJeT9LxS3zDZk6QNcAk1i2IL
4fbRiYVyNct4Tx4JEyfVMMfcXgboNiXXv1QGwPov2nP78SkbfdG/pWqrEHGs/KNe9EZ1B1PtKNF1
fP4UlHhOEPvcbR43dnAD1XSotP+i9wkje6uasPUa4kXkV6P6o6J42fSrPRXfWXChXmQJr9EeKgov
TyhsTBIetH85xzNFGQHAMcaU/aGLlO8MrMvdZzmdJXHjItQNgExgmBybH6QR0ZDCfn70gmPZvWxk
pGseCb6BGYm6ZApQW6gDdaK9z3Zri0DgrZlXB71kg+zKTN969diWWXGvacvZJcqh9QPGzilFxOWN
7c+3SjNsDABpPqSf4uGMuO1NrcUvTWEdmNCi1qvS/Hdf6kp2/N9+ccWawEHEWRiUQIAU/DkRA/V3
R6EUIpNbxBzq/vrVLw1Edn/SoGy9Hx7QjhPVa3R9c5Rm+KoUUn+AFtX6Xs3pS8LOEnuV0NSzbu/+
0shZ8OYZJ/vMhXFzAnpbYJffw9CZa8Z7yZ3MuZAIDqVu/604h50cxaiw3x2UbQnM2/0kbmB+JP13
WWeRH0yCAz971XM5fCT/PojbUt3FF4R8pic9IiM+8NcqNv5bSntrzfJIfrdgpaE6i5sS911APHrG
qd9VB7Q3XYBxP+NYup9aD9NhVj4R+W0wtPFqOQYbLos97kbWH4fuBF79bT5wfsKrQ0apB0xAM4pl
5xRGfQRh59tnWNlANwE8L/785WkFTlHVh9r/gAgQ3sUZznIAs9yyjECE53tqwMC+8NJnq7u5K9Hi
X1cDvX1ngJ31BAF38IJOEJjIqTkFWTA5wb0vx+2RPl0U46ViVZHCqoJlE2AgdCn3QnEFQ2kyNxdg
zAGqCRuRHzRHiNoVI8us+RTTuYI85F0+Bc6vcKub97oxbeC2kygkH4DBTelqycYWGiwysqaF01MQ
ZqNCfLkE1ny6cCetE8q0XU+oWGTxz5bItoc9tgWLf0Ld31uDdPGw4Ae2hkgjtC/gKA8cKBrZ3hK2
qs+KY1RtRuOYxdaEoPFpwRZDCD1tavz94ExESJ7oobVsa0KlojG6h89OCV+oUj+Kv/ppOI6vM6pd
jGTHZ6ooStg9WbqRGz0atKQ9PXE3ihE0qNvGCdK9OkXKV8+GYvCamIKAYfoWDRSSOyAF04aJPhqF
vqPTx1wjKf8jcVgscBLCRTkVcy+hQTL1e3yRs4U5BmClYibr6wHdOy5W19SBt0w2BRGvYnnFHUSz
TsM4z5J4StnsXTUZMzd7pMPwzpYTVaifm/eLjXx0Y4h+NAYx9valvLr0t2TAP+sdWfrzF2i55A/t
vGEKNIUMcAv5H/D2bbTtlzuh8L9OaRBbwTcWP3uYgzcQiV1NtUBALbxr5IWF9VEauPd1Pz5pceU1
xyYoZl4pdrUy95xc0BxEWLDITtv0JazJoH4fd1DoRCLprR7sZNdOCFOfSxUn3w+eFibO5ibsKvXm
ar7gdppVr7OxjDvdVn6B27XDxU+j+/bHFA7xpyd2qxX6fTJ0XWuCkTPm/LQoQ+ryhv0GxqBgCjre
zbqdePNlQnBXkkJ6BvjVc9sdz5+54ip3Rk+OnLg1yDPMpUcG5HmCUjFm7W5OYK9ib9ySl9w36ZQ7
YuzR6yEgFXV4W2EeNk46DlNrRhsT+VcdXbattpccIhR5cKxFSyA3ApoU0jgLTYzWo0YMN5hXKvW5
71wYVg7UgN0gSLDzruJ/ZA3vUdBgtUoNgXtHD47dKxs7UsBwEz6LgASBy37Fm/WwaixIt7WEM7DY
4Xe6b6n9NPmTE2gVTi3R/hSjEhjOZ1Q2LfvdpclwkVTX3NeYxOw3vObclvEmPdsAn/A0P5kihJox
wWiOXf7es/81GI+0T8cgS/ymOeLfpZW/07KIjDPBIQ0Wj/8+wXUsS8Gkg8PvQTakZVFd32JvcQ5s
Xf1wAbi3HoMUSLC/9bFxNyMwpR9SCnyB/Au6WaqCc0YZGRjK2LY1YUqt2NqeJwpjjVHr+ZDDckmn
JnCBIMVB8K3EqoDgI9E4wc/Ada0L+XeLzdpSJltw3039HZ49XlzaIx1g6Z0IbNPlYtNcz9xJVSwJ
nWJrzDj8outNfPMqxHSWbydkNmZb1iKMobU8f47I0tuOxKtpBFJmC4p1bwk2NuYKrCeGfme76tqy
4rzsimJh6+MwyEAnIT9FAWDB1NL7Tndb0MdJe87TiTlpTlKqb6WFr3jCMEP61s21TaOujp/HYby5
m2NRh3Etf2+o+a3suTUu2Kd8Ab3KXw8+P+ZdQ2zjSx6uqPJnlLWRH5phbNUpoYmwrdW3yJ0V3Nkc
jWS2Ps0pw08VIAKhn6PImk/oxnQn5dMt5otSHfEULNyyMZUX9vQFN02M+YwI03yQhB4NdoFblK84
L21V6Gig8IJpZId+m2AeSXLieXComiFzpDjzb3SCgrTyUxfaigT1mhQsF4b6iSPI0KYQjxiUeoj1
5RwNPCLuclh3w0QIFTAxq4od605Jl85UIAvPxoMAI1P3139mVFk6aLOqFkBqr/kr7uOfzh1TflGd
kVxf7ggc/jNQJLUeu9dpKOIbQGpNe/fIXRyoNhxw0+SgttN37b9inPtW+448hgaS2QV59zs1lIwm
9DI2KePzOXPqj7gchzWyfbIJsfWkjTa1/vj5kZi+DCpbqb5MQgyYBopSF6rKYpItWpWF1BLOSz4l
pChB2QgfbGOhvagojCUUEVndUsTLAR9lz4yZoA33hrccyfT7924p27cOpOxMcEg7gFJKACl8jmMr
NruxeolxZcwRjPoUDbgTAAdaM3ESp7ukTeD2JjbWRJ5PGIlIPVPZ4PVphMpTyniqH1ohtYOti+bH
xlDJmUJKXhv0TCw6miDqogjBOTB9tDji97tma2Lb+BnxhXZ7bOb6KVHj4LvUi75fDjVhYDZv1EEB
wIUJV3Qv1kAZ2AiGsw4l5HcodeYsjF3GULkemODjKshPAmtU+x571ruWteFgwOWQE63zxMvQABcO
jS8lR8LZwyXdMxQkZ/5aNxK01eTEebE0eTIz1svGi5LmC7MJhnPoXPSvpKvOlVgcGaHcdxtIsdSf
vKW18de5349TCu7rrc2OsWIb5Qq+hRcSTHCVkDZNqWxlR+U21yQrXPNm07rt3vjCj2yQ911wZnnp
6QnUwMGQCOiGMMrDCbwyo7cQgftnXs9IhTB0LDb+AKywQK7YXhfHvYPE2Xu7K3TTpeHdrLKTJVaQ
9wFCpAnBrXmOfSPSIPu/B0XcdVLcirLQ9G+bcz77r3EoQtpZ95akzy8GuhAMajWMW6gNxQU810ST
3jEhAXLEENJErO8I83L/Pq3nGUwyJ704M+tnebJQFLVhU5MH7IqQBKUPk2S5kz7Ri/F/p5Kkgwdi
pJWP/SEf5+KdnAOhTf5kpo+Q5ztFG4EZ9+Y+TXnUa9RZcqjJTkFjJGaVbxGUr6QzbPGvSNL9Gih3
/eVZgZPDw41dVdVKuY+nl4j8aA8DAXx/kk4fHH0swJ67l0hMiDfdj4cxmuUf3mKMR5Ro8XmN8kZy
UrnCKAFNEN9CvQJyATNlL1ccroovK2uUZEBV3kF2HkylhjJK0QOj2cOMq4LSZvhlCQVHDs6Ncl6p
lNWc3zOsgCknInTlviQq5Qz6qsQVJCmiItCvmXDzSxoKzW8pmlqSiR/tLIW1aEzt6EsZ46C9Fb15
aw3KfiHJ8j45Xq6oQ43HkoXMd+08vNArDtVCKAB+luQwxNEfaja/z/eqNJPO/2LuAk8xAVOw2iCk
teNVP35nBm17Pysx9IRvjOvWTvD6G93MwFNVugb5/kvpa3iyfiI4hJsDDdqsUwib3ceD8baI+tZG
a1HyDTa+LQ5hFB6owGELAtWS5W55zeJC6tspIQwAaXm578jmixib14EAp47KT7py6oEMVodPNsio
0drR+y2PIPjjGpwBQsqwAitjFCDL/ewYQUar46TXqM+/DeTqaqB+GYsoZXn2jCh9TnNgXaJh2+dt
Gzxk37z9Atx8XUw1LWd+0U3cRjQquULy9TZG/c4yJZdjgXl5B0lZnIJPFHmFWLoQCtsiKFk7Hb6a
qCT0dexyWx496Qn0sfrW+2WhNJFksIR4uYNZGy3pM13vBmrTYKBoeE58lQdN0U2H1UPdduJUnDqm
ACLkwA/iNucbTSOOxihzSFgz2El69L2ZPvHC03qucBTAkDxpsEjIDLUODm+MmUeqEPKqdAF88KfO
pBp0e18O8kINZbIJCGf26oXVriVzxu+gVAOTVTVyMod7NbspB6OmhHZo2/SkuoPRHvkins+lVcMs
cA70zCnMosy0vrXVXy1xYGMZQHZ8cnaTgUplRJmRAoQPLnN+aeGOxF9XCtndBIjlHZ7b754uSRnB
qeGQqtBLQ0sUJ8EJ6jHU32mdyGTY7qn0YdrMPDWCotmFllUXMLZ+I3NUmiz6ghpckeL4Ed3IAz0a
xkgOkaCcqBal+hOSvkhiSre3EmNv6sajszEDwG+7/MDPcwZ9FGmoEUHWGgQzbrfqeqegGYBAau9a
omNJbNPWvmSviic+0EybSiCPxXAaef1fwdoI5+Wa5yCjAXX+y7NGkA4NZ7wISJD93jm5dawN9pEB
9oRKbqlh4j7w3BVvCBYS3qAOzwiBGJcL0gFlvbR4A3hWjUcW5kseF+xwkCZT9VaSyWkNz2loraoZ
p7BlpgBqujcucEOKfPGFC3hSw/djHFbbdkUehOBoLN/v98R357WNsxNZnz26sbyuxogQfJ5j1vcQ
UGFcrKS24ggIxh3bkm6BpjmKJWCjEeTSlKLyxQf8Y/lD72opO9HRJSe0sTNYBUoZC97PfC8Eqjhi
ISrAckZPbYEphS934as4ntfAQqX2jpobUhsUJNimZA/DdRX6AIuh111LK598z2AnZqxKmhlN2iMu
F/C5O8WsXJe/cQfX0xKUT63In9bdrXLWpCulENnf/jplllkWVWCAoaaMViSKiisGiuOcD/oIh88c
fCpMrWT2HzZ9F+2nJcz6cNpJ4QN3TsKldX+VY/Brk5iXyTgK3pFdcz11IQrRFFPZWqOjkAAlHP2+
SnXOsfmkmoXyp0FRwzq3yuTTSMqVKXC5MLrWD4DFUP1JY7cFf989TSVzU0J0rDuUWk+Kl4eaT0qY
Iv7yglq/pBhzGmefTRScPIXhgaEgEewq/oMYJvPEAM1iMoN4yUtUMEsWET50VQmXHSUmRhauRsEU
egAKCMvkPSgQIiX6JGOS86ajXdP6zJXPC4+s4o7Cdbyys2a6fZ1CiXOlVMUdmiqOQV03bqUTTluO
OETa2F+1Z3Dxi1YbLud8yXMOc20NW3zaMXcRdm+ATVyAzJ6rFPo6AyaUnGH7QyHSJCGBnuTTnSYr
ezUE04TPK23zwsv1yVcrWvjR8RPreMWm+V+sMf/e1BiIinRpnvzNXJy5CBhafPRKLpMMbPVX3oEW
L7pC4/p4H/G6piKCeUH+eDMFHdwDeMryiYB2tDqm1F5Uv6GpXDRTe0doHeCpVxynem62dnAUFjOh
8mAMwTu3Lr4o1MU3tK8W0pO3Ow+dUOavya3oFVjwIP6R4cNjUke6y2evMCyZS/x9kR6CGOcZySeg
IyStbjqvZdqA98cIkNVSDK8LUwLZxPgC7BxCCPwzlOBNpNxPiyP9Ecb3wayV/7Bs5uOfn0HmFaMf
IJup8cGZ/0Ume5+XpjD36fib5ioVKVmj13HpDvH92QYW0NfIAZgHSiYSBLqyWUN0LjkhjguH5i7O
zTUlfu7EBGmC4QO3yfhEfwcQW6j12EEYMYWvQKMRcgnXceBar7cLwcWKk1sfgYshtSHzDwBvJnap
uw3uJg3shlmncOQeOT6d5DysseiPQrKr77WsIgAwZPpFhlC95QBIIWYXZ/KimQ3aVnhIsmykFOSO
KnajFu66ExMmnNyukAI9QZUbbePKKNt/5wVnrV3n4KXav9JihaE8JXAoIYaig/pAyQw/4PeymXIV
uapMlPfhwS+LP5eKX0STZKzgYtaULtCUJ8+cg1quf7y2BIg+3kJLeqC2pl62BXV7KPhqAjbP4gKB
hqegpaJlUCdohWEFnF8gD3gjJYr0J9PhptRpRq07MCOxkVGDcZ7vFe+inMd+aWvtEmJb0kQAfKwi
ED42FVnCRfkW/H594kwWcz2RPBdYL3wdXuDjAqPnyVkZNn5bfj3ec03AftwvYXRm6Kl6iV+JJuGP
Gw6XbLWyMGuf+lyg+puBwNunNFMdLVT6drKfjiodk/JKs2C2KdSdsyfcC6Y5KBLvZhbSUqRbA5jc
2SI8+GodXOJhkCNsll9VpTWHMODe+Z9VniK21qUxmkJ3U8/DGBYf6Or/25E7aOpbRoP1D0cwg7oS
iWgrRGCnVB2TByvSWgZXzNjOuVwN7O9LHcGRLDcX/6OiC5qRg4Y9EmEU1jwPrSF0H9YHvIRj2kz9
6EDzg4HjommH42V2Xg/JQrljUD8qkbLaIFwGd5+OVSGuBBUgWrkOkCvbvfe+9ScX6A6zNCgTz0D2
z8qTcsX9q/2dvDdthKw+Ud4gRdpoJeSrAk43jwLvwJJ+wG02QEmYdbHCSSxr26G4VEP1q+sFh2JK
pe39cEoLJ+fZLlEbD2SgYG96b/wEln83Zu/s+m10N5WqcJ1J68hdnJEXL2kOVUSFtRtDdJXf0mkY
enRnnrFKLxTLUfpW9zsHhiiEplLjEymi+8TpWHr53rH25xFo6QEE7n6eDbR+n6EvhlONe9kpEoKX
ElCKVyY8NGXn+1xekKaMoaOP5zQNW3mTtdkOoONPYDgZ6A1+8cU8gdkAB6nGrpx5mEc33omha8eI
daTr7kqQgNccN7eS/rD4DfgXFHC9WPskJyxjX71zI6ImEHCSGgHlZ3sDbtMngSeGQ+5v+3JdT18L
bOMFMx7i3VLo4spSa1Rxafrn3Ojfto5SqTmCxIgx0d/ms1U51NZjSkNLWE53WbfGPOd4B6/7via3
p9ngGgF4Gceyealma69lvt8oSWXhhcL3M940dmApsq3hXpRznhZXJWw4J5U1+Z+s9+1UTQ9JjLtr
nCq7n+49uUclzS8vdigWU8uVJBm+3opOdEdV6CwJcF/PC7cqFE2twiDDlLcP9EGqyZs8FfIXv9C6
yFv+rCqIO4xE03hHX13AHG+e8u4OzOLvOETvoD1lmpcvYRARp6rOmxhyygEGIg5irzzjtNrEcvLM
K6SsNhHY7bQ8nvOQP6N9Xd9DHdhlMpV4fMgqJw5YguMfUhGVpgGvhySk4pSSo0IRCAKmX7uOVC7G
+bQtrAmRGKkF7aJd543op4J5wHhiWWmXW0jsxJT9XmQ0chCMuUJxs6bEfVYhIJXgktQQDLspAaQm
GIyRevZe8Xa4Gv9lcA7O4D+D7pdIJfmH8xRmKa35yLAErQWGcOOS9ZCMuEW4E+y5r1Li/qyu5UiA
3WurhXayCjvVPmNpA6sPaWwHF3kRKizUxf1pbDSzZEyrJdTKHfx+kTOOTu8wzrngyzbqYvwv0rzx
4xHCN2ckH6txDJOLgvLMwMeVyD5oogFwo2hHv8n4Q5Ybj1556/15bFp76Qd8ssdhxyOBfBoVd4jr
xGxl1NhExW7pusPqY6b5IEqyh/0MwENags6KDTewkJ/8xfvuiz6mJf39iKzLF+66n1kaTptpxPLQ
N3+4nZHRSxSwMIi5j+n8WMLC4B9qQa1H1vG91Segq813QhQoG2zJd+pwLRv8Kn0/935B3UuJtMn0
R7jZaq2MIkY2AFqUqVXP8tOxNFn/gKF6NIBkc+y/2nCiFre78L9YVtwUcmrwva6wsvyN2iVEWmWm
VP+0af6n2WW7Dxxl6fxiVrO10ExrMwMxeA2SI2jSUmBZVlpvn7aFPYb5BtnKrHcDwWkA2WSmLr9k
Ov8a8FbKDsfjTrK5Qw2jSTBipYWDsVnPCAaOtnIgiu+/LyBj/ByMJBrfynmIF+/Q/yCko6ciUK/G
fFUPtByi4qqgx5FghPaMyos2Lncd128/g/v1GO5o/VTodPiLHbCXB1GWVrr17qntcUjmZaO7vSwe
E6F5Z1RllTHqjTYSghxzN6wx78ttSaTvNGxi/gxzHqlVTTmxiijKmA9t0tuSvXmAjTSOFScvFJc9
KjOPIv3cgA7HVPGA4MklreMJx/aGYji0zkc9t/kWbKYVslGwQtaIeVkPKdQGVQCoH4sQ3jRVHyCN
afk2y0WMAnETOYMMEdNe0QQI42n4TmHZslou0jkYn19AggPATjzXsB8aYES5TKLBy0jyMUs0YUD3
gco3ik2OIQhSioG6/WO1RZM33ms0W+6UIkuAFUeWcL6ksufleHaHACyKlW2CVstvQlXvvCXA+BdW
YLDuwKxz7+RdfZ0JEhPuzS9LnPFnnfINjEBtiOt+g0pXIFXhT90MCt3UgbFBUSRuDbHgUMwAXstO
2cwJBhavvx0F4QprnruGucp3dbxKX+tChtIAdXuBwX9a+SIPIRnl0LsjAIFBoWS2QjxIdtfq8uM+
wM908Xg+bm9fFtAgaqRIt/xsXe06G0HMkhqKK8xCM6FoRyYmAA+M8UKAgaI2cE8W+XWvvqvjooxh
kk0RJgkCPA0JHXJELcRD8/FHCcisWmFzd/VYyce9G6TmkGWkBtDIsX7tj/TRndVnPOZ/rHHYk43U
z8ZVCSDaidavrjKLl+1npJI0nb5HLxh9NJL6RoKECLIk0KiJXiKKsXd1yTCvtoIqZeD24NOS4I+X
1zEnxLUhmrVfzNG2oKmSNTuiOtnxoUnKgl5PAsNknfB0lg/RZHEZfrqvYT/zN6z0Q24j4fI7VrfK
PbNDtXHu0Pxdj3kos7JyYKPADa1J5WKTs/zgdrMHrs/lKPIxkc6i6hFIQJZI8ukmTJw3ZOlOwxeh
6s505vvh9F3K8yoAU8r3AbtDr9cTQdhvfaPbqvrFhsACUgnPozetCL8Me3pG6Ez/2XZVMHRnC1cc
SpC2T50RoXDMQlhSRVmD9Tae4kO4HspvY4Ns4xoeTkqddN+ACHuIN6xOjTZGUqsWfyOyTcJd2jae
VGo6wC9oRbqMZ7OvAyjCA9gtpnBz1H4BMlKpqttL5KvG+0Wx8Ga71zPz7hHWcfZv3KgcIZ5RpO/T
AJZdMUmSWLFiMlZmNazAhXl4DbNoUhFoTLZhQdiJvqW03kVuUbm4EzD/bre6klWpEaVCgadHThpw
h5aIxxjBHmp41DeNzTmO9BWrXvGvZsOCWbHDSTPKQS6rtkZ5xiTiIWmaHTP4Ep1hCt77VsIaf/b5
0XfZTUJQSJ82eW8Ufli8G5TcvqOmzlw8u89pWKHA755OnCdFk18N+Vn47we/4LdVnaUQr57Zmlj0
YRQA1Nf96MITcGjoryzMfwgFrndJCH1TR11XB6Zx1O1co/lClMzMb4TtDxQIwn61pJqGf2YolFWO
cierXNfMdW8yMsiGl3UCFBBwB01W0XO+zDQB2dyqd9xcz12X+YcTdUp+70RWgjMJi8cfSot5U+mG
lsF/TYko3y/OBLLnS3rCnCwPLEbQnqntRmbN8ME46TlMpXNsSJg/lt7vjrSdjJjDtC82SHaNi3FS
8mYQd43kMmyyxrP5LfRdNgy9G7f3dCAH27/bskkv6u95p4ErBDyQxL3IxQB6jdmy0bB13/lVl2bI
MlBZJmtnGzOvssThHisPtVd0UfzhJCLdvqj1QRcOzxKUqh78PG07fSEbFUviRK6h9iE/cnLe0z/D
5JDVsitRZXyMJ5b34BvBkGNSjLNJhmkhKvYetefJr5CX+I0pnaBnCycJTRGtgJS7pes9iPttNHqT
YL/dmwisWsikqJE/g8YnSULfyHdap/2dLRzitBRXOKdBGKWY6VBEf7aNgpbDlUI97/KB8ecWNXNc
F9bEX1mhYk+fLIIf8xADHBYbH4mHrcA5hL2S5Ofp+bVZzEtd9w70b1zQI1C++rrFc91eCSzcku9J
kJn+Hnjs1bNVe5fD42B6bp/ikW2qrcXEqjJ77nZy26DssqzYBxbIJo01o/XHh7LHnfSu6WDj+R1F
mOP5FBfMGTxTc85+83oZvDA+DZxfuSsurE8Ymhz5oj86aVoltHVdcDZgAK9bJT1AXwpMJiK7OaHh
PkjKfNEhfPOumBCdERUqShI6GNBukUD1Vp4Tz1mHDdhE89XXFjFyM5Gf7svTSfEStrVYMGDpbtAs
FSUSCtMRYEfVjnjQ1Qn0/AnJdYvPlVG7yQubcHvWN3MWzT61utBWy2YfkwCZx8kUgRSgWwNyV8zk
ShKo4gp+SrAjdGFVnuE6acsL+R5V8r+DPou0i7hzydw/vMqcvkfylj3JZhqHHlaSsf/zH0XolWkA
STEDzudQcfmvKft/u9JdN4ohiekEbIXqkbLnysejEYNMR7Ppx3q5ps6KYI4CGJ90SzxnDrSJlyc9
6+hqb2GMyd2a75aUZPW5d2UAews1w5uHE8M140V1h4LnRA5/MROy9xQHg7JH45GWW2tR8gyBU91R
zfjbo15ElOwPLb+6VQ+CTMMo2CmM8/1v5RVgQx1skO8JOpn9CtgsRn4OJaOKTV+ascKoLBdQGTuV
ltlY35nOmSzJxHE0a6xhO8nsRLZ37vdhodbYNSX95vlhkDNmmEa1hRqwGwuNju4H5h2ZPnlyMzZq
7kbNGt3zTS+BMDgz1Pnn4LwVHDB6JmPGzS2DY90yeTbcc5S2cOIWqdJWR7aBCJhbqPKNASLv1clS
3mkYBv+u3WPq4nIOgSI0W5YXVwIT1uGRHP5XLM3pERR6y3kYAJvgS4PTMn3W9FAoHOt9vx2r+Ceo
Ya90rvZr9btjJs4DBaMG4FyWh6xyFVS+qPRuWj4euwJEUEz3SojecxwgMSC7q8asQJp/NGuhz7ys
wxnrJdgPhhWAJ17pgh+UdXGqKhxgnFfMZOMqD0/ZFJZv131vR/Uhb/6JfniDxy9UbOQ2cx6qaF6C
9+CwRV3AxnF1iXekxeke0ZLAOOizxogM6ZXK+tqbAr90W5QD7619R22p89Y+BQBAapjDRd0a2Zha
yQJT6Sdxe6w2+Du2cfdLLDEZYt1lxnyc3gGCG/cHHPreWTaXSRVoBqEUjh5KOgbH+mRk7UtNgK7X
syiTWaP/gq6EvIkjcnkOpp1fvlW0jogWhYVye7fW60eo2lvcnRPlb5ggHsqCGFyR//acpDueXDdX
iK0dm4f3CqxjOpmD4fQHmOflP5mYBPYriqg0jtBOhBGPscYBRcmTf0w2WdVlWeW9PzY4qR5ueYdK
XlL9a8HX72vygcl0RTOTvKDVEvgcuCrwh2MXzrUoNQauJEr2pk49vZFYfhdN/84kmva3+alslkgj
xTmu6a+8jBkMzI5OUfEnDE2FEuMjQqdp5YgJpVRrrcO3ogxllBKCcVhlTdWKg4ZCMs6RJoMz7SPP
fAn1zcnjgDBI4aOsVDNy0mv1DO9F07VOPs5jgpZ5A04ys61CyW5+ljhxdNB5iJgR/vG8N7RBc7MI
5wIUhWxHuAsUR6EHFIrWeRr5jlA98iJJJF9RG21skaFEirHFZ0YU9xx9bkFZ7/BjHaCliDLMFIOG
/xaMLTJrO4xd+Yjn+FICl6GEpTvhM3vbYtmtln72x3yZz2vMNkgxoHZX20bhNcPHaeH52ayhf2iI
P57BvuzrLhkvrKp4BglKKlBh1l/wOtX4BEe2OQbMbKvX7ZvN9zuf+s/0MHSrh2ybtB0sKwY5mqwr
D0RGixjtWeFY33bqCDSrIID+HgfaIeoHcafutO64DiFEG/TUaGhygM7eb29vSnccGRsJkTPyTm8P
RYd59/bP+6vaE/T8qxgQMHDll5MhocTNc8lViitvFlFI+f62WhHKB+u0mF0Wt2LNO0Z8fiCNPzwo
G1W49A9kmRh8JepWgNXjteMU7facPi5ldTVJjonYxA3TLVwGEhSOgnlGtuL05QXoy49ClkkdRhDN
dbl3zkGm0GUVu/Z1BHKBjPRFgmj7h5ZX9sFwh0W7Y6sSubGzDcH7Bvj968v/k/j30d21xGutXNUX
nJWuWFZpaA22DCRagF2L6xzXaRuh7tWlSMMnaULzLM/LjVumilK4hBmmdlJmjR+WBcuBT0Q2aNen
K++nb0IXTKkW/3Qm4GgZZ4Hwgw+H1UTAQ71La4bH0/EIc5dugoazHi3/xWHfzv02tPzokebqRicA
8qqY+55VLEZs8oKMK/T9Q7dsdCNIq6qjlOkyLQy2+wn2G8/U7m2CkXYL2pbHhyXqAAQADGH0TzZW
givYnwHOOLzpA1LBKYzTGtwyUlSlP6wdZN9e9/dP+F+TPah8xqsIhBb2iD1v2YN/a7xTbx6TExqc
vAkR/r5IQR6K3KWW52PjC2RTtOCBL75dt+HvROJYYNt6C+B1PSjUXRrBHzSsiF+Rm4OBPpAZrHW7
0UAqMUPHeZNBTZMJcBEWhPHkiGpXB/mgwFuWz3UTBWOFUVpUofT0M83e4jOdJ0QKu4Xy7xzPq73p
gSlkzeNJDT5K6BwRkc8qhKXlS1P4SfuJ3KslC3WaEaaqsFCHGmYYlImSRVzgd/TcO/QC/CfA8Vu/
kRHgVmzCwxfRAn4CdIa3xCnWYwIKnXECeMrSqbXtNW9b66gPdj9IOGwh8RwlOsxywQfhxG2bdPZ+
qKr3ZwRG15gksZkG4W6k0TLp8SvS6oGin0YbQTvivoQU7iqp+bXktcWz1FfJebFLfW8C7Wsc3B3c
cPeh3WN6Ce4aT+ghmq6XKyCR9T1DV6itKWfhT993BdZnBTU87t7KOe+sWk1hakIcgvHNEHc7GS1V
yu96e/3rOO8IQwU+Dd9KWjNJ+QgxWDJ+pqriDRHAseNIufBpEgQAaWUpJLbKeMuZ0uJcW6MV3nfg
E469IOiBTFl+vm6p5aMOO7FhCB8Mi6FlRSXbSGoiEytJftUxBiIeQyDDFF2aN25BzAydM6M0lb6c
PEeypRw/2N9zwbHZJ4LBkztwEwkJYqtUNexydWtx50/FqJzQo4H5PMJ1/xcs6JAypkylFhr6+J1v
l0J//1bjkqIpIeBfPMN98/FJvQIWsXdclCJv21p/WURpk8Ne4R76Uss/qDXjBl6OlYp59hYy6d9b
pU++q3FzM48aTmEnkHHZ/B54zIPluv8fzsOg7QeCoZfE//WYtGsMXt3/itKp/eN4xkoXslAMzD5K
6sLgk6XutlIJy4aGCnAylIIxsVVVEXMhfIW+7l+8U3823mG46a37h3v4ABB5cIduPYQX2bOJOT59
4u8Ku88QQ+gnVG3C3SiVwO0nqBz3unARWD7fKGsU9gQHvpG1CcmV6qJqLLmzowji6Fg1DHLyotz9
FyrLkfsnmXzCoPkLLI5/3LKN0LnYzXgA6378jqvi6S7rrvGGh6RH6AtMMlP8v/qUhne/O18jB+JV
nq/IYH7X09HTDhN4Ii5TV9oruglCAL1BaIlKoLISjHAWSNS5EXqc8TA+R+Y8IHjGYhg2L3O0p3iJ
6vRBgQK4Mt3xdxyFcOXSG7GtJp8KXhKPpmcxsV4IYB2BK7gmbW5P7mGbyJsoe09AUH7RLyTUl2M4
+tbsdbtqLppfVvbKbGTNNR60bJ/mWRnuCirbrLmF66t/l6GVPOoitz9lSZzeM/ByxRhvr/8iRZ+q
vJnrub+I82/d1N6IXNuwgk8lUv9TwxKgOOa+BgfzxJZh4lDq5of80yvTUBvllG9x8K+L/YGTkywV
e8jQ+jHE7ocqSq50OJSy95S2b0ukfmoAvaVdR81WjdGDCX5UJ+/wAvhh7CsWsw9KMiakR62NiDwe
oqJg/6cQON+yF9Ww3cXoUPd4Xbmo4wvKjQafChGANt2WtvokYUN6R4aIEUECWew+YkbRFyw86UsZ
Djojh4q3yGi2D+0ppq7dGvFnyzeP/0NSu4+wg6/5hFAfbLmbwlR93hyCPqCULP1YOhxItHQEjZS0
Gd4hJl1jkRN6kzzMtNEDw1xFo72oFM3B7PgMOrXV7G9gqHtqsb8G3CZqlhqaLxhtAp4rm2A2bjJX
Q0Uxql4YNyupX+p91sCM9w7sWj5+5QmDnks4eBnAcPAoM4iB9T+EZEb3cViDzKaDHIM3ohSmDv2+
L/q3nI+2WsMOm69Cy1yb6R+nsDHH8SYoxzzYycOuHQm4batZ9MEpnyficyiSqXqco9fHOuTYLvjR
eNxc/rAkq2k09kbbA2A8nHyynes1LJ+5ejAXfZdIyKoFfG8vJCbd3yUL+Acr4Z0j9HLQddNwtXKa
kYtHSuMxtpnxcV1Nor4UdlrUHiPQe1nlHoXmg/pY0jS01qJWntMxOkWGmapTdz/Vf3A8rgb1++y7
vLi4UjvYx9yLch5kLr+B5fIrEbxYobXrs8HtzqcZEl8oaijWHqxoUGHgxFN2Q524v8dYthDBY8Tt
B6Bxjt6qr31xDN7QEnChINYhfsO8UlIDinCvDKfzKHmqN8ZCpbDIzwJlnzqncs4Mo24d9JWpHyjG
02800Y7YHVT6UjPdkFqJ+8TCeOwePBenJAbx+YPcK6Yl5SLm0UnW39qwOeggo21HiuloviAL/QuZ
lcWPKXYpUdDCHoTsNQZxORIPaEOBfeX3tpMdkSpChArN1GkJ7msrbLN81PXRXqLdjiuVvtEOXnbz
hFATMkOEX9FoKYQDEg+rL7EZ9yXiAviL/abU4XWzLQZolyuaEakvriFtGgK9y39P0DO52+Ohcglw
8dS0Y9qCGTDpNLwSius1sCql0tv58NMGCuhx++vauUey+maD2M0KZysZ8AqlhYqsQu0waYLPnoSX
WLN9TxT/k9+zKUC8iJI+TB1LSI/JTv6m9sBGDEHUV8Jskb4lBGT5EjjhLXmBS6Bh81yK3tXGjhLe
+cnCH4T24S+YyJZSX8GdA1yv2IsQIMWISWcBN4SfQgCVizfPz1AhxW3p2zZM5cGB3xB5485MYyuJ
RoBzoWG8Hb2VuX1gOUBUtfFPEGMvUgajk4pDBv0YSYK3DmNdgCip2SaLIFqjGNWqwyrzIhU326ok
EYJDK+f/PvvkesiFEYmN/NgFgLH0mhXm+nDr2BfmMmUmrDxzZTR8KGK5iz/AE+yivsAP2P+BL4yC
p+Nu79uVTRWLlJzZaw+w9UMqSDwtybBC38iFEof+hOTRUPSve3NqL9IuZVX5PmVF/B9JOvXAkZVV
e0YvFDecbLurqpP79UnUSBCBBrgGiOQnj8TNmTxdL5S97cv4p5aXuSRNj8OwM/suQ1TVKASVigbM
yAd4eQpvEUtVGa14OkpAEQYFbIM0bEyzoRnLMnP8VMgNCVeZI4laltWJZDigFz85rjj9+KfaG0k7
ESX4ll2P4Z5QAxhj1lRPJzAvIkd6ux2Kh4xsNAz/U5YhGY++kZllU4gczy3ebs42geMlnmndvzro
3TTRyRJaR1P5/iFC+omO91mJdf5tBZF6J2fQz4UCpu7fCj/QTZVGVacWzncCYbKL8FoZ+6vD087G
DllNWu4BZedVJXMYet0DoTp1r5bnydLn4G7wonH0T41SpOLY5hEdeKC7e0T5yZVZQcHDMikCS9xW
cFufQG7sFk5twiTWx/hNyjrFUBh69rXyJeIiDxB+dMoNA7Co8Gt65LAiiDo1Ia7TXiQbyGrhD4my
KAjtNaNqiJEAv4C9Gxwar0yAoPKSdSetdyv393EMCTv5r/QqBPixfVXEhzBLOLcTO69ukgx18DIp
ih8VyVBeGw1CegQ5JtSJbYKEjiTb95vbINwwmU+fGISZ59/T1NUoqfIMePyfUFaO//6eIed9bo2m
BUK00Fz7Ore8XLAlP1m4aI0UKHeDmmzWL+V/gJMhebFA81GKgworFw0+4hLcGCfwTaf/j9a9HrT2
GLZFqDImTTvKtkK4Aq7FVysUPsvY2iX8FMz0eM2mYDPSfYpD+QEtHsVq/uIuiw+rpeHhqIcc9o+W
9Km7NQU+4kfi/klhSPR0/nwTxM01D6imPckQwO87ZrPSiRHACYjq++JxwP+XpAia+0Mzs2qJLe1I
a4KsbTNPQ7phodlU8HzBNio0FE7tYu9+6xJdBXDOlqaEsrXD0R+y1TvpjumXKe6zijS10e91novK
YJkG/fVhIta7cT4lSjdcT7jB0261azALVi137W/8eDMZKQwT3Xgk2+Ys6f+EbcedQPIZMPuP2W/D
sJYi+cThTjJw15uuOaNeyntp4Blu+p2y9lq3Gms0ta1BhRlTZBtFwXUXgczg/dZ9uxcbS0CiNlZX
xC3EhR54SWNnfTtXJwTq6ylX4/8I7+wrzNVBSJYBqjscWZ/baD4z323ccz++RxuDDdWRUN+qQCMV
ka/4AgaQDJzAoo70BXY9jWb+Yx1uq+2ftxbNQtzrpxmmIeAA1grwjc1kswCMhrdbTHHIaatAY9R5
tHqqRvV9eoVLgstw0S4P0l6+iRO/q0wP8pq8WYrkUfoNYIjPS9V1266eRaBUkPYHx9krqMPjbF6w
hSljlr4Jl1z4Tz2W3mxUaKNa3W2n9yyz9tWBIgCXDTO6PHPY5XpLlDK2FEYtnFq476rnKxaLLnrk
p3nxhpPivjBd6mzQtTzv4+zxU1CK+iQUQsOjX3ixWcl+VRlYDKBRVmisIHpxyO09DuDtsdRQlyYK
957hxZWLxdRT/SvAQbzyMABBL65ZRni+O3VfShMfcZEngSzbgqM1GmmyF9ntaQorGtK/lgEjKUI8
keDdtgLd1D/lQaCkMtl8aBG4Q7e/yqgWxAfgSGIWSAPJQG2gdWrVx3fpbab7jC2DLGsTfp4gPhJ7
NBhkCPOZjnrMV2x1Pr2Ff4g9gXXHpUZipKi1Hm2auMX6G1aF28OfrOmMlLQja7SZcSBxceQ8Z3LC
VOqyf2P4f92uqrekX6xc2+BhBsKZ4I0Koj4mhqcwTjFe+6SZ83eL7KT3Qm0iQ1nyAP+pZSKcdza+
H2FUhA34/NE97Yigy3AziyBVxtqqjaZZGGKyCfbP0Imw+GVrj6K/yiF9Vp5uSDnnYOakX+z/kSCl
GeRGei5ZkGx6yUPFURBvT6O2kCRhvtAwi/UFr4nIQ8njynYYnsKF8vLKdiddceIuUqS+CMknepIG
9WHdbT2kxLZHhDVdag1nuaMOdk6RMuGX1Il/B1MbiBwM5wktnGCYghaxKcdylD4mxBtyyHBiimRM
rjEZLk4TRcYhn7ushMOc3o2ZbhRNw/1qZeYJpVSKtuLIwWR1nj7+ARcM9ycxi62+14WmCj+K7RC0
7axX2ucqCJ0mRmU5o+Mfbmhk/CB/ORGsnXn5+/IOAOugWVHsuONXGIkQl8ZCzhfIaAQPVj85oD50
EDgt5ordtT6mXRy1iu5DRgYgB+ITQn1E+hZj+7YTkk+yI79GYjxMqOB9Jo33n4tLgMrhtgrBgfst
fwOMjhO5TMnAuRrY9eXT8+A0R9/9RCgOd2K0vqMu9S4VaE0yocyM0bKIsPmlPLYpRegCdaqhAGW/
Iiplt/94h4jumYtl/onyv+DgzNtWYfSrIaHn5AEajWV9PvWS/TKmg1xymM6V6QaNbuwFSlKhatzy
/ONZQAsYFOtUMlKm6VnVr7HVIzK+L5IpifYrhUsJKXCzbxuW1Tu2gqIk7vuyFGc7xxSPKKtmdeU8
PpqN4KE3R7Snxw1NdzIb6kTHp4rx9YiemxMX2vR/peKg1DAahC3qTTXQK32iCDMGPBwlHf6U9wVW
Qa8jT36aZkfL9+Mtneqf3DwhsjeJvoNZK3e05XT/G8mJ3BpaHN3Bc4JpjuwxbR1tz5ajKBxkf0g2
/Y1pCn/fMCaBSaVYipTMxstETnWYp5jh81A61yA6LbW7Iwv5ycKNCmlO5F8JI27c9Nf22/X7SG43
j70X+5nze3UjitqBT9BQr/NO+t0LaRdxq5lxSxugJaEsR7BApLMo9Ds2/9KxXHoUW1qDmC4701uO
Cv6uxwuKwtbCAzq5GhjdOuXtL3xtKiWxJocuTXgdsfx7w/0L5OtP1Tmc6aGBU85V4uFwsEmcddJc
BU0CsQBWQXLqH/WE5YcijXgQtK4qBEcyetyv0tUmb3OqaepE9nXraI7ee8kwQKhTSwT6JGj7hFN2
bhEivkBvYd7+GVNNjEDA+bC59xh1KosQWAeGdAShKfF9NaCbE84pEfprB9VVAoCEZ1JMzydHMqY4
rVuInYVUWIrxS4Z64aplj8VES8NX4vI1PG1CNP9M36YXvrroZimK/iXV/JLUV7VolRpvhv4qRuy8
pAp+oMDN1ZcoC1L21joNE6HYN/uj2BnKC28vvGm1P+jl7Z4VYoZl9eB9NJfDyxmWhTwUQbiK/P5T
yiTi8CzYCm25y3CpfbqOZsCIobESuidjUmobH9e0LaU0e1EaIvuMHQnnq7cAmNZoWixg9M5ynBSJ
J8FoX1OEWL+EL4MGqq1JQkgHImI1cT+12jcvRYx4h0R8r2DPcFUK6Wvu+/1KliEVa8c1cGcgnxju
Baywkreuvk4ifYGdlicV2KLdJcMAZy7POGThMtGWwa43C74O94f+2fj83KZuV2coTQ3AmmfhtH7D
39jTCU/Nr0vdSrYng9iBTux5RYZ8Nvg4Kea03trUD7QNJcb/5LmMJx38wod8uo3GS9aaBcSR3UTc
iizbEbZCxeJMxur5Mp29Zp5QJ8Ch6pSUjoFLg+aTu7YIwZr6l/ErG0c6fIShMkQ/8VR+pK9DCtnw
yUNbsReA5Ix6ofZSAU8CqwUrvjnNXjOcwYN5QNZ3bdYt27Ehl3yzmXogTujCji9fRT8sbEtPxahS
UWEXArj8VHCjZVVwszcoyI/EQxn3ckIZsoNqfEDur7JPhkoG5SebHT/DlQzqfcZpLo/SGV8mZ3zz
Ljhzt3J6QiPFRw5UTlJIVcPPH5eE5uRVTD8MtTUfNUMme1uxt7tS8Ijrfv8LvoF7kmdvppCHw2q0
hGb+xz2QQxBFB+KgYljqXli+VpJh5GqO2zubwWgNX3LlQKinhsgsTE9rICdLkshm0gMRjfRx8DU3
/lhOIYFklBLriVlK/zthU/ClXjPkMW4EsjBVZ4CTlceWmGF8vwDI8Ogr1HFszohpumm35w0wazm3
ZXEMSx8me8OxVVmunbUtT3ewOfzFnlMvIozAuiG691reCbafo1u0CRE7rNV3sM9EBRRIPUHoSTdr
rByNWxUQ0ucYirs9GIKrortdhnE8m/PJ9etH7nIha2WPC6mSE9OG7KmJOKVFlnggBBO7re4ec4pF
cnF6yKd3TUq6XotDU2ysM8Rv9uLZN8NTUf1ewsVPB2pRdI+m+zJV8O9rrImUoUk2mSQ+zQgirbF/
yzbAH+dd//hn/2SDyZPwdW3xCyMfSMmp35IhsR2Q2GAU+3Ns+bN6YYODw0URE4jPfjl0pd8ijNvo
+dpnsA16XrToaqlEl/drwb2olEeiZJTkmaI6LKK5xUcJuPCDiVTbCwSNTqlgu5wsH1ljDs3cUK96
elCbAif9Co1nvcwG6pO56ebeZ5S4X5hK/kZz3pEMLzdUoxNfesYZvPlZgaNifZmYOh+fuYKrvFRI
CI8glpoVJXa6k8LVJzSrYbywMXd3rezTs/Xo/uG2qdl1CkWpAzGeVbW+GBbvMfHH22LYdv1Hc8Qm
Y9oGtkbadjuVCwzcuRQFjPL+/TuGX81xAyCAIuFHCBnEO2hjIkVpvzID4U35FLtRauXdOEhHgsz6
uy8owTFri0g0TYy6VZr506x5nOP55z1XZfTkt1UwJIgnrqV/apjmCA5axonNW6bqzd5NzNqGPxBH
CeQQxyeklh4YeLqGlf9LfUNkcTg7+4/7ub7b5hLXr62Tesr+w8e2n6ucIIa5T+4h4Px+w+Shl+i7
CzzRK7B6MGjvBPiHgtFoaxH3b0VFm/CdsRJRpDHGljtoC20eUrf0JB3JENWF8+YpNX/T8k5GxBwn
36JFHF67huKcslOhBLd85TA7LCwQZ/qy+3DhW3beU+gmBI5O7MaJAmZBL1DNATflKJ/aJwzJbwt2
BC8OrIhkgOI08Ad3v0VUoxdleE3TmI4PbPWSPfSEUQG1YO4d5zTaWSUqwCm0nkm4BS3xvi09+Z1e
EYf9H9Dr4MIGSU/XRg0uxYzjejqOdwqNpZJxUEGtTqxQcxeIR/XpmokCjLetHMN0sJBxIXEixC05
kGyj8T0uoUhmCXVWxaoedAuwbUMn7dTMNEvT4OXQqlYIzRCCgCb6rrQ6KS5J1hkaiq6gMdberzK/
Kfwa49iqVbabEpC/tPkNa1ShRoMGhdLO/3ZBywV1dYtneufFAHUBBQahJrKuyB2VqXY9fpBiK8Pt
0HeDSPLVQMbs+kL7AzFO0osa4+teT5hscPOyaJ3VpMot85m/zAEffJiu4eJj1poWphR42Tw4SkSq
XIBdskE+NvRHEgFPEaf6E0yzjJ34lVIawZDoxty+Scgp5v6pWsgrOHXlwyEc7gvfw6WbFDEeF5Tw
+GRNQgxkt32ZB+HCgSV8rJ2rjkRj6MQCsbNJeqqY5srxeJJ/eybOUSojzhu8FHM9CrgZw4o4QQSP
QOv7PlXb9KF3WyJBUaOIy8Qvsn7fXJMkfIBGmWAsnAoOp51qJmsJ7Z92UWxox39lW9DupRFeWwY1
x/ji64MsMyuqQeBlzOvokpLccXltFU7ZD6owblx48u39QSlF8Bdfxn1KP4BppAMCMQVT44QdQa9Z
7iKQaBKDKwgrWR5OPPyVd/9jNxDV09UK62xHwmRSzALGWRoYZJA3ge9jCV4Ysxu0oXdsUIOEOphu
V52mUSh5HPVVkpnBfp87jlN+ImRHDB15QvaozKZWNXHVSeM442oc0r0qV06ucgm4GvfpnhdvyIHv
RdOkzrBG9LSIT3LR3eNm0ZEGJjPo1/JMgYlIRKfDvX3JwV5BjWmxtRbM0vR75sFYfyH9nUFrAT/h
gbdBrxjSRWopvk1BXneZkoalEe4z2GvJdiDTe+A9ZQmmIzggaO264XqrN4ZVR0YERZpnPNvbf1Pn
7S/XMsGtvEUlcOBJsOmHCMFpI3gDR6aZmkcEewDnGPP2vVm7xLl7opMP7QNBT4BsX2MMVxEVini9
7wJIO8I2kaJ/N1g94QH6uIKvA5+v0+MaspgRtg5VToDrDZNzVF3sEYlWlL0An8pIpF6orUnChJep
HeCwTE3lrpoekrf6rjrHuCf+2C+NwvkO6zbyoV5qD3bfuQBInVOBVIxpwaWfUwi853R1iVIKNgFD
mGe3EfjrGc9HfSs/Do3I8Flkyln1Fkau3YHjjMFYa6hiungNUpLly31c8e724wuBNRW2akZhypX1
UDJcoN03YFFEny842i+n05Wi2PFyiKb2sSL3kOlnudokoGsPzDLZ/lhoQ8TCp29X7T6uIIPZbnt0
88HrrYW2YQ8L2apFpZYZY15LDg7HJ5ZphDTJe1XYCFvsvd3vXwgeCa1dja71XRDepuTzGyYr2Pjp
ON5oYbmhaeJpzHCL+QanBX516sQ3kzshqub75lLZNj6a5Vjn6A3SuzE4hgKmosrda1/WncvcUMC8
NVNZCfAox1/Ho0ErWk8p6b7noAqSXSK+f0ehs0EtlzNwVhWgguqMnLWIxrGOLh+oXUaucpoQjwAq
sozmLOv0VbPCvcEg1kxxZimayoSihpNWvagzwvvhVQGc12jVqiXjpkGmrRHCy4YYAj01nw8ymm0I
CdJ5d3h3K5YVlppiZPqvCTP+1cULBEFAT3KW3DJZLR2iH2s+QikicF0RVW0v4mEElxYOvvAGFToT
m8PtDx+4kvxQZ5Hnpd4CvcXNHOeIMOeJbRxlA6LcTUljnUDNk7lYJeHPHTsnwnGogvwRTBks8upH
g8tPsSG5y2jk0x8sCHrDxO61Wt80tH12E8uBfrQAFHDl0bAHCg4DsUmrPAREIDeyRdYAFW7XxR0Z
rrhCEEDGTzPzKPMNIhApJm0XfopElmeqa1d85MwbqlYH1fkgXubP+NgWLdnXxVIJUeUogn+xMRZA
Jy4Gde/DCTZfSorvHS627wXLPH1gkiM+krHLDNuB3D5lo7rqGTy87syuJW+GoF+hxRE37NOQy2sY
262RQZnWY6p4Jvqfbk5FyhcVpVA7ifqBI5bNoAQpYjLcD/LrhaEQdN4/PIOsbpnLpe7XR0HhCl8h
hBUYhMfGbYm4DM+HyeiPzMxF+qdRwOzpLlbdWRVyA5Bo0CeXy+5x7RzMLoDoIDvB9rCSZtmp+c5Q
LYbcQwsN4NsNXQTK4A/x4WtT5SFK0WmaAlO5rB3J4TYVYQiZbhrAuT0JFgr1n8z96oMw1QMPO2jO
w1i/j3H7hXjJL6HbjjUmwfKX1/mw5BaT5w6R1ZUbZXxJwFSdmOB7PbH5texFlq37trZbBXsr9fVS
YQ9o3xtj13KxJ0gV5GKU+W9BWnjgE0+ElWgOvUBK8y63+UEbBHL5XR6aHsqakus/rO3LhESvJEG9
VaM5TToMhpGrMh8IquzUbhazyslX9+Hb9ipTtdyQd3tCoGYFnvzlpvs5qnS0p68G8xxVoWQkgi9o
zL2bDYFQ59i5+NjAbM0Z72CqU3LduuvDPHLmqYH2YzhycRQj6X47dT5AYzACW4U8OSgCJHwUeY4G
UHshgJ0DMVbzp3gnl1WaFApxOcr1eGkPFgUiikACSe+YRCG63kpFlt6MfgFilOLUrDE0+n1hMkok
E7dBaWwJkP6WKzglUz9fWdidaaAZOkcfTGhlODH2Ma8lplz4Uumn7jC3CLl63bcS8GCj+vXT0JfC
k3u0ZbNbx/4sBzGetIAs8R1WTd1nzmT8z+CDZX9ij9UeSAMzYLzrQGvZFcASfmAyM7pa8Ll6AeeN
kMCv1UasMvyBfIHorOo49NJz6V3fTRDMnbKHSORsbmiixEKkiJRRx7pv7cnW/pP/kXMK+Tho7Dc0
au/YVvWN1pt37Qnh5Tri2TZjmEQuHOLN95piQ4ZhpZlILn5Qc8JvWP8OGBcTLG6GB/sZa2IirAuV
EGU+WSjD3JZrt9imx0f+6Xs3ituFtytJDaR85cVGHlY4DJgXbzsdTM3wwgKnVQjehf9G79e2baCm
UotGaQTxn3pLRTl0nXJFhR6g9RPsKi9h7dKhJ8jQ7YXcDY5XjgN5XotSw2Q0A8+AligiWtcRPsYA
4ww0K5As9W524q3zgMipqTZIJO8u68bKWSj0o/0jJ+EgTbXXdz1J18VbS/OZ/9G/b9kmNisbqikt
PW2Utva7R4WOxKa0omJwRgCQ0oKwYv4HGhT+R0oT9KrqqXQXV5CKXvPL7OPENghVn9CKUDmNxrnt
fHpfg4y774DPCEi8N2haNvvSJg0do4BA7c+ITNmhLhFf2PEbNfyYdTfoF7qnUk8/qXqDfo6fFZF+
eoTbW9qDowA7k1llAFIVGRWQHulZPO+oZDaVhYieZXzAGdI36Htf3faSsS5yDSDF7wHLbV3WEDgZ
2TokRU/fLkO5RPnzKYS6Ypi7ENBDMhDqfwLikfSV/JCdTZ96zKitIB/9egcmX/YJYIS9FmYLxjxE
U86tkdKdT9IHFRQSdm6kZ9EHD2jmbJTnjW0FZb3qY+5nyNe+tzKdJw3VoNLUO9PUk8zZKd7cJkwX
HArwWuFmgRCwT78s10eX5F+XlcKw1V+FEOC65ve9XPFM5RghrQA8xtdTST3xWFNdQxyI/g2Q4s+Q
S8bCDXitnVklg+rJKZ3v1LSyo5MCW4h848+Yax5qoyrkhU85ZyjIrSZ9drnueSWLjBnEWcK++N5f
9IDTRofpC2bdvtljyMJIN7bUwhJ8MNiJceDzWnYQIMU/9RMqlXPXY4uKAHhPbTn9PHxWWjUzeoA/
5cYfXgk+52xUvMJN8DqsPp2Ed6qHW1IjIek8iaKhTcnHOe4I2KxP2wib4WuukVIFNV2J+NDMdtWe
VW8JgmmxtKkM4PBI46EvGWLGtkLg90OMoIvmoPuub9VbZADpIz8ytJh+Abi4FbsSZxATt4cksXcV
BPqNN6uuRibsL9WHiBQFsQ1mmn4KUEWeQIlfRT6GiXNSXzrbDSasZVOmhaUZE5uZRXMUkvDasecX
P5ktoR8VC8C79WgmXIsGNuw3YGdXXHwN9GpenMKSTa0lQ9/APbkUm2V+AvPyfpYb885CaH8nT8GL
3gZPnzum+6OdVvigYcPX9XBALvAiVhbTJSsUL0IeAr1hm1MSvenDu33rmsnZNIB+bIwABYC+/g0b
zuFQTcg+c7Rydd5FwXwKFFEasSH5sC/+tP6cSLYVE83mZDODMj6A+dmEsCuzRgcf+WtLLJH8Jyjm
Pi3APxgu/hKSwxtokXCIulfcJkgfn/j+PNlLeyksN3TpWg9gjFQSu7xlYP9tdY2Co/KAIz6Nm94D
/BvNn1rPHECqt/4ky/aSmvxQ53XzB83CuNVTyTzuTCfJY+/K+jhKGQGR1bPg0V7gP66qMZ+znh4z
sMN+W5rNckGR3v/lmrv7PBvA/3QDSlbsTeeLmtFEsBvW5fse/JZVuzKO5eh9XrHOrw0Ja1seV3ze
bPdPb9KI8YgNEsYWBJPhwJWNjQ/Q7IiqPuCyzevkTtJPwhM8JJFP/iXS3JqIx9ryNLmsmiX+Y2Sb
oQ35VlGRs9LJ7wlsjFmf3sipPMGJBWEmit5oz3onG4SIE8C5jXAJSzkNE5fzIzzWOrjiBFl6ova8
bIpWGti3SyDh4iD1h6/VzeuNvDeWdInYtlZArY4TdzJzas7tZgMlvpRjPHM4Mvv3xmFUUiP0FABW
7O0oXYi7gLf+weTIhRe6jiOlF87hB4S/m/PZ9H+EdjVMCMiYfec0IvQeGbK2y5+65NvbcfD/NyV/
opcWsCh6gMHJrHKSek3eSEKY247blZYOjXG4KeWuMVVsNxaw9rjQOQn5tC9kNdpHbJcSBA5Er+B1
vZ2BV9QX0KWcqhFHuwavoANLbn+2CLn3nw9wn6aQHnFa1NnOI/VjX2/Rtmrnr9HviKYIbQloZQIb
tHz4h9K68SnZgTWivIvU4ImfPo5JbjCI7zxNhJ1l9i/l73dWxMFpz4WVjW3QNg5HYIz+YK/kkmg6
Td8A7dcuMjwqCTOCDlzaRYplTPkYZ040PU/GYvqHRjeqFHz0PJKu1nCcGRjqJMRta5THwHmsd7g6
jbu3G9wEQNshzpJyYPvPpoERauVgb9VjJdHCN/YG4uKhkG1smJr7Tiknf63o0W9pJoAobRnMJlgd
yBiJ7q8gS6TCjBm+n42iMgYB3jzbLR2Q6/5V4nV7SWkmtZQ82dFJDZKgAfM4gesOgO0KjciKpSHO
dzh9jgJivfgj4Y3jZ0dQ9X88XjZeI7P0zmOApXjPxO8qfqaf0jSl7gMTQoygSzdSPj2u44/wwX04
65Zr0JtRHFKxYX0aq7OEjm6Rm1xqBseiKHOvJNuOKg+UKnay+zNaVkegHRZqMU4FnKeI0CZxYPRF
sbbKQILuJPwPypfr8Y5EIOXI+x8DWa5v6V1IiEFaB8VYzNWyI1irZxyoumkX7lSL9L0zmX9iGoMg
jwJi0+zUEMVLu10i48PljWqsd19nLwgN/SeGWIjE6X06uOVRswdFpcq959BYf4sBWlk+MpQMxbWm
TgqnD2A0gHCUTDbajbe44tqXTEzc2wMEUUiJiZEOBgzg6kwGr8vhq5cJ2mt4m3Ld5U1HZ0+UnCDS
Dtfzq6HgjfRV3d284FGsDJ/nqCxioaAQ8uwskaqg5Ss6LkVlsSf/G58jbvAMghGJcxjK7v2cfC0T
LkBWznpLNC8zgmNSEwTU+l5lua8oe7AqREiVjktxyXitn5boQREIx9reqbPcJtDLqHpstOnEGE81
JbXMSFm8AeTBexGNIvwS/Sx8GGbxNbrO6Xo9KmVDu8vAry4YXdyfiZPXj6GzQPG97EvB6rcHXUsa
bpcBSsvcaxPc3RGcjtyNw8SUa2oHJaUdkz8laY/9cE5CKYEFAE2iTF3+oMAa/eP1cA1AaVa/GTo9
tcHvb2kxvlLxTzm6UbstiSB4UQcF3LowbyguiaJSEt+OrxbBSNJbgvDU2y90wdbYBkUrS6dqTLwh
/T/S4yFi7PwejFx7p7ch9zW48RDJ2hQckDN5RQj/2IyqhY90qPOodLTrL1NOXkZkdtJKStG6a+ek
GLIPtUc3nMdgbRJ2DxmwsGBseDGz+L765aj0Ke6KWorBiAl7VFevF3gbHrF3MwInpD0QJOQALb8S
4q6zuWLoCujGADv9mN4UBm2wLwNqsla1/9+9IlgrFlV2fA1oZg0Je/ERpPqFBdPk2FTJJmN7AZPa
KsV4e7oWyCI8SkmNYeWUZlHbHtwNj8SQN3bybQMz13EuHh7hPw1UKHR2N3GujSbdFkPFPKjpFMPx
l1di6wkbMRfpwF3vJm2KwD93pdJ2xaoz7BTnn/2gdhPAEY7Phv/GTSGzYzCdiL797dMACB3htdFb
wUWrCj9Y4raxAKqhgxOOtY0PNU5Kou3giQdiq0XdlIApsK7rSRW0RLGEqNPtIbYJWe7XepSRw7L+
QQunKORG89sRXzApP8P1HJN8/vXAxoBam3HIAtz28B4H7V1tT17/8cpuJXO9arGDDC4Cr+dYk6HN
eCr3NTfH8e0BNk5YzHXNQtS2ivTUfZeSGlWb6n11k+AXtA8wdsSBfeR8nChWTj9JJFkjtsKB6zk+
HIofkxYkB7Hb9mZ6fSisgOns6pdLRGZSeAqauz55l2ntJNxmGZkRhc31QJyagjEqrn/K7Tg6+mYD
vA5RwYMagFqJu4Rwr7gXowK+Xt/kVyrVppedVR99x90dMfUsYMAjl40z1VTbX/KMSyHTT7Uh+Nje
IJmbV37gG8uGTdIHc735B2XygX45Q7NIQUCYMSW8i1wZivC74QmzUQeJAe89owXomBIUsgW841ff
NziOvGOFIWUM04Hfaz7h3GDN8VKPbPrZhO9t32gJID/5rD6vjYgx0tlo3geaOm124lB8YnaZeDPm
MnVkaE7giBDROvFRS5LuYV7rqWGPQZVAADlUPFyaUnZuNWVoVfO91vb9QkfdcWSEZebXZt4ZCxBb
xsffAz6/oCdy8wWLir6LdIJ5/Wwh3s/vvYWqwVkjVyKvMXDkUr9GQt0CFR7AQy+DpJEeIxEFNniO
AA3J0U41+Uy5xn2JzEiUwzbMuWMq6HitPYFXAy1tGG/eehWCHaJb4obvcsv8tNk5TJaXeBl07x4M
4pVK1tDsjI2wnovso657lbCHB/+pM6z0spb7boJO8uxKrZRnFQ0IjXD/AiQh/izKRal1rOxQnk5o
5Pr2HmU7Zu0a8f9XqHzurQAFVFKl6M41UxRroLnGev1fInsSgp401kjbhtPogio9QUgZj5tKvUYc
wvKwPDJ1o84kBkWyshA6CSZZjTNDr/4ezk2wzArOjKbXT+XjXL9UgCH1HfP41xkPjX5xVV7Dx9Vh
3/VXkMc2KGZ7UxiFIQUe4Zx50P7ZKZSH51jc0Bpw1Ed8UQQBOmF/NcO5Syvhu4KEswox777f4wDC
r1Ww3KMyv2Im9Uf7IHLVDX091wXm6OPDh7wceIr25pEILn0l26o9yXYY6rZb4BQRp2gBAU9VRu/1
y4FHrodm0DHCtEeP82/w3ILotFtPVvo0WoF5PPk0fFkCuHcWMSGeEp9SLvD26taVAOwss8R9f1Uh
cBewWuvzDpgtw6r/VwvFlwBlLPGjPdj/Ytjr3v0PtBmsyXgced/MxlACULhHYku5hBEtDkEruRCD
hSgmFR7K7UGy+epbsmOy6nWO0QpnQmHmf/g9DWG4o1Ejb4VVNdQicRcPo8tvtWGWapbVjVJ+URJZ
54mrrjFrjAFjvpD2hyabxjdkfOPjXNyAJkzBg+v9zEB/yZFHIHGX95Ur65xWyz7Z/ijoYfxBcqYc
HZgZJWpg+e7AQCRokwJgTJsC8DY7NNrV3pbbzQZzVv+qRNjdo0VZkgCrXBVMlyyTGm9LnKjDhMxp
apJ3Uu9JiHyga9aoEysxixTNZQfAelPgmU1D5XTKO81RK7FUa2ASe2Vtmix5OqXKLmxkQJKk8UnR
flBU6RevAHiJExIv537xHGpURtgL0JGfnb5JsbCKjpVbU3Jzmjcp5sMVA2tbDs0kAiUwCAiyVFId
zSpLpxMZa4OfRYcJiBxCuJ+Xn6RTU7UpSN6DhX+HpUcnDmq48MCiaJobBJo2cQakpC+q8vH3OjAI
8UYR1jAVeUSVoltCJXC36Eum7PdvUS6cyg40UcyDtMtf0hapg5AsY/kTLj//buNe7mAc/6/s8owB
lhuS9XtQ9I3sa+eQ+LFFmHGnbIkrE9T8Znvda0tyKVxlZHcmqALAjKr38qtdWPxduJAkJvuIRljC
WuSxu1USne9x7nfydvjJrl4xZJI0jH+n5R125Hd7bch76Z8B7rRalAiCmPm/UuZJgsOqTZrTMhqd
aCQZhxy4qPQKsgBQvvFQf7ma8nqbzRgoql7ABwmLTTuDJLt/kVYDyYPZ+qPtgGnssv33Z4Ko0EpL
R/OVvQtlvX93Q6WbO3b/lAWaXSxmowBMVxCExTWYZCoUxyspPR5tayiZrFb93zseTRrD/dALPrNQ
MSA8ful7kHfjy88Hy1nkmEdDQpPLfHk6jQ6grkgZCDEMBcetVORk6e81QdedkrEGFNxXLcmxN1A7
0i1mfxSKWrI4YYIyDD8T2sAWiuX1eAqccbqeLKIwezPjFPA9dYgNUPJZZICv3e0o2e3bEKYqkxqs
wc/+QLD6F9LizU1F4AmFNMwgKYYhV/Bcmj1OBkNnbTdT+yR6gQIWkLsHeSIkJhvnGVwGJo9LylpS
VX9QzrN1QjZA+GTA7J7sxIvfzUur55nuleK2ZUiJwZmfzu4skVtD2/G0E99kGL80FsxYqkxZ2dqc
AJIoGb61Qk9F5l2GfdDCaUDUX3x7z2fn55Q1MPi6GEpE3DSgtxzZntrS+Rgm+7fEMNPvhokAIFto
3hhvyd7NP5GKNmMfZwcjylgO1w2g9lCpyBf0NrH09ajvVfKXj98hXLMWW4gIsvtOXGrOWqKoPIiP
CzmwbaVbaKvRX7YJpL7LfHqGcGDwt1m6wKTlUeOZto2KnVULb3Voy1YVTqU0AhtMeXKWpaoZ1jfd
/cRIwZBOiVaW/oQqhaCggmWHcWZa8iCUEM1atNlEmFeLY8oKkhjKsYE8Rek4k4HSilxQF8541d1V
oKboWdxud5/V1Eamggw1j+xgrIqsYZiusYIAm0AwdGvZLsYVn8D5S230TS+MBqOdL7hMhuTLcG5R
ii8wzo5lqh6Mb7svcTu51DQ45ClAiO5sKL1a6Uc2Tqq8yHUhiGmDZzzoPVH3r4tRYWa3mHG0GjTc
Nz23vJG/Ct61nM8f908xyMbXqVmUJz9hKqgYVsi5RYwLynvKfOiY9MBPLyAAGcMS2I6Jl4DkafmA
bAV19zQnfVsKrt8OmBg6Ixlpg/ushdjMNkFmOUr+NLTRz/hYudGxsU4N5nnX7/T8s+ghDhTXSpZv
RUBcGDp69o6y8wnqeTObK8lwbnsnSELF5Da7/wx+At3ss9RCvo6wKO+JQAGXxVgg4E8tqgckkNy9
I9mD8G3RkjjTg1tIO91SE/L6p12Km8e9PTMtjLcV4FKOlHH/y0ecCyqVZXOv7U1I5VHYsGC/0EcU
ucw6IZMIVw+dohtkYR2vh33YAJY6T4xUPeh753SDy2jQrWw5rCYpbuPzO+XT4Qn9/aR/HhcVCPgo
ZrNH1QwfTEUV3K2SmY/mgnUtxo4mpbYJIVKMQXlzgooHGQSkkUM3ylI5q5vkHw5JxfIogI7rI0Ls
bOYo9kr4AgEjKivmZYavkzepkylC9GIh2St/xhswxANzt0iovSBSohf8lUKAVbPfHewfToM5ef+Y
/tF79HW2kPSb9k+Io+DuFQLq379mYJX4EY/Q5g2itKEIIdwHaXdBnYK7WsOz6dRUhJnf/pjyS4jj
66GqJIMy+QacLUSE9084rsrcCqaH9wZmd4lWrgqCPkt3v2Z7oGkzAF3HWEpjgZi/VqtEo63jCdwq
PE+OjlCyQdgIVYg6QQXHd4GPHUXmNz8dXp1iYA1AKoZ55+MWqKn2SbFnsqid5t2AGyeSwmmnM3BY
ql7Ytfc1eaHI7/5vdZFMXahu2Ml/5H4zoUvpq8m6uDZcSrE+RjeKBZa48pdMYvQWHgRk57p2q/Tc
cKaH9HNsPKdPry/ezT/PmUyzlAwvPrRdtb8JTiIKZKfRPwEDtxKVv/kD/MxLSCwM4/yaw0qr5C/i
vpmukMb6X6UJ00WeUAmsaMyibOIjBu7XR4AEtWrwUbVJvtysI64xTGjmCQBPp1YIZKRj0YQWDQN4
jDK5Z9pc2ia4jQOFtgyQuNnY+eQfcWYRQ73PgoyIL7ajTeiLaiSJ/xILu/EtVZxw6uaYrpF4I1gI
eOFT3LAKVhs4WwfY9WKa9I/E81AIe9ZTHCnyCGlS8JZraGf0Jdmkk90QOTbMZWzTri2gcv/t4QLd
kJ9nsaci/vFYSZo1TgRiu0DycQA5HqbVF7Xx3nEbNbu7kfhN13IhNLPWTAWL6L8++ZFOnZ88Edvn
1j8UQarhoiMIzzIMEbDLb970DMwkJ0pI+Mn1NEp/Qx1vGll0blTf/7s9LctPegH3mm3Ae7RhqoUx
vvXRGF3P+2UCpq0AbzfxqrZYFf1dTXUIGKgmPu77w6u80SXoV5E2SEn8QftPSST8IQHkc2Ir1/br
AgWiOi/3KeQ8vcPIDpOUSm/EHHKCAWrMuUVIEKqOROgo7PqjW+2qN3NKTpxCTzm/HR0VwIoWwCtU
cWufONrHZ4rYf5DE3TW4x6AcDzT5/tp22dFTV7oar/afBqEezeUmZhgMx8G41/J1BN0jlYS7ifTt
aDJ2/8AU+0t/7Y7KvBeA788MpYDUB6FF09c6FvYb/3kcL1yFf2TTRha9IFEi+6BRdfCXbYOshEJc
oY+dBgSXGQGj5mrXEwUSpHfWNqi1DD/bI8Gp3TIAXUC8cuA4tAI9RP1Kvt/YGfB4jMN8ypVN7Rcc
bIIxeqsHsyT8ns6eK5F6yZwAjkcApkA0Tybm3tSIJbzicEFib4lasynyzW10a9GfbHGBLlhg9RXu
ZO6wWIxYV4EsvRgatEXYOVaXl861uoJVGGS517hbIMRrLky9McCMB+XFRbmBkRQN1jXcEeOtxkPG
G8f5kDHjJibYa4WRhgWxge6HCl+PbWrRsNl2S3CLGpLZnrX62hIoedy/BszGrRdX2xvCIMQP6rM6
N2OlzzDhlgpb6KdUpGJW8xJWwVghV1hHeHy71icqbZtMFoDAcKQP9VTgxVjgrMsR7dsiu/x1cro8
Rda3z26arIalWLw4GBsi3YkT6wVLG+eKCD72xGLAOaElQ6wz9V8NtmWZoEi0iljPSSwT+l7Xv1tt
x/L1NxeOt0n3I4EKLBVuCGM8b/dgKqOGn3ecMbmz8x3FlJrOyc9b9Ct47fP3+3a498L0gT0FZztJ
wQEXi8eDvRAxajs8an8yCBHZIMrOACoEXuCdfLltry7dyFoQXunrnozAzA19fUvA2vf0ozZVKeFv
3hbq9uqLZsdRua+Xo05OpI8sAV1boR9ytaWRbPEhILlc8UVZtuz0sJ1l7ab91SEiyNb9C0VGzUAb
Ysu8DtOBHzAcBbQWVyxuQXV/gTytDh2MZG8p+oBIV82SycCRycyurWQplm21SVS4wrOxzGSzjN3K
/CEfYL0/2Xz14l2zkhm9667emkq7RDE5Ldzqmn8AlVV48pINgOfYg2+u+j0EutFwJwxJvNHAxAXd
ZM3jd4yqf9HnfRfdaQt2lXW6Yq624K/dXmPEq14vZslAi4mVfum19tUHILREa1Mh8xShS1ouoQ5n
A6FYPsTqmYQeb5K0UfipYv8qRcX1P0bhENenxKo6D7wnA3B0+jmtpS/yLcaOMAZUiE5ZShStCABc
qJ4YI9qCpjoBPs8DoO7QDS/S6X3uj3ycPt4L5HV5gDS8E31DUl8MGrbK6zsFoQE3ipmwZ01LoqEO
Vofdaxm5nkaL+wcTFZQ8MPxLmpVZFD/pvuWBr/bVGrrRIT5fX4jJ+Q5B8sG+wgxY5mBV7ynZPZIa
5biCetQtTD54I6Ee3ZSc3wvWqYsFL85SAvgjmWuZs71Z8UUZI45ffunVq0+ijmgtO/7Y1HiqYbIR
WB4F3eXLjiWeJOzXVpcTLTfoItoAh2OgaDvWrrjSWk4HljOw+7VN31g2Zwpp/mJF3h04rsHMJ+Mc
/+tSH51XP0zAHJqSdpMNzsdh3me2IAqXWN8Xhd7nbcjjBn/ZPcNVy9Iua+JfWj8+KsbIOcJEiF05
zSQkhMmuSzsqus7J8S8HhTtcOrIBJQp6+2DwPsKftKU1mnGNXhe4OPA2CS6nGbOSv3gpNVZ4rwNr
3oCRAXD/zm3qSfIZOJY2RZYgkdcGbePJxGxXR6ZdBH8hgm8ZbDQKkCGbTA0Iqo69Qg0+46mNPNV2
16Mo1xLWSogFW+jmayr75DITh47HHKrPzApwYt1O3oO3/aXDACjnTP/Oc5HMhnr7uBHL7LuF/qSO
NDumgN9QpMPJh64H1qTZpFDiAwsacWcRMMoWdnSMRxrpG1CPfFvG86Ar2LnxMyho/GnRI62LsQra
xuswfWMTkKWu7H11Jt2VlQBiLAtvtdFGlxWgVCH5O4HR64DRVB++m4UI817nOPHp2zQWZ1QXUlyp
noYBKPgGHpDSTWmJszPEYvbbQZKAIVhb68MDgDQ3jiwAEu53yAwtNhWa/jp19XGiB63AZggtQ0Yv
WFZcyQje71ztLvPjCGCBHIoojp+jxgZf4v/Q/+gLB25pLpSOysLrLQ4Q0lzNy1HaQytiOn9h+Iyz
eT96MZhNiDIK3qkVXbCHS8ljD/vtm6Nc1jDorzUcs3dWXj0L37dqpPCtBcCnTmDVeJaOCZzPyFqI
EP+Exup/q7l+6PYN4U85LJG69n6d1jfyz6Jf/pNgmwLfzS0vERVUEJD0bSeb77/4M9obuTumvmhu
W7aLz2w+imtcpPBtz5xsCBDeppvr5Xkqqi9Jwuo3v8psxSsaLphIcHBbSNvdOjv1ghFB/baQdbW7
kdmMbI/warWUtpbwCuUly5dqUocBTHWn+AAJlNrxzY3plqh0KuGxwUaaRPdKtIK+7c/UQ5YsQATY
x32j9C00hg4GOyT92S5nQYFXn1z61D/7Dhr46LUFFlIHvTgXPZ3vOJeOdwIYpk9JZOeBoWGi4uY5
UmN9HyX9mrRed9cvyjK41YyJwYu0K1MUjaupZ6k4K7Myo9OUldJM0Y2/2jj9b4qPhYpTzeu8H29i
M+D7fL/yIVoRwVJLgdL+XXloPtDn1VPQ/8igOdOTmp5rcDOFa8e/bqfDcq1tAUOYB2sBVA+TEA7O
h7YzdmoMjRZm9jGah3PSLY9YC9LkUrVqTaMEk8s10zNF9B6BKyAFrmKusCdd1CCZc1+eBRUwACra
f323uiZeSD8p6At///l9TpdTp9YzRMbKyTK0wOB+7FNDOuFxzLYZzkjwJ1vpemYAkct0xeV4wsV4
ME1VXigxJR/4SKmpHOiE+7h3rEBxDpWzxCb8uYt99xqpRae/aD9b+U9j1eHi5W4kpRc89QLD0+mL
mBmsU24vf2STeckieLBerw/d5tx9suE9HdmA+pWcJeBCJcEf4GokhPN52+ELTHRfF2It9zWZ75Er
MdOo5gooa7qNp+qvzvwgyo3hd23E9D9keuYng9r9XZUzMqiz7vsShWVLAR+b4NIK/8RvDRveaE8/
LrcDsah6AcjwURcUJefwOxOs8Bj/euLHfDrW0DSVYkOHocG0Po0V9D8ANHLXrPWs7HnC/+D7CTsj
PH9L2FyQFBF1YvPr2Ip/1B+PZdIE/7SpIKPmemhQ3a8hBjLVaTM+8RBkBZzjRdM7a+9p6QtimRKi
WUU22eedMPWdLllcZJ12UMITzTeuvwfAAKJ4fznbIBQto5Pag2Hm7Y6njmNudqVtqS8DfVN5QXqN
z83MuKE+VUjj02QG8N3k1+Bf9q/s6SGu8AdjxGAr7j2mV8NQU3lNa5ZBDkmOJKbsNnDPzFfG3xIv
Y7XGIKzfUZSCpCq8A+io70iJoC1RxV9yLUSmZijv7nXe3h73MuEeWdyFuy8xGh4p34DVbHf/pJlZ
M79nXYEKd2F9vR+KQl4nMCLYeQFwmHTPbAAmohob35wk04RUIpE3HxF2aR1lqD/hSgvP7d98sK6U
oYGwwnw6nFDl5H/x3or2GW4c0IHIFZfY+Sk6cq/PTMBUxDwSw+QvLWfDhuCv1/iEcnffuVH6zdLi
DprXSIp0Q6mmWss5AgqWmEWZxUEmQEW/gWH4Z3Z+MIgsGVUgnFw16AgzLhvfL76JkQBSkFdjCG/p
xz5pr1rj9+HBlF1Q+zka88sCIK1bmk4vmqCIrNSfO7ztyMvv6elu9S60WjyE2pPdbBWpDF1AXk17
twWcXZ9B6i8VBswYUJzfNGMQezUNBZth9e9b655HSgVgWJ+t/ZABNWLUTtUCt53JPCDJfSjYjO3D
ljcYIAkliJf+bR2WzvFEJ0IsCE4QeELWdFmbLYQNboq4kzBGHfBWAHI7jAiqTZbx2a6r+BQIAFHO
/LiaCOXqRsE9D3AAXxQOqyIFAoZGgv/smtydBOCkI8s05JfAAIlIlGR/HvRyq/rLLOZvnlV8ha1c
0lbM6WCtVay6GJfLMzx7ZTc/QARSoWekZxKmlGZAP+uFr61mTvGCf2FTbRc7AvYOaHQnbh9Hi0DX
2AzPA6T1+jSmZtfoG6zimfphmVzDFtuP9EDGwK5wd1rgskqISfLwSsKtJwD5zXaSeR7X92rYfL1U
PgIAszlvQHJID+e4vMdhi+h6LHSBstGBEUJ90h+hFnBqaOb4XSXjGxbTBGGQfpq1wnRBNwukC0U/
mrl3MxLS19bRiRXQLMuKH4dbTh0qfN64YnN7Hr6Nfa2CfjGkO9vk54yDOAxib0NOLLsvSxK1H6tD
EFmlqD/hrAlI3aF781W2XhAOA3+/q2mqu7/uZDhX01pMQPnWnPfyiNPiCbV9wsgpQKSqG+z5dprb
5nvV+Je+5bUVQm0lFEinwoMf0FWKfivVK5F7fDK3tDK4FMNWX0Mqbbz3ZeXtBCDo8crfKq5gN+Hg
oS4R8OR5kn32hXL6+B6UVLEyeASkwEUW8fk6EisvqvoDIM7zyM07FNNd1TV+ek3EJAMVXlBRYimX
hUYrwNydRcWHqzpcKC2MmSl9H0TSzKCiO510eqaCxwdAPzkzXKx7LrZlEl6jtnk4NoBKE3c/iW3M
a+i8qQ/+EWQV22QUdgtzQE84YOeuHmvm67ltDu2Jf8jXsaymday/0gQaQZFAhs6WWtjWEeShAZC7
3XPiAXE5uaTBy6rO4pXKAuGTwFkb6Mg+mipPrKfX7f1hLY57rldc6hTLhkpg87AWiBAdDoIoTqVY
xrYhlCO2w4ufUT8ReSEba6KkiB+/pvrh4tXH4DSoFxtkL15RCjaok/CbMToe+CPFFIT8SW5azPfY
7e/e5BaNRvXz/+A3hmo/TfPC/Kanp9i/kuHzZtFYThcJ5auMfLQLHEbr1v7Y5CFF0N7ICmpmGjnM
zzGtOQSrQskciTQPFQNrg+ZbHIzDymTYVvipd/2Wp39mqb8YKSSypQudT8u2ojniDxHU+JxsyuLR
FCeY1Wchgz8D6Wmu7EhD3T6/HCpZTvRuP2GXdeNejlWBvZ0dFjlGtAuPPP45pfI6oOauZ8vz+Sbo
DgRxn70l0OPq/+cA8L0XrBlZYk51d0e/AvO4yAMVZoXcu1uAS/Z3jpLZ0mn3EVKgQcstGcazNIqu
TfkS/BeAoiKJA6WHIzLqTIjrT3kmxQ0mxJCaXPRNHgb9kAVse5zKGNkCOLbIWfpof2J8aeAW7Fib
x9gGaNIMdcASjNJc0saEj3/zrZeTAGJ3WUakjKhdks2nivGCzW2s2v8xbO3rGyD7EZNG4/wIlsL6
HzCZYpr8FlAYTFNaJDSMnzMW2OYu773RFMM8C0ldiNHr696UY59JGu1qymSw2//RWKxlsI0uM1ai
laZeVUxA202yZFIUgq6PB3R+MIAXSx5metf1dF3iqrIdxppdd9fvYAeIJabAIS5qwkz4bn55lotx
P2AzqhypFi8A8P4PLJzdQ3l2mG80ul0FP4QrdsUBoWCWU2MXdHWPkcRObIwevlOzlJM9cpYp1Kjp
qXSxIahCu6gPwRb9v+DLZ5nGRPF1ZOM3OrIf7t6BVEkFkH4bCUPP1E7MS8jGcwfJ5Son5bPpQnkl
Ss5zaN9Y/7SpoO37g0U5nX8NaJBRh6xcCqUSsBSQ9JnYF1tsFXzRF8kbDyttCzpo8tN+rg5Bo/Ge
DaNwb//+AtUADQlAxdLOOwkKx4V0o77mc4JF4GwDtzOFUuY0MkUaaQuMB9IiMlPNA3wC6T8Y6fXz
mrn8HcAM9Yz0NQM1Q66Y/+KjkoHRZ6dzBZ8sucxVRtY2FjgcPHtBX5iZYVzRvLVazpi0f8S+fjX2
iT8IOnvyooIOKNHhbqRCs3BMwbD1ZwZ3ik2jxQy+NKLDSSCBsBZu/fdBO5ZWigXTeE1bWzr1lBSK
5WztrV8iu3799YomsWe2PEa0acBZEVESuqBeZWP417cgW605vZL4Q8nBbM8Lnn+aX/SrgZO81tqM
gSDsV5r4HPA3DOnGwScif1526QXTFwCuRTyQj0wuDXFTtkwqaF4MikF2X3G3NMkn2hJjnAiXb6IO
39iPCdHOX0popUtgptZ458C0BHzF6I1//sJEVuPyZc2QcLjrWqXjtWQU32iri+HhmuYHvdLfseO9
3TpYkJBDXYt2kHt5VhvhN9kc7gNBpd7taX4BnOy3TFkArlsPlQFImXnklfXDLTLVOAoD79cNbnY8
Cr53pGrVGrCywCyqaDumdzH+ZVPPBAdqWekTTse6lCOlx0nF0Hd1miBhZt4M4honh5C/wPPBd/lx
OX7yAF5sHyTIchQXSEC5olzNZzDdl4PJti6rv5D+LNUyor+5+7XmUYAbmM/HTmAz5IaaSBvVlHn6
9/xhBXR5UfM+FFWEQen12sYuIYzwETmWzL7HN0lJ3F0cvQ/BAE3SdeOpjvwt5y6nnnVefgWCKD14
oE90Qa33QKrPWu1D64EOC7qc3cXDdL83X0CcwU6ieb5SNkAhKWDKhBTU+vit3LSKCM5OfqaUdNS1
9A2gLXR9tpY5+E7rSjmM1ULuRT5rUZLVnZMnPDVePfKv5ng4/EgJYYnfYMWyPx0f+gD3uHHNObFf
+EwxDgdpQtTxnTtOFXlGUeyRUzFrESSLf0KVtBYPt5xJXRfb/YzgH2FoBq2bgAUnQNP8p9NwMBNt
i9qD2mxsrSFk3mK4XnBQCjSTA1DLmZyZ+40P6g/bz3oZPeZaLVISLGVUggQ0o4NwILf7N671YtQx
HRgytvwgXEe1UZqyBe9AZ/qSfmgxGDA/dqZCATP5fTrspbAKqIr5YLmUiX6whkzkmGOoQ43n/S+B
ManOZhxz4mxYs0NRBmJ6ZHHJ453VFttNHItlNL4rfTmlg9RtUb9EJWUQCDR5uCNSjNTZMO3MbW8P
A5HbF7FTH6brKwVMnuS6S0+TIu+GYp/2dnllWDcsWSMpWSFNk8ZFv1q9UitIl7W9gfiKtFlKSfTV
IZUOPIr7vzb8ytmoIf4dYLxpaVUP3+DhQ+QSgxqaiP3iSx8ybKFU53cNlJ8dnaln/HJVfqzAmhFl
FwY/MdzR20mQpFMOl+y0Fdf4Mg2BFfJTzxxL/xvQqt7YnSI1X8O8uZLpQ2V+EEYpSdHWJ0RovJvb
AmzuBevEkDT1abuTyW5yLOQqm8Kju7zedV1Nz6yLRwUAFTW6y6llLSrxE7SCxM4D2yLDHpF9JHux
vsyRKANWUVLzyfzljxGuR3OYwI+0ofRRhi3UEqfSePSVCUkeZrrxzFZgeypiwFA7tk4spo/hhdly
bmpzF9jvZqLE/7JDU7Jp/sl0T0IqLG08Vt7iCxMNX7ccbxapolTycL1rkfOJIB5UZw+dQIKyQZX1
bnD+dB0aMREwiaON7W4z/eYLtAnePOvlIwTP02j6YF6rcyPFuoYUUizXpFO8tXGgnT6RvJD7GT7R
pD/YP0P+HcQO9UB5EUV5B8AhHkeTi28Bj9cmklwaJR7H391pRUdFlEXg8M/p615Q5ZS9jxxVG+53
gQkIwFM8uoLaEcNLwi69AbIXTYMYeE/F71uFtGDLDFtAuGOuFGI5qYQ1dIj0BXdem4v0GVm5yRcS
2JTkf+qNEUkKQcs99k7cbH/MW05PJ1qCKJOf9FoHzeiOi1WTICBmumLrXFS6iSsZWVziSHBFK+xa
gvkffGjTCm0g0uXTLoW4q6qUNRnBiQaZyAaij6SOojMBkzztZLEyIHedFoUJmEwt7M6txvGvF1rJ
BFLi7zOg67qxl/14oSdkCujKgvZ4pW0wi0qYFyJlgNkwnqOfivDeeBehmMQJQMd0Q514B9G8E9xn
VvsYu8ZmYuz9sKJ+61b7spxmMSHPolMOM7Vrob8hdhvxsDMk/v8o3uOj1WCGabRHsu5yX5FMWA6z
iPA54Xfn2VDfd3wJopBS8A8f3ukyCa/BaU8ATRPBymkazj/aydJNCWNKIMqVHNhbyVWW810OYvhf
CJCR0AzMdr1jt2/UpydgQz5/auiPl7TOPKNvkv9JaaWydy3QTTxhTvEyBuI3DZwXGpRwmsXXd2qu
a6dMFa0xu5yJ1BhElZ/d078w5LiGJtpymhIAhKH+x1cegvWqDObrbObWrhMyoJIgsDK+NARYs94f
dhpA+cChB7PYZs4S0VpInDjLZnujEZgrxi6zLOFzzZ/uV/dRBw54t1IFVccAvODDlapAZXU+GNe+
bO/5Z7isETizj6Px0dZXoIW0THJFZZZUNX099BlkeDgqGBfEa7GSQ03wWj7pnOlcnJPSBH7Nt6UZ
Xm+1C1XkT+P3z/PYmShXGuIUOLgi2ZO/+qEeAwba/wTJSMFpNTWY/nII4Kqsrd2ZNGz+a+QAL+jx
G2kd6hesGbDMSO4VMA76zXQZ2WKCZ/ReCoMECMx/mXrFZgfKFG7gOKGNKChnvrPJIpO5LNzy3LmW
NLMWoozDMXwxtnjpQsuWGGYseQyr7mTTEIYPnV1BWf7wt/ZkUZXVXh0nqWfQ5fJSmCNudTD2um8J
D2sf8sLk0KanuXgnZ1n/ivnTFnzpUUI+4rwNG0Fc3JuTyHcAdmm5lUgb8oWg9hSqT2frAUkisCTk
sINb/jZbY4gu5eRPQKEdw8n9CJfXQ7sGhIZ8xkqFbi85bn+ovvCfdImi2MzoS+kr1NKZZQRkfEmF
MVz7BJ7bWKhikaf8Wg6uhOo0Obrwex4U3oF7+BAOnhvyfqvp8w7l+W3FqnNzRa1l21P0fFNlwk3b
kCDHnoeVNHfb6zDtHBHh0mq+5lkdydTP3k+RuCxZUNaivBRVCpqzmXoTeztlAj1d/sbOLT2l/jza
RyhYyOxzvvgXnigMEKMOdIm4jMlNcFhK+Q6Yp9UWP498oK/AVIz/LuFB1s612PJuATG/kdoG4di5
aqKyZbEo24qJAVvl6kifeUZ3Q8q0OcjOJBUqJXvNwf7y/qy/4B7rvQy5L318uVdhB03z2K6fWsw0
U7dYvCkX3iMfrbG+uuNI/ZlnJiLoVCDsI0Y9jc6wcNg90TUgJqkzln27VU8FE8sB/WhI/JDIevM3
WxSgAutzzwugl3XSJV9B8538L2oJjc/m8/KGQWHaWLIaQQl3Ftv2TjbhYSY26+8amwKdvZES9M5W
gHW4nh7ByxsYmXha3SJhhobyyL4Z2yOIeQtgtclny+S1r3Aszlxw0+afSnnYNJ5N1XetjMu0/G+b
Ad/ZseQNzw/Kch3N68opKtb6Qu+PwqDjGCqS7wFhKNLGXtgHBZxmUCfj5EZW2grxCIvnSDZrWL4U
r+j+/OtA02WxZdbuDiP0gHqfaW7v6Ap0dbZVJ1vZb2QX1CgFSg/k61nx//trX1Lr8iDiYqXIz+E/
VcvRKgYvdp0uAA8/+RTpoADypwupVu7dFyznOueO4e+bvauGqtP+tJqeAwvL0m9tEPCJL2lvtRuj
AC3d9+6xof7eBo13UmVWsG3tP29QJEk+ZnssZ9HNwO6ZB/wXZdFjgE/oHiyNm9S7aJzsZ+6ALUXt
iWcHWuwkpCHlloZpCEtVKB3vannuRGCXIsg/E33DbbdaUQAJ/5e9JJGB3lzHh4E6ULF4Q1P/dQxj
5zMIvQ8HRCmMtN6D65AeQXQnDYoJUE3rNgOLPYSIy3EoXupHccdVuCBoaIiKkqs51xhKP1X5Zk7w
iEwBR2UuiAjR0Xqk0EGfXN8HszQWy66lWDIBEr22wLHqIKZ57m+P051MXLNZ4Le7OXXLNC97QAJf
5R5xSwjrZ0hubSsIEXSraghu0+Xr2rgGPoAKo4sAG519EuGeZfsQCnhBWHxS3KE7k/o6H3ZcA3Km
IaeFkMdEPIPPUePcb8DcqZbh+dmNnl9CfwvW9ih0yVBiv0sMabPN/N1+/eZYZ3EUdzuIsxRTVHse
L+ojcridcVpuP8J33IN2LAqLDqymSVc+0KzVRHOOT7Bb3FdJ6HP3/I5jzVMVdBHxwQ32Q403iWlv
VCUJjxhDsXJxFh/ZhXAaRFg9pd0wdsdbzq93Rud6kSGNkutPrGcJbmggv1gUjvtO3+yEu0DSgh88
PxART6VoA02R7vdvb6m7bty8CguLQkifQj4Pq13KWMF5acH6LuXMc0IebIT5ntzOhmwjhEmGPYh4
5ydK6k+CpyCcgCGCqHNRobEr+bryi3gA77piLtQX61Ne35a83l0JTF3k2G+QBEECLwzsDZYimBN2
BtUv2AGw7g487mG66b5T3bTafk7eRlw86DQr20SzSUEh9wiQ6dy37+4vJeHj2Kek7eH8lHptoDuV
iKRIyjl5ZicOL+usnfAx5nPZ9scrWFTKu9X0ce8mx7bkFBqP1kdVYQDiAIRe9Mw5YXdbjNBYEsBa
zdV/csGN5nYE1DUmT1rslsWEqY2X4uxal1c9qiSRguYfN2B8Ua3UQLPd7xuo9Pm21q5iJ5ghQ1IO
UIHHEjsK3j9HAND3J0pRJkwSnoN5xe3rA8QDXV1MBzNXKbprmMZmuz1G+KXuxvl9qlRHe55mX9WW
DDWNdAE9Dhv83zqrKrAPyN6ghqOedAF0URyzVjECuNOUsHjQCuVt+rEVPU9H/yXJDBsg47LF4v8s
+AC/DN55LzspWixVQSHV16IcXB6j+hxHiXRVabyFje3IHAcdlH8NoBtIxDmcsi9CMso/CnzV+tCo
dKgOh5f23rTTzIExc9Nhy2AU0Ladnp+dmyY+IAc/NR/6PVB4lJgWLq/aJqu+7T/rZAz87neZpylu
kbegmpqvRzv2WblfSZe12j/CPDs9FOBkXr3xqHcCPIieYguVogQa1pfET7NTPcNV9Ijndq1sVZ0p
ZJPII/vqWT/a34d7WTzSilbgYCvusdlRJ3nxnUE+/18c/uWlsUoos6/x3I46/LDZ+qVm0FQ2P6O6
LKjixA/vxng8qYyvmFxsSwWGWx97u21wBFBhpYWRCk6nopcTZAxOKrUbath8sM5+XrBo5sAqQW5u
PbJp4JoogtCKIQD9Gr1E92KkJf64w6LAjOhoa+Xi4Zf3euW/S/XiKn0YOyjjZ8qk54mZUQgCaqVp
syqlOB8x1njDJLdkFruTcpCtjUxPgiyDScakGPWl1cjCyicpiIltb3XD/nCJ0PJ0otbPLm6qIvXW
RAw6aK78icsOlpD7vThfOGxLSYqLT+Wrn33JalEsu28747Rv7fX88nG7hb6JA/ehVc2DjdInxkz0
4AHywrcJDfLWfyFjarupFwTkiUwjU29lRaMsOedaiueruxaH08hIKPX9cXQPAzoB7uWe1g28Tj91
YntttXqpqa1E3M5de2HySTXL+N7bVJZCc8K2nYIdSNz9SlayrhwqnvX9cQOMYAL54tuR7r6JA9C5
orf4WhagtbTL8OgmZ1zYo1jy3JWeMH2GWxY+/N8H8lzMauaLzQolt72kvbuvjAuCZpaKNJ0bxiOd
lweRTvKCcECiW+NA74fbor6azHg+7Sm4ZxPmFnN1FTr3drnVL3jMjjzsBdWrgyq5FEyl5hG/ebNd
SzQexeQ4oLiaiDQ1KTEMRDsG0bobYr6IhYakL9/S0Tohx48ms+mauMD079XAD/QPNuGtiiU8/2t4
JwHdbT3z4qxF8P5UYmZ+jAKZ2Ww+SXXyFdAYANkBMNFo+BwZUB9b06dBkCoFrcfuKI+seHxqsfin
G0vyyxqHa8qu/wnsLcct2T3rTI9KZTDXgpfKGLQ6oUkWsGPW2C1XrWOgI9u7kwokOui770npyMmk
d9IzNKkcXPtECc6gi5BTosCNYEfXdnwOjKT8lsG1IoYN/S1OscTs37/wgONy1xPacAvi/7N9yVGc
CBy1SpK7Dx73tzhS67gyuErBIEmJx0c5tbtHPPrvvsOxijF8OYH9LRuxKpb//iBGSQtT7QqnM+GS
zniOlKTnhSvZiC7Zn5zZpJgiaQI7o5zPcJhKEJ9Px8qAzlC+t2qTiiMPM2gibDH+yoCDHS5XPx9j
PE67lKkYOjbkuD7/kFrKVmYbUi2JSfc/K5k1vWeknP7NELRB++4diiXLPyqYgwONeyI5A8rdwx0J
7EIMYJgU+94UPemwjT49szLv1/zTflf+jK6fR0uIUCLB7xO9bN6oJ9WBK2WQeEi6PVsrAyJfnHri
lmEPVROCU2wQhWwbkLRtIg8hq8T8q5UPN42TIVUVoRQl6th2VKiqljkA76Dd5yLChnfI4hif38Vx
qa013mJxd5mS6n/MV/C0nuwVJgJhZPagpQi73EnLx55zd5Gqo8OkgGv7JF0SXG0Wc+wpei5q3N/s
E8ilZ9c0YJ8F76hwMvzo606mD2/kuPzr+0e66mt+m45AOQGV6NFqNiIQoHZrTaAgFWSNwBwoOU3L
mk9J6GqwQC/hl92tFxGR/mP23y9uC/5z72NEzrBAMiMzDWMIdDIMFOTVXXwh30RB7gxltnj9wrb3
sb8ZSO79KSHlF0urDF2qKACmF39F1M1gMhg13ioAt0x7yLabkegY8IKiY9WCsHVHvjlCFgCDKkEZ
QNGOAsUGpOKSxHV1F41/zoPqg4ctdSuEUnrAsx7kAvoe8YLvzGBV9XG0628ClAXA/7WjegHTMzY/
xmVEtNNsbrJbnA9GMtbah7EH1o85ZMGHxROz8o+3NNRQ52N1NUFbWLJwiBRS+QLuANb5Vlz/br5D
aknWZDayzfMb3vP7g9dCKM0W0ZRXrRZm8wbsj+skF6XsXLXv06HQkH0wd66fGwGlhDdKFJAPcajZ
dtqIFK1Q6h+OqSNDvyX7dcWJjVcionvUr4dXJGpG4yc1iasD2YADIhw7vziOSQo3kggeZ5mrVelE
/5qEf0XQZEEbGyQsyMF7ok87CzImS2xqq76i0du5tisT1OPldLeFdb9olcAw8l0t2zBFyQ2RnmM5
tyiQMTYJahTtsCZsGVvDTntrbhWKFbISDJWli9GzXeG5FRaFReJBkdkaBWukKoX+wdsonKZX74p6
WnSJZmddmsz3ZPIkUH5hZBReu8v1X+2OQDZqrkxh2o+O9rJQLbUbGMCaEXciPh51T68lLqu73/ul
YbdM57PGigJ79X4FSYjZjI28HzgMUWZoAFBOARPJwwDdKN9jKbV0juwyMM360RJKHrc8sWiJt/Ii
gPelKeaxabICmmkkLAoKer+w3Fk0iYVtAmiK/QzhJZEXN6Fkdiml7oSbAbcOltt4/fAyVml036NB
8E8X6zjE+slbYWtgn21Z9Bp8C8uAQe5HNaLS7j04jOdozEcDzGFoabFnoKwBPhLmzbBeBle/wW2J
JAYtOsH/eb6CvRuZFsPC663mdxebAklm6qJJv01zRobrPoRWFetVBzEJYcYuR2tHx+SuMxJZBSGM
aCeyDu3j77I6Q5CLuuPdn/0ipwtc84ViT1ZlDd9e5P1ufF9/bZ4TFO3gusEtpf0n3p2xmBJhnr3d
OwHpa9JsNOCXXeHOm3CUJxP79wgTNvAeefadkMe1DnLPqz6eK/uqamp78XOEm7I3i2h6gZ2LCPzO
EeJBb/J3ftJpWJIYfNQ3pCl4H5fwyI0vmK7pxquqiSnPKDBhHgbsWe6PbkbYkODIAua2uOoxr+HV
y8dUhZmuZtjYPS8TFmZYLIMVyD1aR0BNOAUS6YWeXpmLDk8xM3OM0dh8BHlR8iJ5py9BEsIthP/q
ewZnHtrnJJ5CCVUu7nYETPX3xp4vIN3UouccJyvkS0zOkXhuhNh6Lx8ySj3fgcGwSUKDzfeSfg4h
gbSIHk7Q3KlS/PUJFvqbXr4ehrnH51V4e1PplmKj4DAoll5Issuli8JCPlfx0LWVdrpA77ShGqzn
MRk07PQyVHxPvq06iUzmzljtb5unvhuus3JYjijLQPo1JiXXPPxX7MgM7CJ/Q10aW599QOKpHAD4
aNGxr6cAV+8IP2Dk4b4cXk0DrngV45T0AWuBqkfKSC3HfM0srAedyScQLtfd9BbQ7IdqM6cQEJS/
v9HBNsvsEZFHgK3c3o+FllIc44w6Eed2LCit2YQeXuZukD2oEeZ0VVlhFjaYNVWDWgyUFkSfzhL5
KdZJ7Kdrxh+rnmxjvqR23ncKRannjR4HEDo7b2V+JxeY1z3TnEWE4AvLQVcJC8Yahkh/zHaWcxso
46H/JsxC2sIJvIqJAcDP/2AJOal4cTj3VORLo+Qhb6Mt+2Z4Vv94C+3iZUpwuGmxCFiX9l7nBEvi
JMIG3aexxpn0+yFc9DnhucMekBFz1fDhnYu1LMWvxlC+IS+HVgM/kv4vpgSDuB/IcNIkuTFH94dO
hDf3Tu0Z4uo+vICePwEJSo2rDF3SOsPqLs2Y+rWYL+fEiQjCTWjB/E0sLWP+394yjNhKVjWjfn/n
EBmmNi1DTnF5YgzSBuvsiufJ9kcylYWH+CCcVcX6weuzH60XDP+Wq4Vip2WtD2sbKo2c2KRdzi9s
J95PfKg8Ve+sx84D2qiGl9mCx8Pdkm84O6jD+KFeoHayIkWzFCVkE7NJyFyB0iEAOQ9L8worR2ez
GzRjzPm18C/m5+SZnphYvtP7usNpQyNPtwQFvNrTf+Qy27Q5FZKDqFxuGSF6Whu7O8Y9qVkOGEHK
6QNRL8Og9vBHoq6TVHBC9XBGZzHg1OKJsHHOaitKn6nBkYldoVQ/wSzDCC1HcjD9o1zzcgX8HV+y
xYpYutF8rDqGbcyI2HoRMXOJ39NmLrQmuxMhQuYR+DZgM8x41B1qPW3d7mjQgnsonfQgHSm5mba3
idki+F2jYcqx1JhybRsm42cBj/1c961g/UJ0Ffuys8VCbEIAweIvMjcSWLdxA5zPvk1dGfVOxJrb
rhSUSY9qo6EVxcq0BbF9RWzp112XDG/V76ppuAkhxrY250xgEVN/O2LCX+J8ArG4ywk/oEu5gZb+
vc2buvZUTfncmmkXCx056cKPuk1VOnvkDGaGD2iVJ+rcWlKQnuVIlKEpm933avYmVlZmHtTwSTyY
qZfWA0WhXjMgGyzNaVsXMl5ufGOAu7FgPr410Rs5DlO6gRicNGlTt9l6dy7DcVT5O/bG7XRbUOyd
B9jJBWHV51U0Mi3jT86FZ0gce0OE4Stpze9dYBTYBtd22dQTGzFXBsAJGpDsGVPe6piDP1odZRF7
MsH6bBBTGeIkMs4R3wGdUeI0L8S2Nls/0KwItzWXFUgavOXJfhmvymO/clsoKJ9zb+tyAF1AVonM
3WybXq7+5xJO5HDif/msjoaD0Cmbexb3SumpKT5SGR+Vs2umwSWB+EU8yMBgwwxe4mVwV9jgfpPS
zV+cT9Coh/cM7UJnY0Dg67RUMTi3QCSALaqjVpB+dyywEb9Zj+/i/6s7k9lDvBY3c9qUenvQikQO
5T7BwjXiiTjYxwQs/Xvmtz9ByS+E1AqMMn1iRi/BUYdkP7OPaU/rtM6nmOirVvQONBqUQfhIqQw3
nNczxr1B5VHe/7Wmkgrla5zCsZQ43oTZgbsKxS6NwwZ8t64THm4D/MD7DFJnxo/8/SdoU8EoHfa6
yukdGAtGZx2HfEk7lUus2ZcZNvAkdP0Che+9tskJbSNiZbL2gq7AkNe1zL/T3xQtUWLqoAs2pE+a
JHrhe3luuZlQe+OH29Drm3u2jpBLt4fSSE0bp65iBLtAqAu8hVodRR0JBD0enBHTvGCpHudizPSx
ftMpgL4pRJq+uPVsDQp4wOXArgTn3sV9s8mROyz6PT+Kl0x+VIySVdBpIgzDmshaps3dxqINpoT4
MtLKWsM4NPopa2CF5s5dqT/uhZzbhyb0dMGAE7kwekZ/rLjczOQicuBcf0pPtDKk/h27giSZDEWA
mlsoA98oLFV99HijoLABF+Kqzj4+C+iZat7bjzExniQl4HKyPyyXfre79KEGf7a0MQkPMMCHLpzX
CRULsAARtkPStvY8zLWgmPz1+Uclc/xhSWtQJ3BBoAEVxZ/0XqTijRGuSIMYjczsqIkqz39In7N6
kHcTo/g75z/6fjGnTMcUCaCjiY7g6JaVzwqQHU9wSS5Awz6MYEXy6W4yCgiuTxwBez5CM3RfHJcT
LwJ/X5Wx9F2UNBsBjFJrdngURPSptjvQ7fIrkCnxENpImI7V6eXudJpDJ5qGTdDcMQXFYP7Fk87y
+h45t80Z2Yktn8TOGFsv6fHWL9CDniZ9D1azQnkjVgUAi7M/MOU1WuERgLcLn0zTScAslCfp10fZ
GDgTERo64d3ym5mH4cPcJNpwK5b63If9HpUW4WjIJY24sjWIgQW9Tom4qaEeUqZ4FjSDnXztDLZP
GF+nqjdEa38eRfETGw7GxtFHw8JNhsEruX/xkw8nVraATKcp47JN9vmyzq7g91TqYwI4gswI4PJM
kXuoX50mcoD9wSpWhL2hPztaoEPey76Lk+uu5uB9ETQgUsQNA/ma6I219xoto72pyIuNHML0hjI/
jkEUF2oe76OutEGi5qPD90HBR14O0V7TRE52uFd+c86D52I12z/lOjqcMF3gvrhBx1hBp2LIUVI5
x/0wshL25JOCMBGjxjAR6PKPUFUVdKL11ZaD4SYJFJWcviuBziBavKk5yTdBBYKXUmRRw4xMlzEe
ZMJRPGzMH8/uDXabwo/FVmR6woMQsP8bzCJN4NdymCuHI8DT8C/fOg/4TRCP4PL0wjC/cjKxZuFF
YVihGoSa26gyokHKUO6EYXSLRreHJvJcdpNexOs8ukSycefDPL1WUaf9XF2nXPTsR2s+UEIaSWIa
5MxhTmrwtcns/gK425XCpMLz7aKA9yXk1hTmOlHHOI7PGYfBwofU/5A44HhCZ8KAHweQqzi3I/vw
Wi7eXhvuuBCbR0mq73Qr48ewdz7E9/Ay7k+wYSNPGnhY50ymIqPvPjR7vJ9V5xA76G2GnR3Mq/8D
eyFKECQgvR56fH6KR9PBrhq4mVnSdxSVIDOYixlEu/xQqm6fw3PX2PAkR5fZ7nuX73HmnmKJW97o
myD8XVcklrm83JQYsHDmSXpX+h82o1Z70JEESbF6KJwhZPrg5s5gH5+e77i6a//S+BKxAzUIk2Yv
ZSlsACP7CbQLKsheczUv7k0n5eWLxOWw29zOCt2tAwW+g447V4FT8Tp6mvdTozG584N+B+7weVuT
y0JUEdGPSOVqWUJqw29YPba7H2eTG+2OHRC1ha3DovUFAT6CDwqbKjsWJRqZpW5Fd0qc7iIS6Yds
1cQEO3GMgl3skJOfXFMgFAiCr8hjqS2VtdSj5T2GuUnr1pSzj+0m12yet1IqoJOYJQUkxHoMrRW/
ZWs20ETUvWt0JSnLRUHpbtfEmwGn15XpwXXrxfJIv9JTHUnxSu98yrHj6gcIdnEw8w/BYLcvANh6
qbqUmSgXDIexcEr8IX/4gsvALBimTUPKRREAi8MthQUKjFjsQd/7PVkdfArBO9oiO2yjPhyd2+bf
Z+ZRcS9bUD0OWJ7Rz/xMcX8tylT40IUAs6aDvFOkNBgbq6Tg42gCDVMuDRiycA4urU+65YnZ2tDW
dgMzSI0/0TXHTyFUccvlEejazs3njvsO0OtgDN98RpouAyjy43PHB4YfZPBiK8UxdfliNKWmUsOz
9rY2N+4lbNrpLvLYiV8jk4eWjRdOADrYK1BNzatv7EXr88eja/WRgBjmlF4oK9ORlSSNvGOilJwJ
KW5gRqzha2m3u6KmjAoZrdOarFvrkp3Nteq74lEseKooH56lvjVXzZSMyMFGWjjtfO0xw1h/10tN
anuHn+U9cr2EpmchJhAIyaYkrcqGfuC/AMkbgwggfjB7tWZcbVc0MyOA2x8CtuZvweZNkzBHX4ut
ZOvUdex9bdEyduVD/ngK7Pcoyggj9rKZ0lSms4OH9+AfvATXmzeGKuVzSCZiADuR1dlF/sIlzrm1
5WGo9xt1qgmOyCSnFr0Xs4sE7sY1U7gfSsAfEXti3RMCkHFAWZ3dWv7bPukq1xJjnebH+HVnTzZy
/0+uDbWlrXjgI+yKNVDrTBz9X0zCPaCyx5TajNyysXCVoeyg0Zz4u6JQvCoJClT2C2Wslr9100tL
qY+KtIonfog223RYuwhR0p8VehhLUrz58oOyrZm7NXyWEfjmnPCMr/gxYSb18br4KeQR4QTnaTuO
CrrK3U5zYdy4/eEDjjLHwdr3KeklABTD5L/rQ+81O7/dbCoBnZ62Tem4Nlg+SKN19HYAZ4U99eRB
+wYhrR1QWtmQl//qYqwFI4O9BdkLnHR0hHMf17lesmYk3v62tjW8zp7uhuLLASN83RKJXyfhdnMB
VswG/baBlPXDVnSUSawv6tvu+mWtlmp0UOVXbne0bMRkg6YlcsxZeNxyeHllZWZsETyWY2Umx1RI
skelT4mOn/4nS7NVhuU55VpsJihVUbHmsm/I7kerz4CyHYDe6pw4v77aUsUe1Xs/9567QdfJbb3r
5JYXEsVRnYhqnqbqrGnbp/Rw6Pa9pOK1WH7S4y1D8NxPl56sfO4sD5PAiPCocdXo3rR7LQIXaxQW
KBfAQedgDJvVLHrzc7V54fvvLC448P7UlcHBqRg05UiMutahghzra7eO3e1tG7vZ3lsRe/sRT3XI
ty6R1NFp1CUCY0cGb+gKGUwC+2LB2ACQsGR32KDllcm5zM0tpDpOscu9/Dw9SxZsuv7yuScc2lWr
dVF4inLGl39bGzG8TPcrbqiMNx7GCck+SZm1OWiIT8eAoyvScmd9fTYc1fnq80qdeLqfJFAdGvQk
BEYh6iCon9TzUKfFesA6gGX2QBYki+T8xU6SFLPYdgCPDFe/n/ESK2fwtZDa8UwPBlY4W2ZKzj0Z
nwDDdSyUsFrypNg2UKKgrUsHjOLWWm7BclnQ9en+CnJRPhpEQORS7ZtLl39OxNaKX///87EIyUF7
1S0+nsM6gEGrNME9VeMXP5lkkzwz1JvG42KFgaB7gGip3kPg029mrydRrWtJj4Iko04ZCjWPJyto
9jSB0dNre6pXILrMUWgbAuwWeL3bOliwCTo5oqir477T+XiKny8X6HXqoPg26/CTSFXzgL+d8NYY
Vo2hTIo55TD4LgwGTZWHlL5s6o0o4+q9+DBBkixtKwIOciq84IEmllozzZ3CkEfT3SB6m/mK+3ZX
3lNl9fRWU0X9s9muZj2YlmrPoNzBmylSiiFxm1zTG2N6J5GWlCItqBJqB3XVKeFlNGgj9N3yQ1bh
ydoTsKZtAbPm9ZDUMjgWKadyhdVF20Ptdel9PBZFrD/Vc91Pg9NFKlXJ+/2VOLKZbEt5ZmYsb3KP
TvI2gq6blxfVSCV062rvC664dWlVl/Tt2WD2adyG5od740BIgatz96a226sc83F9VC6corOs9+xZ
SFkEhpSjVW6Wtfksfz9jmAwMkBmXb+kI0F/r3ZUAyw2/tJNlyAlM9THKaEeAv42weKoLVdpdqem3
e8bEyTJxZJXHYktzSWL36xPBlPXcN5i55upX7Ua0JZrM5YYWi0Zi6UjbsILf39wklFwm9b1EeIBx
QO7ogU10UapLAVVs9QlrtP8auptHs2EpLs4zQ8Ltn05pxfgVQ0bJH9UsqWPcfZpdCtK7a2KYDmlf
5jnkyqFnqm2HOV2+Q8ceL8PtImukvJMaU+dzfEfi1+UbPc4VT582t34ZkS7KXmflyYiRgX4f521q
b79TSD2OBYHLmbiOd83C6RGOtLodFMs7YPYB8lKIylsLWyAywnpt2ctRdK5ceL4Gf/cS4iNLJeJL
Sx99KoydGH+Ny4VrL1yb2/d7AcW98rqgAPPHdZyTq6PidL35Tsx/spepdLcIoLISTSLZhQrnu+RN
IPaZ/ZVz8fs5JWY8dzmHYV8m3aATt6R4263AcmRrVJ6mwSJHVId8kAAXkkbZp9rtXDOJ/s0Kt2gF
0/p8ZeKlD8yaO2In1K9z/oDmOqG6ZwQ5Pfos1jJYF2j2Hl6PArmVQCGCyzKZ1khVTmzpLX/uhrM4
XKwlyEA6dY42UUV0fXdwBu3upzEbfW4U9v3xwyBNjBdcJH+A05R4o9RMPXKAPiQyVOhuqpmOE3mC
olxGo+2xGZERRce3i29/5IKc3imYyCamgy4B3qxOlz4Dm/NJIgvlVtJrACyK1yOke+ods8DN7sgK
methwpCnNLWtgz0gmg65skCKhsSzq9yXf0n3hpxbcjqXaAZovhs8ZnbutP8QrAXVN310pMY46JdQ
3X59zvebOpD9D73aZPkd3PHPaGES7pZp0OBj/TEVy3uK1qaWzOKjonlATnrDndK6+OrwY8WpyhJq
m3O/U2Y2RDhGvZa7yb8hfVlyu8LHvrxoS5sHUHHmO3uXrpFa3mOjCcV7BuBdvay1BwI3qoO7INXX
C9mxl8QQKJZkBP98y8LjtHDbKoKT0nlpW3EzchckKGebZdXIGFyQN1eHhu+kTYzIkPTXE8z8eN4W
2boc8acqL+hP9ARPQjarBsvnbybSPJr9GFo7Wa9UWe/QY0L4U9dUbuWZH841QffaK4jo0XRQnfXP
xRfs6qRuacxjwp7BGLwZu0Znt22AK26vwkL/tK8gf+gHFGr+UiHSUdNo4DT66M+UbaVwQ5gFTmOM
KmvZuAIva4h0hNiPh40Bh0uKabPZD9YZwomD0y/wqOYbA87ctiOTZ1thwg+AgGqBwOjcdk7H8TWl
cVAj+s3kV1MYSWYCZ0+V2vMbVncAy71SIJ755Brd4ww1A737jDhhpl7/CpdeiQyuRPU2IrlrL/xI
v8daJ2AfHsDFLHp8PcGp3/6+R9pVd/q189enTuHRh6fdKs/D5XcB3FhMzvvJLN2QkaIer+x5o4Cp
JNifrZLJR5Bkz54kP/4cJMyZqCXiKWnhwKZm3fdjB0iZ4SsOq+DLoeiO4dMeBfmwkdVYUZPDoF+0
R3TXuSUaTGzeVxUOSt2UWnh6gdf+udY2P+JFVhoNtU0QDMkvbnkn7F5ZJ3naMrclVoEp3Yebl5Au
37oLzmZsCNOsQomVkS/E+0nZKbb26aco6c3NIyuR9CZ3f028BNpZJms5KejTFfBVVSIeU7i118bX
z+eIYEpbT5JwfjbwFY0plqUwqgiH3pd+wxt64lV2CJI+/tjcP38Fhnrv/40ye9ZAEpfZZfjkmOBp
KPhTFl1thEvB8v8uVtspNXd88UBfepu84fLe7wsseDMvG+WRzZeymDRHLd0kIh9VbqUQ8wiQvmc4
lCS7wSSgSfPKYBWmtf6TrZVzdz7dcuv4IU1uaVuKDgO4cuWRZ03hsuxSriPvnRONfXEn5Ukcmcd4
vfUky3UsWluf5rHhjdajvJhJHBwKCNm7ht+Jb2m/fUtbdrTyg7mzkGfivXa6NQIUUOJadeVBItC0
jZItDKGVbyVrKFgf5Lrk232eizfGBuLiNfSyi3khjliUt/YnbQeWISD4ITIzwPv9osdLyIBMxgdY
FNhkMJu7M2h4etX+CJx1CDEa3fjS3fkBfswhfq7XHj0kP3J59gGFT/t7xeVCpHB/DOXvCKuE+Qrv
to0BptKtqbE8ZliUog9oZrDJH3VIb3NzFZGW/YpcgEjJadNXR1Fu9GUP49QyeeiQqmAuuIA3/a9Y
RHgbnPSiBXlISrMfOWzNUYfF5UWWZ9/voSTLaATuR/euFzR36PfdJDlvHYHQPROBhrrrM/EWkqri
sW1YJiwnVxL646DaGpuF+7C7Wsmo31CCtaAZhe4yXET7rEnrb+C4x5BrX41pVVR6LTAIcmVwP7PM
AGUIDQq6dVHStsKEg7MYURnKUWHB3fxg4w3Xkms9sORp5ksOaqo+uG/d0oW9W/OrXWvIdAW7fuc8
KxurCUSAlBRprQB4iTo0oKuFCoCMYfXSEm11VSOSO4atrcWvLCyQiTAGLWIPqrtQ1Rd0CMA0Z4Lv
f1kCH9rptEtYbvV1Mxrj6ghDyqp21z8vVuSJr6igkS1K22/no2OM8Dm/WtGHvVzWomQHCSrWCCB0
zsAM6AlGin6JOgRjaHkaGVhevA+vPYVic2IQhP6goyr666YTHqGJC8y+14xKiHMAOURUMul4DP9f
F16Xi+gGmi9ShSSSSdW77RR7AzfkVRPo3VsqkGnIxpN2UvN9dkubM8RDHIljGI7Z9vGVipcdTIUE
+TZnVJrhj8H7oD60yi2D2RpiYW3Sc4T5vlkB7sxtGm7r3nyN179Iod8XaF+TYc6XZN/t2oIhPD69
KmTb+UcsRQyxcCIu1vo2buGAqdr+uJLlqpByST8q41IdJXFNibrnwlucVAwtHadmVMins5cEZKiD
UcxHwPUIK7SiHMWX/arb9fLDsAT+YneStsnK4pUPNwS+Uw6i3tCDfbu10W+Q/eaxQNExxSuKMQpo
1bxL3bhzmvRnqTRIRMV9W8DJP3dtZqCX7WXBV4VdgyQRtip29mE7olzt02xbeiZ/6XFAZEDEfOEI
JbPklK7XNnWB18XgamMhabMBf2bBF7z9yHErzaeTp9u8QEWz6TQ/H0o8/OxLi4F9kczvG4+UkDwo
4IJbdWA5fBf+SdJM/LE6E+NEBfd+T5jBsDUPkcvYmKjkTqOmRpRgziFxq5f3+hJxuCtxoCTOeNWV
7YnieAQwc9t+aBLx/DsgscHR4A5GVLlz1lCxgkuik/wTu+UcT9oKZ+agOFTx9ZxJVDq/DHmWZIBb
XdMp185QsI3q7qnNv058uqgui4rynyruI67ntunIFhv8XAsTeXH2cGrOfJGLarzQFROF6lP44z1O
xvtS+sCL58W9GZZVhMnFWYN7ZeoI2i+ZUA7ByxkXBldUtm31twcK7ZgAkhQH2zYwvX3guELYeTOD
8VQgJDhTenSDN2LWvdLNcVg7MNpKuoNdfEXljajWm1gJYc0MjCM0z2aApkxctoLkWroi7ipF32OU
K5ijRPGYyd7UOGQY4CTEwx7GOtqsk5trTfx7oEc7+YUPBf+ACKi23UDBOa0Nt+8+rgh7j3Ro/pfp
oB3Orty3X7GhCyNgWYhVmkPAOFqJVFuWaOGVAT2z9WJ7GwMip2jSndgqhlNOexR46NdwX/c7+0Xw
TGRozcRbsTyT2Sm2aGH4odB5MkEUPBlx7CX2SesgfPIqJGSNWToX7gfbP8x+X0EFxhUoqLsypA1I
uk4EhO1pk4qPeCYFmOauhv8TY6nsYGB1AlShRyx3iGYXHpBS6QKiBPi+BxE+YW7lpYnULT34WPiN
4pJgCnfTophLLlaiHGur+4/jzUOyXJSB7UhTBOsmR4dwnIhh/XM/K1gAUJnAIndtDJMBQxswncye
1S18TvetlukCJLxLmXm6fJocSxxoqe/qiy9zJ55Y/ejJ/u1B7I3K9T8sNpUOZRdRmt3aTzCDdjK7
R69+wt3EP+mVEHbQ6c1kpv5iUtmp4CUzG3vT82uJdUZNzzKQuaTeMOcF253fXKPg5vscC5v4dN13
mowIHT5rcjRhN9fNHzGjeowGZ9iy2Od6IikcI9av2AzeZZqz6DeBqQudOsY1Bo8JdPUblfAP/p/P
tHm65hMuF4xXCA0jt18XHKS7wUlWKSCEXoJl6L15b9i1h6r4G9BA+32c8cyWg5McUxCuEhDf+A7D
xpHNAng8WH1ltUnGwN2qW42MzxUn9dp5ZhiW6aMoIDWzIyEVLY/KL0MPSPI+99LyloCupK6uL6mp
PcNw1WR8TgXV0fSU8l5DSttR0/r/h7ToFv1Rw6aATY/1wPyFUeu8kByPgBF63Y95EEeBQrtFCfMO
hLPmoneHdZMDars9qmDRrQO0sIOHlq6N9Qpvqxm4iP7YDJjQ4FQNY8E6KPQ2L9QtNFggqQxG0MYy
IZyKJm3NTp9QNU3cXZp5kMjmJCot3dpDZFiEs2hdccF1sQWTr3CJKsN+iTEBygmfe+IdezYagAjM
zvjI2oR/68RdTUvQmK1Fw30hqJdfg39AVmK71WBxkGWips/ImGiyFmKaI0wg4k7YQf0vt+HUdwlS
eJKfkwHY/ibmCNM25mlcOh7fcs0nXsX1nqr7VPOW8/jEwh15KUY0TKUsXkh/f3jNFADwcRk9yKgX
yzu/RgXsfcP2365327ZzG1X4E3zuCNcwKAiMd73/XzgVQrApEki+DIAjyTuVgDqpBqvohxJNwA84
SpB0jmwyK1UamFAO3Q/RCcGXarzNoY/ppd7nQlDTLWb8vFku8hBefxiW6NYSOKhGq+6d8ufttYpD
/yBg8E7KYL3PnzYJHZTWuAEjSO6mr/j8rEMnUirUtC1OaRirp80FdLrnbZFlJFZMhcc7/ofCaHfF
BxQFsBxH53bw29vRcw2yrkbjpLUqpT0w0rE9PHOelfGtNEzYow/evRHXehxK3B+DVwXmRaVWl5l8
eY0CO0icjxXbTUMj5KfYy5DJ5Bbhv39MN93tp2WpMOf3GK3FnM7zkWhsI+G6IGB2uqRumfm10nN+
htA2mAjgnYJOSd9+iu2Au0HIrGwKI07Ru4T7uUb/HwKTFi+pnJFwRqR2nhXZtTWXWjQ2/k7Qn1sz
LRd1da4h+f9Sg3/TyTo4SFryB8DHZrbBGdgTnJtg/Tz++QPGTU1LAw1pJ7xUkot3cySvQ4yeOcZ4
Ux1few5MCzW+U+W3Br1jlOECk9P9aZjwK0LC1h7ebRCsQy4XEOYt1dezzKwKV87Fvm5+Ny/d0d0a
0zSoMPpul7lvNgDNc/9jNrperAKlZYgzM/sjajZcRqaWY9P3EiCtLfw2HxMc5VB5lIDQh/6fT9Fi
n0LNGKi7VUH5RTR14vXv/7g9D11kmEPFebdMDAGRmRTYo9eIyV5BVn8d2fRATTZOgJmpoo2/NvNX
ThRQ2ZTRgmm7y28nMcWGzEf6gD9T1fnYRNowAc4f2PMzWW1bgT8g+zDhfOindQ5w6Y123WPYwd2q
sK4cUfBS7PT77YMaFooMZV401fyKwOVvI0FmMUUE/yk6CFvaIRkuC+DS83w72dYLRzKi//zWIk2G
c5JY54+R1Eqok1zeigEKyio5XwIFKjKAVMlEgM70G7NglG805g6i40kFA6JcPpyZX5c7iNXgU3+H
RIppmRRNGk4FMZZuFHL/gxts6LiTZJdM7FzyF/ZhAus2d1y0b3t4hQsCHGVW8OCBYg/ubq5FgvoZ
+EVRUvEMbvrWDG1AvN7lm1sZemjXc5Wevm/Y2fC4EwPGRSSBrEhm9S56BZ7Y0LTsxxXRKL+L5DJ6
11xNZpZjHpY+C1cD3+h6y27HKRGbpMoOcFg1U4oE7fkruVkReGPOPFsdt3jddY4yCZ9EydOMIWNZ
H8qvQGIZnBgNxBux7e97pb/j/dMXl0tqYBZhrufN4qRBgYc/kTsxzLOSdx2rdlRb5EPT/2G2OG0V
FWkYU24WHu6Fy5r6q2yGmdiX2bCWJ9VnB2stF7A5p7IJ4sM1jUB9mCtaRclrT0aPXXZ1BPYveZFm
drxPzN5xBezMnfS6bbeU+IRI7oeO4gj+oROZw/CADjNGpPjs0lPSByINYG5qbCCcW3OUz6YOaIdb
L6bbSFCFNK0ySRF1Jeda9dYXVjCqgj9eMoKGrvEHYQV5ywD+wCyh/PgWYWSxeynQ9Zy1KIj2Baqk
Qtq+4dsvCDmhMwnZH+sYXqYyonRJr60pyitl+oVD2wNVnG9m3q5aHTpodt4pZyivMcwDuvkc7soz
6QM+3fcxPrQ/e3Ue/RyEOtfcxI2rfXZNIxI9QJT9EL3YoF8tpm/IEcvmc1RZBJOI8SCCTKXqFs+T
+6fX/zexJAUs6x266Q8PcD2yta1uYbqH9ONo6ycqtR3TXB1IHJHH4tBhhOaD2Cy50cpnWyDK74Zd
ovfuxokx0SBg+eDh7JIOKJNox/aFoKvobwuX2ebGu+qLwuUFID0ZLldaIOirpSIk3BFB7/iAhdfn
gnCfBInnax1PQKqBh3QBNeHE0LDvV1Md9yJ4c8wF/sa2o04BEFf5eWVPlZjIivNsPATkBkTjcwMC
FgCE7MEwzX53jlxwkb1AuskQYS3IpWDlJ5gguie7saF8AuqhBm2KCGMix2eP4puVybZvc1ULp6jf
FZ9JKFvRQmU/E6OW2NZAqLsnTzBuUkqw1QAgMXY3jWHF1OKU0fCcXzbOGw2LaMYCK0J6YCWnUeih
9/pfWUrJaf6x5NvCTqKGGdjlaqU35IKumWj8UtgXq4Q0ahVRhZN3xw0mvnPbCPzdXlNNXgPhVT11
lg/VgME6Eqwfj0pIlIm4IAEMnONPNvzsBiYOw4sAJdx9eCYwhLvLE5kujmYRa/45tASI/r2Vjb0H
G+SqwKtoly/UzOoO6FIOgUZiNmsHO1cC8h8t+TCpHZ7Hx/1BXF1LuQafGpOCj/7RHVwpXg9/yNVj
ErkezVNHMj13vKV6tlbvPjx0dw/a/WJBwirJA6XM+KWgRaRNk1ztynauJLlKetTFyEvwRKHWOZ4m
pNONEAbRlj+A4rjLXV2WlZXsX8sdqMEWNIR/tq22i+uuAR/q/NmHjX7K8F3HMTCXkZGNOIBtnaAd
hrtPu4Z73c2kNMB3QduliXcvHVGiIjQZ6LfkYiGzBaR3KMKP9gcVhvJAWDFOniAGbeKS+VOm3Qja
lrRvLQXQfRgiOc87KGpFg/x7uSZ0J0Ygj7+/sF7uxEkkJWoIHg0IaU3GCA8Kbs5qrQwCtC0PAhAW
5pR9BS4tMNNrxVRAmZd8g1TXY1fKjUziLc4ksbkrRen7BuRuH/cXhgJG1fo7gyvfffNZgHGmx9eL
2ild0/iTjcBE2h39Heh3/LQcdMrD2V7HC4OaBA6ckzpl2pAKVR62i49C7/H2nnKUxyY+IAlXC7QJ
yzHCnVkMOQ3IduzURt9fLWQajDn55g5c9mWBjlC6uRE9DCmN6SkvtGq9f2n0PVSPy4tqXnySqxQT
QRUIWyCzPKb/7bejhsCedIEUJDOrJIjWStHjXpiFoYpd2TBfellZqFNiDFN2RQkYvbizymvfJNoE
mOk31SN2VFl5lYAgQr/Zedvh3UxUs/O9z+KwvMIxHxndm+npZjj3N8RjzxXfoh7sHvaQIVP7GMHQ
MrjAhx6UyptI0DKPLFt+u5l/hTucBt2f3cwOVijpqMyQJI1+FaiZHy2qJ+K9aGXLMSxyyOBQ4ILX
JTaFeyx0jjzn+cAB+DkInn8grnHz8RpHP4gJoxk/XcbT4yBaOFN0bKH6zivAVw5bfSub13F7u13U
yhNQw3uyMkt5JDUKQ2q6SOMhDAEXJMHyfUCi1nXuqOg4SVFcyo324ou3ELMTdvUILxZZkpn8KuhL
7GM3KJstg6pZcHUjZ0WPd0r7bfMGODJoT3JeVP8DJXYodrKmZlQaTPQkZN+k2LcHVR6QGWSvDu5H
jWf77V/CKxsIzynPl1AbR5WBlxBk/HfVD8cSJwD63tNH+zzUbOhnZMrs38Ic1KePprMOG0cqDz8h
MspMyudLJ6l3QGuuHJucqL5G+dnnihTvaLptN2ksAS5wf3FgaL6+uRnuvfaGXJKLv4RbgnyQtIq9
o73GI4oAjIfrxhbT87Y4xmUpvDQVXMOIKfB9aCM7ovwMESkGgyczAOroD2ztA6jFNvdU97IHd5yh
Z7MHMmOYg6Dp6sWWIVSbEYDcKJgVd1jo91zCF4ZWxSmStdHlTngaCmoVaASJlvVdnWBxo6TvgkL8
Nq9DPJOkry7d7xNlS3cZivzjBe4ntp/fk/xghaa7qoLjCZ+DM852RvDQNjvh4LrXwQl7XKvVHKM6
fEK7xjTKa9fYTCYDJ7C1et0nVLfb6LeV961rfASqgEJ6o3HSxzMZEaWvErLj6+MfD/jnpBK4EeDN
c9HP3HpWU6RrtAO7hu0atCpFkycW4QoPVfMF+5C8eb7+B1q5VWMXldHo+hX7+l9stcKozxW5YqPa
lvRU0VlwBeThBA8x+F2ZramicKIbPkif8H/pnC3XyWE5ViQi75L0BQYGPZ697t//58UGVxUixKXv
ox9VFpf0fWuOp6vubPxuhaNmUIIBNVnQF+zTtMhJsmyhhbTSiMaT0TV2aVuh1wIcsg30406uyZ0u
Zvlkjtdb9LV1olvJ0r0gARl7TOGgLe7bxMK501yKn4YmX2vko1SVVU5HI28bCxzB8Ktju8DWLomq
wb5apvwFKf6tySYg942SVpzeQUA31y0DM1/+aSmHohtgQ2YO+T9WzM24so9I1Z1ZSWxfEMWC2duz
LtZQ2htZHk/jlyoIqJfuwsjymRuGfq4stgkjBSjSjqTAv/WZC/WQ/Do2OECuwIwmQ6jwE/Oq3YQa
A74vua7BwQwOHaiBdSUlmZsTg4mV9nRltY9kB4ckfFaBbWrzSXTOvrtFLzoSoEyLiWUzW337/YgV
bBgmdXbTUErr97QnbRGD0IR6XsJhDFYGpTXLDFktzKjmOInqtB/v5klKsQmbOnbPpDJCj0DF3K7O
HOtHl/0oCFWx60GbDdzjHayXfiumxQapyL8pmspm0x99Tz2M2BoavyWeLD20+GR1sSBMm3vTUOWc
MKV+IGXhV7L5obJ0kj/Ohhfz3bsohO17yDjkZL/2CQn/RLuSnDiVdvAhHGrKqZOOBpJnlxEyY5ZE
RYf2DcleESyRUkgQyyMll9euPyHEsn1E0CArwTyRucehod5HPK+gvKELxSCq2V3hGcWgIOEmTsyb
FnF/ej068AGcdbCXhXR8p81hnU6MJ11uZ/cojKlkKnj2QpemYRkrvxxs7K8UJ/qjnsqDw85RYHIB
b5OgX7UiWc/uHeWixt/7o1P2sKsBaQIsnuWhBk5qAdq5Fag1F+/rvKgIrgfNLkTb2P1S5DhzpUK6
Jt16W2PyMUbkAK8w7rYqMqkTOoTnvEK8byj6SqoQXqUXvwQp5ZcaHTfw7H/PusdnU38IdBOuZ9ZD
Wb9Wmmh0PEbsYtQRmbZLIkT6kErIyuNBlUZeLNG5LkLymDRmkXqbYUI+w4WfQ6Q1xRvRNPUPpGzz
ZrpPKuCC/xTLotvcJ5wp28xFxTNZIim7fX+SYQCQzmNvm+21Y/N4IRBWShM1j3ITbFsZ9eL4Hobe
tKa7RsJvRcSInGCVBARdp75DittoGye9dDtd65KX6zzlJ3gAFdkSEC/KJ+JRZOWbBXGifbNd61B6
lQuZ5SRsORRi6ef60VRPEi3EvVVC5/sMh6QdSj/IZH/ch/k0mWMGQjGtN3QOEC9fhyhGWRv4GiDn
R+1873zLbSvu4hWRD4jrUoaWdy3JusfCtURn37z9pjaFPmefVUQLVX5qpyx6ZzfCQ04gCNdAiEyG
5keRjHQc9Z9Guqvbggk4jkP46OJHjqPQKlUFbHcN3IjpVecEVgxvMlq/yJFTofa0b7Zvi4uispFO
mH0fnpEgp9L4HI+QQfqRZ+Onk3U7Z62mfomfl60xbHgX1bVQ8wVbtuRYc2qfWI/a1gtRXQGQjrPg
rgUbTOBExrYKIwBySXRqQX+b4LWsOskgjTC5eY/U8TB+q8D5oSbl1xk7q/O/0AxDqAlQxzaqgxHx
+KEr5f2cwBBczC9QVY+C32izJsafHffMUj1OH+Dtc80CMD/cA4KqoNmUBmc0DStuYIqSaetK+IUK
YZ9jVHWJ0iWuEMsjXa8RotAd79lqEIR6YWux+IYRH33icbGtDWnvYj0oo9YTeKThrwJ33bb1Dc+i
6MqWMkpX+F3qLAe/YXB32QXeGEDN29+9laeFmUMuWvoTzHV3dY/QXHIeG6YSM8/Z6BStqn7wFagt
0k4/0xshZGcXHq3erUZrcte1vdotfcIWumRL/HunmqRTjaqnSZ5d0eFO8yyCYnP/VvzkJBGekc4X
ZbBako3Bg8Zx4oJnPPa9iTvn+eY2qaJJqMxnE6uodkv8/1ZabxOWA0pHaerdMJdIrY365sXltxbM
wf6aiA7v2mo0drQGK2oqgvBWS6+lg8QEbPUIERFpT+2JR/k0OUaMJ66qIte6qh+OiWZGBvj8HBVk
KQKtJabOqve/xn8sdkhbXw+o3fZKbMk6Yp4aGjrxv03QubB7uWDLPjReBwPJUPwvUEuZI6TCixx+
ShGsYhejlOflMCUeGD+kLK7rKVc9wR0qpez4VjrRVH0yhNu4MzP5lgiANP0woR/FxvnSJY78Kwzg
5on3CzPcxr3OnGSA5pzq+Jo3hoMGs/FPkhA+nNicco8oh2T9W/TD22wSkuNd9DEWz/KfPS5cwhty
YYxBgEMl7Y4zNbNt4pfrTKa1HvZnwp2OgUFT9eKGFYlGTQwAq9+ORqZ7LH/Evt35F7BT9AoW7FD4
dDBSl+onYhaxKBAuAWGXGNczt4+Z5o7qYrPTC+iGPBJICy6rxLDpILBhDqP6PEpN48iO2OYShAIM
r1zdFE/guKjgcOUIoo5sTlFH9V/QvP93ty+P+NmSlUpYRJSTAuumedcfFSivOw7lnGsBbwLVF2LN
vKoKcFnx4bgmSBdkxHQ3sG1RJTEULm8I576RCjPPMLKY8kTjGxxjRoUkHkyFI5cw7L0dJ1ioTMxX
TF0Dhm/smySerq3ko1r440VcTNY+D61l9D92ZpIGu1sXCJn3GVRNJp9Y3zpM9GiyNhS+Re9B5N05
TNRFCxL7Qi9qBEnc4GaaXf6UJQCYK5n9KxTojyeI08GwlmIXygGOGkqdB1KoPnNaQPcLorFJhyqw
V1YfG2grHIBE4PmpqCJ3nICZRqR3b+NtP9SmJvSU574hvxzZIPZ2W7i7EV47WjXAQFaUodIzw9V0
0KBr1vqlmAJMJfr7uoIY6XwH+h2SZjdDBXZB0U4XuecPYXs+bL5h8lV4TjQ7m49R5TN9kbXYcIxW
adMnupLuw9mGJ+y6DBp7FQRuKtnki6nCpiWDbS80G/EhjOBiVim9ixKC1au7hUZOUt88ss4o+LLf
KoBfcULHmxbQNJLXjK/Spo+0J6OY+ZKcddfZVwMiafNn3/iGsSIeO9ubdR1ORZ0r14DXg0/Hjp3f
X7qjKEtpPlHUE23idSIgG+3EjQRtS50Ps+RwwEqdWEFcBsIu65Ri5Tzw+Yc7BcLAN7UY82Au6tDm
RHE2jnQcho1xrp0djIPhiybKBwdhMmvoVngERQcemLxZlpAvlQ6T9w/ZjA/Et15O8+RDcZAYnRrw
dNzIDtRkpKDXqyH+Za8mSCJaUpbY4hoeWOV7Al8dH/xAVuFszEhfD8c/eEUXW2wcJ9wgpSA7/y1u
bHVdG1AKZEwSl9SKEyULPy+IzOHLeQGfGPnQ6xtnAUzn+ApaPO+9lvK0r1iNmt5H47PzWmb1EU+K
t4vxZTBV/bKKsm1gfY9OXJg7P/8WjwsLQHEk3cEYb8TR8fpqWyt6IN4EPvfrywsibQoYrUoRL075
TxkFFuPWWBrYwowfFNY7ycbiR/sH1kV2ehDnKt+vOW4sL0sv9IpUmz3kFWIZZY5u+4LD6u4We2k/
CSJOHCDYkBHDFNjpLSpv5Wok8MWjIpXzI32A8qaj2IONktA3rS5uCBsbey0NfXGyNalzc+aFlRDx
VijVV1JapobLthKeg81SHAvlxJXWzAlOdyi8FPISXZ+7L0sA3hfkRJ9Bmr+j8f6c387gcUypimmL
MS/1IXSlUe9gaq+pliqXYri8tv+5CiIYfPO6TbKYR13FCiUE8FeVTjpPfK++FURR1GzJzCx7It78
GD1zR5+N0F0Ys8ocR47WiODlw4PusWCPqxTF3LDMTi/qFSESrf1GcsQZiuhi+kfVY8Za0wfX5mxD
um5xshihDaCuQRK7bN6T55LywEAq5TlxTbTDgR875/8fJzApM7IGBp8yBItmI2LIAm/JXmwKmcQe
bPMy2Zid5ryovpZvDiw5A/vePAAdHeImXC658kDrOLbTQI5O/8HOkiRDLKkYtFoo8rJPg16f31P1
vwjp1sByHOv/NevSd5c1PwqWxLHil2wzYuI1W6pG8mnSFKBOabyLEtY/AzjozrlxbO7bJPtTwM+9
yiZmyJHmn0Hy6kDYlmWAshVgCcoHXIarxjgjvjz+89M1MMBsM0Wih/vX4BzdRub1RsxDuQmrfv9D
15bAq94/wPIH8f9cs4YsFPySxRYgatbT9IgdUNY5iTKRAGSY4b2ELNVo2mH8nzwtlPC4Xxn4rI4R
B+vE5G5bMedNh6Lzgv8z5WVDMgE4P9ez8tgfFTHKcJyU63Yzcj64vS41bdcyJ8WmTQqowyOjLAKi
52G1drxmxl7YJcF84i2Tx611rSd6InD97emv4JxixTuZlZEh0lBtpwqr9ulbxApvj/vpLbQFG6Aa
tMhGyr1tzBTeyGQ4xKMKz1oc9p8QBsv5K8nMUqt39LQfK2NNwRjIsle1fQwuDtxW8o+s4X/rrtBF
U5iqWoUlEgkU7DA0fh/HtlYa90h1Go3gD59D+WXgr+tcWsY/DOxZuAm0r+CCXMJPPxsZJPcKUStS
M4mmoWP1L65POlpyd7uo5WexyqTOdS/MkQQPPnD2HO4FVZF95ikZknoMuywB1bGr98ui5CzhlA0j
EFn9ctO4mmjceK9tFjyVdpz4AjeVF/+Ht8PiozJ/tOU99NjK0Z5zN5hw3+TnNm3b+hl4v2jP+NLA
ok6YSa5hAi3q4ycgFZFdA/w3ebLImza68QLSwx5tw02y3KjsDXwqnVJK0/eXpkEWbQ/qHqyeExSb
BLbWviudhI94YLx0N6v50ESVQySeKibASe9cYDA3w/Y5x+ZIBqPYT/HgzU8k//+1Ds3LajZlPptH
cXYfaShFOylDzr3QyLtYm1ox0zZirCikffYqsWyU3ryyfG9pEB503cc06FHGFPhK0nRIl71eb92x
Kgb2WlPRq6klgEk6cl+SkCNN2u0PPUeVplDlYB6y8XACzhzHPyWp6sg0eghM49rc37je2ZNW7ghn
ZTZunYrdKwenZxqDe2DZuhdUnuFXOHm98m2GEtAbbF+C/MzEUNeyyj9BXGs0QMJm+I7t93n1iVXG
sCxXCjJs/lFzZss09mf+SoV81bQ3w2muoYsRWjIr+PwkpwaYRwUGXp66dO8+2PeOADiqReBjj/1s
EtPO0I1dX5q+LCz7ULGAjvW35CK33vziWY8lARQzw1s+shLo+dfYMlOfTfxsjV3jgEnjVplOUmrV
EEP6Uv+WLAIppvZaN5c5tUU2crGm2m3BXshG/puMslLiADdVonHPscQPbW6gwwZJofmKbHX/barL
FbHG5TSC+q2v0rCtKQQC1c4UNuCbBiLDA/1+QEHQFPxLKui8MNOcCJF6kZzkQLa4AV3brkOEHTXt
sVCnIXeDkLlXYdI/PCbxHYs2PjSukEXnhhEKR8+Z18n95cKTEPD05A9b/nbD2bntX/YZi8QTaRa6
IZApPO1hek62kc7qbJyrIQwA+amNs7BH21vzD1+O1cAPVOiNFM6RpuP54EPJnPrzvSiOLAlcrcPa
uzRje3UKHq1URoOPGuQNlUJD/MaUC/qRV3SBDJg9WXS0l2pmnsiubL++W/eFMj5d35aXA0rwT7d1
GUzBzqbZgGQuhR/sizdI1r85PJwI+QD1TFr0id+diA4HXe2s96vShp0hWB8rkKpXv3P40zQJffp6
pPjgxMYl1dlXrNSzCMnScgh14K3VOewt2xlM8FG05j0D7zGAh886apyhwK27o1CQZWqKGn8THheV
c9cx11TWYnDRTSK9k0LrCDoI2IhRzeNe4m+KArHcHtQ4NUqtFVrfXFhLkh6rSh89q96If915ot6I
lMd4pZGHXrNZ/KoivFhjhtKAcfBswLJr79QTKoVeycl/oysI7ahGZTCIxPY2nJv3lz4qDUiEoPv2
jxGwOLwx5Z4ivRFLo8NdDHTZ0lB6YaS96UcEcQIVz8urth1PeDLOXs4XkCugFuAFD/qMZXFyRpNr
7BW/gKlNpqNHoNfvUknaOSCKba8WxmJE3cXtHLF+D4WuBf9Hcn0Ao6Po9BW/+EROau6EwK5GDTna
rAkvZeSCOUzar5YlSaihtlkg1nfL+dzQIA4OGVxGj7zWQPNGahNXceDMRGMNQBESG7htVnr68546
XsN1uBfNVgYD//CL/uewNSDjUrD+b2oR57IS+hPsq/7lPg3GTPb5UbG96xj2yzHQtVruRlgA26V8
LopsYe5XaJHMRBHDIPEwgUoQAypmERPw0wZTrs+nExUOGYYBF4DjRwt5aYQBoNh0za4mYuJWHHR7
gqv0r/rIjI3NA/m9mKgI6kNNbhc02f2rjnq/jG2T2k7GLNKqg+u5oMaRmo+gjutAT2jJoJTzmcBO
MxLl8wwXgjFOXLp1i2pRkfJ9r9e5K6JLFY5Q/YOkCQjyMCd0l6Efx7OBWRhUfNgCgIM5MZWhIZF1
PbXPwlViRbe6YkxH3iuKSWCU/dtYlW8N78JdCwjSOeQvWtcRaf5+O9wtrOnbYs+qHyzfjzBbW4fZ
N4Wkwtnqcc+Hwdf0Ntj+5hJlJiKyZy8WhmzjbBGUjWqyvEJPfzyjZNhpWdQ8dVN44WO2nmDkDQJ6
8an1pR43eo6EcfUxO63iPhb0d6uxS2EZLZQXa0br8W1QI/yyVWXELAPFV7xLfmcIiihCBEu7NKJr
JEAQNWoKi73+rPvRZp9WuskIhr8xdVrFXKiO4Is/QzXUVdMbifrt8uZGwZL9EgFVKIASL/BhX/hx
pJyzq7b03YHVTGrHh/hIpalU8oOTyHgJLINitJglMACiqbWtrWPOuo+xdUSWm/iikqq3vsRexQU6
+VsoJ86h3Aq2WcuG7Sjkvo0EVZ/DoUHIuKUkliVrIgLW1Ovq8brKrJiWMboE2SlXEtU2dZhC4aoC
ZBiBRKw6tza99VIyetClCvhRhtI60eLvW8KAvysUB05BAq9jx22ixXsLYM4H91W/nJPG9egV7Z2O
cFxUqyN1C6y5YPvY5/7Qq1Fw9agL6NLmIJBmfaWI6ZovN/6QGylg6hR6ZTwoIcF09bCj+Ym/WHjM
MXdKM5GOMd44fL/cweAV68ZjKRvvKhl5DA8p7F2RV5+lEkb1CYaj7Ul23ehPXkwNwoqNcZjyV83s
0HYl7/bpt5LdGzr3OyiJTa+OvdBpTpZytJNZB6xTvgUU1yyAw4ZlG3dBFyAD7S7sXohFYYyYX1Df
d/Pu4C4bexghjji1jEs856gJohX2TtDe3XuAPJgzJoWkFvpEXkM6PG990SNSuQf3+o+7hp3006So
+FsBCJSJ5BbpaADPWDy652q9U1b55fWTVk/ih4Wt3WNtgwJLApQo5dHfsYC9tYDHdPqMu5JvdLAW
2O7+TJnVZ0lxhFkq5PcDvNZVQFROStWPR8zxYicU2nZp31q6p5VxhO7EEoXrOskvFxarKkQl6UCM
/InahYyxqVIJfD7PU3Q67iF0dmJrGNJrjWGeLL6ApVuflgSoU9TqCTEZuHpGUHJiyQIa06yD5SwZ
9iqViBYnDrIq0xeBjLVEeiZyuTfwbgYZySecHJlIyupGfWD9NhW//CaUMPlz4DVyYV6kkTqqWLxG
ogcllmzZiYmVYDESCogXgLLQnGSmYupBuiVH7LN7mc91S9w2OxXnrvud4GSwckAoN+IPsbEBO48s
q1uPuK52/38KkGvZJ3JUJ/Cm6ABKGFX8lZQQc+AAXM7NZvdJmqKel6/fWNa88oekaTP8XpYHtYEx
KohdtFRpyrDT0gbLMPKsjb4jKK0dBAX/orJ3TFZ8OYspN05elM9zOZs8+CA/j7xGH+7wmWVfatG7
FNvULR9gpqo2wgn1NAn0k5JaezNejbIE0ZDMdmUQy7qGpmc8Li3/guUw3Hles81EL1cU4vm6qatZ
xjdPTvzcvgMmobYx5ZYM5e8YTTDCPERMSkVivkoupLg4tmaxufbPlaXq8+JBkh4EGWO71vCdNfWg
NEKq3ur3nRNVWIsWe/ttY2k1InN60Ia5Pos3LdoHx0JqmNmJR4+90eiWoIyd5cQeeP+sKVunbNPH
V71G3ifCp8Ym1FbIxquWmqzyWbasyKmm59Evn2KAQS66dfke2pHjxZ4YoPrQESuhB4/UhLDKiQdK
ZR5ytBXX2rRytKnlc3DMfUU6qMO6/I1CrdA6urNKUfRBS70URWEsk1J4Fxh8Li2lWQ3Z99xhVmpr
r6Twc5z55+SUm2BaqLyGEEYoy77NCksfmYlOJfwpI9eqCaY8cJ5zxkQIRFMnjlndSN2WKdZqX+0u
FbjlGaFzXF53Mc5gHOL6PP3JrGcNXXxtThticBpgPtzl2TFfhDlkjdoW5bItIlIKmD0fzlFInNFY
yKLeZnuARU9ECSqxpMka89JrIJKv3pFxWrzB4N4PVculOEPjjgNEIVhqN7sAdAmaX0XFfixPDXis
VME2Ts1WjJkEDIcmIznZE7T1kJMDrUdnT0lojQnsfZSNYvh6PFUFh9MdXc1x04Fz/P+mLDvye1zL
UCsRRRMJ81SDM0G65LaGUnB6vgLWu6sH6G79oVCcMv6Bas/ONBfGvQQlQ2mronsQflospYS0l+0b
mt5qBPcp3Teo4cSPT6IFei8Xkk0CiLYoKJD9E+DWQ9sinWq/uecxYAS8ZqygZIiQVtjM9N2pt9Ie
AwP6NEh4N3/JeqdixdiQk/drC3HZW3M4Gk93xzCdXyJkQpU33YV5U4Hdx3UiSN8t8+O476dcA+in
X/K9BrX52StXS6nAhoF4QvAzOncNQs4JrD7iocP5FpFttIEJghr1gGpMiHdjlHsOhJ5dPa1mk/mk
nofJ9cpiFY9iNtXGNTvYZWvYjhVqaacGNCSnizb8gFLzBWcxmoUl/bs7JpEZEBwgZSDMYz7bbU4M
5hWW87fLpFdGuped8af9FpAEKHreXBzbBSpu2Pe36u68gnTZxvfOxlzVXqQPAZNqQVzVGZfZ6tJb
/yD7g1jEFfgm40MSr+GG7ZV3y02VA2xCPWv8nCNfw2b8DnbXj+E6TT5/7O2ist0hAd1q6T/qgaoK
YZbNnmmd5HnqDQ7W8CWDdOCxtPAwEAXUbTURMrlTcPEuyqUbFvFvB4k1mT2uA7rx3I6++1LPOlCA
zg8oqqgohh6vSdXBDqPMhHTQUuklDL0VqI6IhBfUcDoKU8Vipjz5ylNkDhZvnhcIWYj8eAh72Bkx
j3h7VKhvDMB4nCJCcqz32Wgfg7OtgGWOP/FZWRMqbyqxN0HeiWnM8Kz0gYTU+0zvtkZvFCslVHvr
80UV4gVniwrg13hW53x0DJG2mqnWgKjOByVru+ElnP4MiBYWRnlyOkNxzEfM2T8zU20Czz0OFl2/
SHuejLumH6j9nMiP2i4e5k+bAn9qXOcsIII4c0IWlTSekI/1D7OK2FxgDfJiWkoCZII3EUcBQBOM
P+3dhZ/M8r3HifmKN+VrLwZT+d4dWn148CAilTPJvDwH02/FQXFnA6dZgsxgw/6JZUQwECOCVUM4
PIde9abjt2OeL5pL5Jh9pD2qhQfRRlEw8hXWRAZsLo6KmXcG/NRQ3zCV7qLXad8fAbuq1rAEwOh/
qzcX7sTTCBGWRieY8SpkzbLivyPO9jd2lhzessATKhKOFG+Tn3a8JvLBwa0gPCEn61/gklX+sfVP
HfcGh2n0clByCrEDEJnGHgUiiRUFTJzpmHUg9qkDsJkFmXbMwUZFjmsmw7/F1n4wztzcUzWGmMFg
Y8IhqVMQQ1/RNaVNx1sVvutd7ILqXWGbkHOq5Xvw9+3102Th3vZED2D9pJxiW9Hpl1nojm0qCJHz
MZ71o9E5YJE4bwggv39xDCT1T5lxKPsh9XCSxJV3b7cB8Kt0KpigMY5TfInYoY7NxZmNTrVvZ6J2
BO0OXwk5iXoo79XdF/DaRcWEd8Lezr/cj0R8gaVOHZbr21rkJ/lZf1oYESmQIfYox3arFFLu0MNp
ZcS/hAZXCPFx6mUU9AcLtsl8BDZ41rDoMOb2SGCxpBOwJOF/y9xvg1k5O+u2NH0OPJWPfvb+QALm
T4aNvXMH/rayQtWyiEss32zOX6KnsYgSJJXaOnu1YhzBZ/ru23piRmXw6Vr7aSnvs11FMay7F5eN
PsgyqpdabD4HqrDJyvHFUqIq7p328bY7Q/xRBK1qriRcTSgRQYAQ1zLE252xUb/RX/5fW+M1BV/l
rSTzA8nstBxpU9W5UChBfhBNpTU8NCbPZEFr4Y80cxCtWLbvY3EL9RjUk7uuYpCJhlAkCkkk2VDk
FDFqEekd2Jz+lSTRetZVScEHUEdaN9UdRVNGIMSRrhQtAndjhEiUjXngTxpTEa2idSGHYDxzkUyC
RIh6cGWi5JxJZD7luDw6Lbj5d2cWSNJgsDwW+uPQyOkJMM4G7VoDBfszCo2YZPK6DC6Tt8lSu+qb
y8Px0DSBOL0FI9GpQLEEqBUk19YMmnnF+uQYeGKGSqwXDhOQ3lgIgFat0oxfpAsgLqVbTCvA9g3V
dA3j7aGSb+j2vjPCwcoVLqG4hRQvdKprrzIt6WMw4M6qF6etjX4zKz0OR3zbiupeQ3BPUQprsZva
mqIn26Og0NfFend0KIN2k9v3Av3cf0+hIf52b4xTRYjTlQ8vC8xY8HvAz6e3aEneYHUgDVJlkiBw
I4/Xb3inKxbU3+oJAWgqh++vhp6k/p4bw7DBpCHYXUb2VtQeZHaTxcbFxvJOCX5CMjkp0JsIjHS7
IdfuYJU3WvR20OYCKkgJZr8pBeywjaY7DVWnWW3vPZ4UbsVlJKTTdrozqqXNF8iMT+R/RGHSVAaj
10ZhahGozGuCI5RrvhjCeZR8OPzF0at9feo8WGEAU4uf4l8zBdvUScTQiiz2fsZpyk4h/5v7888H
kIf52RMjA7n6pe2l2AoLbEwMW5iJeG/qna7NlVCev+wNkaMuC61oTyYvIOC3OF4ATyIpBfZ+ARfS
DTc0pAcxHOxuGa09lUGD25FbdZFexMTkiv+lr/wYgTKvt1GVNh1IoAN7+1yPPQFVUfOcB6utQ1n5
pVA94GFlaAawxhnEjsMyzLtSKagdyx/knjptV8sgVi8jrexM8qCZXPtQpO8Biv1QWJ7afJ5mZiqi
YKUdu+pdbnZCrTnxCv7eRl85QM28c6Wh4HDMdsuvWHZHKSyYo50tQWYDD+gBHdAtmhd1k/1gvGWp
sSL/WXSKLocV3+t82cGu85N/vk7JXm086Niegdzy4FMlxIHtzUhIotUrB4/CM+D6V7i6meGGsOCB
rqJSOO5yB0vVrnXcYsbjnTq6f0gk7WSSZAeDOUdNiEkkW0JDT7GyHbWEpyxL5kyuFt/wysSE8o07
E/8TmMYoZz0qspGnD1IjhzE4wONWDUpNpa49zk0y1dHD2bKfKLZDe0Vci4nxzjaRPEL48EVtdI8B
p/yr9IIPp5F434hq5rvBFkXzASUAZRK7CW4EIqXTLg/xYqPlO45SwcIjhKeAnmXTJbg9sFWzMFAo
NkZEsR09sn/hGhuN+s+lfNrKuZbtDtaw0goxPWB4X4tDTH8Haehr3mzyDzJlxPFsouCdTO6f8JRh
BOXTK3AxEkPAZ8x861U+SEGDvgfZAJ+qy/wRIH1ExM2HxRD+tw7Ux2qL/yrk3aejLa/BScvfd0r3
5QHu2gc0Jn9l0GLMaQRZ2yYxciWMiWKPhBMHcMl7KMVBMsL1dKSdDFvfs7Agzyg/tl+QxB/rMW7g
03UfgNE9OQR7DOClUNRt07jQp/o+R1E/50mm7TrYUeHSEhLwo+bRtqL+9G5Krfi7JxMlOLkfvith
0HkhHR2F495OIb2WQ8d05IAAydIjGyyRIQPhTqhfmPN+8PTF4fEOsuAHM/FnnWNpl2JDwl4M7sg+
sWHVmoEWrLa73E4YL5T5H6YL7xh3wyYPBHidkYvJPqKqeYV9SP1IYG7eW6I7/bmvUURb70W7u371
e4ZUcaOVMK4ukgf1eyINl0C6bdRb1pNvZlA6pspf+Drgbv0+B8MMtCPWacI7L+pzpzisPLwk9ZQK
iuvUmihZt9R7eqqOVXLlmLkuDfj33hl8pdgH1p7VtBKPLBssrxENFvr6mobdAMgDFeaRjfAKyDAf
E9sm28bFp024+FXQHRfWSWVr1eEiNXC7xkH+LXdV5/1nRhq37M9PNhdwBSqDKZXRdO+tRGceDTEy
tpDsxa7+qBpQqlUG+qOhDSSVT9PGfhsDJGMxWivwWHFS7B+QDHdcQscPGrBSJbjdeYYqysnpx936
lAJKkClI3xovKJmS3wlf9nxCZ+4L8ac+RPNElW5JmIF6IzyHiPbp83qZatde4KlsOVMZsjDnZHnx
iDZ8OvxoQPrzwRd21i0ql/hzZJdYXBW9fKduScjGrjJpcOxtVcFkfvICbd3vS3p8i90oHMar+WM+
2uS21JjxBK32oACF2w/9LWJG54zKcvVnXczgLy12E2TpgBh+D/q1gH4RMagyNUHiyy6LK4UPUNr/
Zu7apy/4Xm+0a0o6j0fQxOR+rPyPFKTCml3fJXC9AqklNJJD86E8A/vdb/4LvQl2rsJxcDGsk7oY
RyXlm6ov5J4hH30YSU5LRvWl4dwdTz0oXWU+O27EC0aAdDLlJp38LoF4glzZn6136F5A9UKjjDMz
tExGuxSSap5ppvVMtC1E9AKdTUk021hp9Wv/TucDMNye1x+EEXeucg8KXEah2NSTGg35T3XRWS6k
G8JWkp0iYurOxPc8GK0dd6AIxR4E7reLq///8WPbYERiUOw8+cH3ZbuHOtOnHkIVXTmX3PIkH/b0
oV9UTWtLkiQMAZJiVOrqjohMxDOWXufn9cUotMsmwiJB8pKa64R/t7rRtHS5bt4xPg4GFHSGYzxa
dQGVWAnO0MFM+N0dEl5o02tECu2MHx36iwCzsousVax8fFdWAiVGj+dDdUR3JnQIRRY7eeABcutm
o19aJ0Y7uGaNvxqeWjGVtMlvFNr9/tymqYzhd1ydMoc8lsKnOOpNV57IsTDkM1QmB/LTBoXp2g2H
FE1BZ2mMyT+zfWQLktykLRc57f3+79YJRhYxCQykOxEt+aym9a8DiCiZ623Dj91SvadD8az7Nxy+
zU8JMF22MwWqX6XzPg7KrD0/nyi5zA8Vl1NQnq0EcEplYdmqdlZl1ggz5FsflL8f0Io8UPjQbpEP
Ug/1xumUBMC/dqZhffjyL9AwOoap1MtUM9UdIZ29dyRritFul86ZjkJGAst63cZ8YQRwT8Rt28ws
DNR75tk3KyiXFl9FlgWDo5VRiT8x6YAasjuzZbvP2cDgINYchND8qQ98/WCGPDeJnnn35DTmcrGi
58dqM9e49VzIhp2f7U5o+EJEz7UtGnCA9YxTRVmdGzXrrjc/yCiE9Ex8nW1skLHGK+hrzV0MNh9S
iowmZp2vXtK/HVFjU4/Xd/6JC4+Tu9yBwpjs0nfdb2cyUWVwqI237nenVlGwEY9DXBWNQzBk3UaH
pBvZUDqIKfgaC95Sus/t8Kk4aoNJQ6obe+IgQ85LLW2HKTm5ll+BCEjQzyZxZPogZN7N/v52WiJn
6n3o5nVmtNEHDrB0QFSIII0W7jh+Sks1htofpvO+8tMeKQmYRym+IdMGXL/Iugk8au4fuGG+U82W
OGRUbHtCgqMoOyAjmB5QOX+GVR3QTvXmYjSES1PvYgVyc7Vcgw/hBSSzmXpkMmO59mo/J7x0DvgB
HjpBlQ6DcCD7Me+6zIFfuHmhnoTWnvyyDMadmnw+ZR5fUjfRwRikd5A6ZOZPzhUeRbTv29Qp8gsK
wKMgHtGSxrmWQJxkO+awv27mkBP192HzZL34AAWZPHKcAb4YsG55yzlXAn9pjcQTFD9ICGcQryF2
3uKQXUw8nc69kO5PubYK6pLI2r7ApwIGGXklgIbnPNSJ34qWnCFdDWJ2p0xCt+BwRjYUhSP5uF2g
PfpV79y3cStbo7M+/m4vAL4CQI1IaduYKjoJ6lawe0FTvz1be5pNi6AxzVs5tb+XQMzdrscQURJn
U22cdJw61Iq5/uBhIEeGHhVEkyKWv8A40YgvbXeP0p42zkkPFY3rumTR/WcvNz0MgXMZzfPLf5WX
waoy0ropZHeYfkudV/SQocKkTmKMevIh8lvRWIhiNIyiJjXlI4Tks9Fcxnf25BZwVZgh+4NDNQVs
Bi5LZ4iADmMUTduRSDyc3yPudOsK95fkVgeQjdF8Ctw8RVj3FTBQgOuOExlPI+hfxsrW52cEeiAX
5KTDRwkXP45rsAoLU15njC9FZrYtVqeSOTA82yjAixXkS6jNefrhC0Q3RdxDJixfbaa7v32yeK8Y
pyteMwdegO/1pQGiiKvktW4JngIZnsKFyOmZKv1nLZYTcMM19YGgJ/Ofg3VhZcOXehM50IpX6UlY
MGOdhezluTYoo5JaAz+r7I5ZJUm4skHtqj+vuYNHmj5nTvWYkdgUJysg8A6GPFiZCoQU2FBaCl+S
5O/23N8yZSXLuDzKJ5mkXDhXaG/FD+DlQqHCSLkOjB6bjq0iq0KBuf4g/PG07DWA1mMxoBZVwe1E
BNKYvsxgRYOkpgd86+pb5dsOmNWk/EgT4BgdDI4k6kJ0Qdl/CvlbjpcRAg/ObexsRPrWJYdtXjwl
oVXlqb7lvqUjq7rLSS7U3rJIBWdv8Bow0Hlrs5NphZ3CeF04YGIYG8PxC9ZmYxcr1pKpA7r5UmlM
hsAqzojB//T/FRPfDfjwYu90s2CaA/LwM+ANpfdtmGYrwOYuQFVYmaBuRnVYk+OewiRhxrDWn2FP
cefB7VNfJ223lCjGIqsYsOzyzx4/IgZ8Fc6AYJRLTbGH1LgiBB7fRLz+50lPAA9cxc5BiabIqjKs
zpBptZMSMlBUmYSbw6Bm5dsanHpXnxp4GRj1T9z3P/S7tn2c5qiBhLthw81fk/0U/e46bUXkwhAH
VfQJJz3dlASae35IqYMA/J/zmGn/01Z27ATclNSAEbp3c0oTGt+fOuCYvG7Iu/eGhn1gWWk2UWbo
KUp6+7GtGr7QykCOC5IdYYLQCSP0m+d9D3z4UGE1pML+CAGPRl2pcl2lokYfz40yZ+3bqKmLBv2E
8S1h/IHRQBVdXh29kgEr3XwveSeh910Eh59WlW6+sMg1c7804+p1i5CNZ8OnP3fm1hbxQvzw1BHc
LQOQkvgsQmncpnU78tPS9AuBwlsncVAjpfp9Swph7DwWK7USm5OxwcEJ7XnghiH/fokpec9o5yPr
BuFIs71m2CupU2eH7Zh1b+FLAwESAnUy770JmstTajCHJmkRgn3vnbPgpC273oPsp8Gxl1uqbVS5
vR356tLFbgfFbPbBqeoO1ioPYp5hTcHCw6WGZ0kS3Rog/YM4HJOGzpsRUZZ2hfK18YURWhnEQxDc
S/OpJOHHKVd9I6qkfY6B18xo3Mel/OSwwInRfM6cR5CQOj3D0OISzyupZJhDqqHRcRgqrLsKaJg7
aC3S+NxMk6kFBYf1SaemvnZrgrYBaJpUR5TqHa8EDZ9ZLvNir08L961emyYJbblEsxgq2W8x5cM9
+IJVEMsMK4oitPlm+ljXE/mIV6o36O0I6MyrK+hdyktm8OR/TUEAUpMd3qzfti09YIwUqfMTS5KE
DsQF4LFo2G4JLHrFpm7vWeNFYBrWKnXaGJ1ZqjYQxdgzGZxxGrfPsWg0n9zMSicXOuqPE9Do0b+o
zLcjjRgtQb6gP8UeqtGyzjT8q2FoHo83EB3pggmITPU1pbh3wQZor0IguDBHV3r0Bl6BG1dtWJ23
4Ru2sLgZXGVlGkTzBY+47xzmf4x1VPbG0JmMqkwUruVKeoiLmHOgbh1j+N+ou2lIeUzM8cYbmpTH
xvMyr70xYGeYLuKvmSv8eJvp83xJbfaqDTTU9NpL8PHjDHtdgOazLan7odYPBLGF9Gg1gqi5vtcS
FIq1k17md9a2VS69R+3IWQfZIx8JqjRhOUEHSpu82AG7ZmBKKniv8tNXC7RxOctHMP3UhLwAmDCb
RYhE215moSOLqiis4tmKVjlppOqHt9wO+bdcHcsDZP7JtrWbeeZLQEBnvyA3sVzPKvNy0PpQx6Ey
d59+vAosRcHbHc5yfIhpnMgMdaegSCe8ftwvj9efcOz+lNsDyyenrNSfzUF+hqMS/Kqag+XpvQIB
WkvqJAh5wWG8yAcoqDEuMzQBVf07w2VgRppVnCP+TnrlCOWi+CD5Zjf/nl4RH2n9GyyxtConOq/l
zqmZ6gyQ2UOwEeCtLktsFqwsMdbbfYwzsNdjgwRq3T13Jt3KwFXvzakmVSCTuLEyMVijiBBmfuOg
vMVmtWRERq0PWW7O3XXQqseeFoyEciwRBotwijT6bx1B5xn+91+iYsMghd6Kp7AojmW+TYYEhzXR
bbKKS7N3jW1vi7zW6oP7ToA0eZY2Y5PzzCAvbhRTAyOuiucsQa2wWtN1bJrc/dyy7329GKmjUYeY
Goys81xYl0rldOZnSBQVtp7M9xZzT8YGUfU9Xn0qcAnwPi2MDky9zMImaeYwRVqwcFDVSz820X5J
h+e/7BEakB5p/u6Q2m2w+aNcfOMWzdG5k5AgZk9ZzniQ+Bk1SR8CyruBIVk+gtaoUuyvCXF1Z7Dj
3a3YOKLmjI7LXumm/7tsmiDew7t3pp9Z/LJn2WWusMM2bzONvEdBM5leMcqhirmF9hxXIanfWOwp
40OKOkSAM6X3Psfhpt+KWwX4AAXr0UoEVE0pGXTaZTLGQi564SE+Sfil7sbc/9VzX2s7gdio5//t
7aG4dUI5wi+lqBjJd1Gi31b5FQhvGD0HICOiTNbnvnrYvWeV6PuUXRRTnqkblt0V6nMDs0y96bA+
P57upsNFegdqfbP4yyZuUQetC5WkbF6wNrApvm9eFD+9vJ6rBWuVJKMXpz3gTovzGK+I2lQgH8cy
Y6vZ39AVglw7UD5ItIhynjwrtizMm8UnDhKiGwmFDEd3O2OHEP7Umr4uLBP7EG9kePcMH8BzXTMB
Zor2TRU+VR5hiDIAAzWrsJ0EB09blm848df5G9dB5pQht/oSH0QFMJSsX8qB1ebUbppZAlFtmy3r
ov6nhTZiOSHz4ek4Bgfj9t6WmVXhCpn4vYuXzKDKi2myOQp448n+ALfuTKu43uB8VMdqwXlzF6KY
ozh97ESFrvU/CC+BiWIMzYiI3zgG9B07IpRxfnJyBiiJi+vzPGfRet8qjraeJaDLoGNlgSJJHa3o
CVpHtj1OPA8S0Ijrw6ZW/7CK/aC+VvE/RLe8af8VStMs+8xEfg1DJw2aDZGqHnBgVP3rWezhOAzz
kIWT+JmAT7yAPKFK0HHJXYwe4V4lLqWe6rZ26omXhSGEaDUXi2FXvy1acVe5A5brw/3MEQjeq6PW
934BNozDdox/+EpT/9UMNFyikVePj7tRg7JE3dENcNE9cC0OeHkzjPe01E0XRtKwuwkn4N59N1xU
XSBFkYPJwkeI0tg5aFNAOqwALjAnA8W2XNhvn+XTGZUO/S3isJznHkUtW6OoRzStuFN/6kbDHdOw
ZH9BPXHshk0UrSgGy4q7wcUt/KTbzgaKj0xcoY8VZEH1SO+lE4Rj05MMzIOjTWluZ1W4c4ydHMD4
/qkWaBYJ3ycTSPQ22RM3vMNanNckDQKhIup+BhWEIldgdS1dV0SIGpn571BiBJ5CCzh+8Ea58v3w
kM/CybDeDm1fbrWVv9+x3NwlpN7eyyQGHD5wXZpGMKcTJT15rfnpLkGqfG0sMwOV8wWTLOwYh3ok
BVZotje1BxOi1agE5tcjm/3CGKepvXl1/YKVw172wgTB2/VCLqlJC4Bul7xsCS6V04MTHz0oFhHX
O+Ci9yfR6ACntEgT3SW9RTIX7lohUQe63WklZPsfhZ16AjsEtl59/Nyd5whhmMV4cGRkktVD2lah
f+uxCMbFgcqqNMA6+iXtS9E6x52dIo7E/GWQI31i9/xUHQz8m7WiJcBXzUfv2Kf7lzBc7XWquGcA
0dPzi0xKh5Ukzvn7yXur4rOGOdzROLYUjwpol99+VvtsjPMZT02waXMcua31+t3d0ilwllX3YlqN
POz4bLU5hUge6Mnn7uak/fZBP/xRZ9ibQK7xDUiJSR56HpK7YIHryImnDW+hrU8A45EhCkQzfO0C
fnBzoICkaeMSlSUB2NSCmHCA3MnB1SMj0Gk+Th6TiMosgA5LSWXYCJ6Qiu++8eRP3kI9LJCHfOMs
3vdMTDbu0XzbRLK4RI2lY8gHwtJ4T3rkwl352LyH5R17lGVPUNHcmub7IKS4bK40IP5yr8q47kR7
35m/gdL/4OT5QBEeBxcFKo585k+D3woIVcbVwTmSgkalhLqsEWbc71YE/yh7h0QbEY+oxqmN34BI
lHL/ZjJT3r8tAyBNWlITEwZLdliKoAsngMdU3iv86dWJiG2OMmU0uZQPt2RaM9Q6sTVmLHzV6QQq
qme4zbM79dKDPdKbcvPOuG2ppBj3YJNp1UMiiICPMWxSUVJjSJOyEZNg86TbMlnGz1hc0eoeyFIA
/nHG96s1PMMIG9dYt7/pqShMGUWyfrpDVGNVR3K6stLXrbRC+xz56tntPS0J5a+XCDodZz6Z7xqj
ok5BwjFSpgvQArmWQjmVWHpVWciXZameDUSqK6AjGHer8tc8de2gF8CyBFdJ1iVc7vhWW9crBxLg
4qJpt3vBXAEhdF3KUbXIvVW/OSJL7TeX7FoW1fMmKHZrtE15a1uZc3r0yhAAeO6R/FNQlDEiUJsD
D0DWEl6H2yOJYGBLJZeRZYsoP1ouWOyoSHslU6s3PzukUu1D5OGqLg9PR+T5dHD9AzvAOZvJid5t
QhflRWO8t9o1AN50JvIXqDK+P7cJnHih5JhJ5DcZiSw30xjG9wAjq+Xwvt/jBg2oCX5RpNsczLUS
23CSSAM0bClo5V2SHx5RnjdBrdzB6HWTGIGx4D1OPHQtX14svVcDSVzaK67e1h7jGBIJf9seWHtt
FFRZDNbN8cyAOP5J9KRBAHMKwSCXev2LayFwrRbdkLKzrDyZIA8rI6ww13cZLy9THSx3DZPJBNtb
8tOVUBMohsIXmO8CCknZV2TXXfp+bMXF2e03iSgWB+zYiD7OBVMEcaRzPvvt4P4GGOyHyQFITy1a
+/HTJidzLHAKDm2G9wIhHJ5J7tYF2ONmPdO9HySFoPF8vfrSgGC0EOEDaG0+/Qnc6vmflyywDbDE
/m6Us9njqwbMrSFjL2IJvQcyrWDp4BUZk02HBoG5b7pXe6p0gxET4+sXmKh5+p/DBPiG6tQ2SklA
kz4z/a6ZAVeia2oOb9if3X7cZ2Dq29aCboeedftgXT4W9rvOf4TSS9n1ygX80AgnpZVw3jSHvkN+
BXzZdUKkk4Bj/8QrjSVWeTq+McOyV/xr38YR8YnQ0uPD9hgnCf/bTEVyMSmvPOedykaKyaR4fx77
bsjt9EII9d91jrJGznEgL9u9mHCZD3nYawR0n/GHxkuwPzsCV3eP0DRGaHm3gj97I5S86MFMGo/s
aG65IBBqo5hkJK5GGB1C56lUsHIM1BZ9yPkH+TBiiYWy11g06hTu8nKuyDWD/apT1IhxWNV4V/hL
D78hTgkjdo553sR5GyHH5PUBpV4aRb8c/E2vNYyIT8LFlwOvHFb3cZJPQChfwJRoNskNOohMFOLE
8Bqt3KY50XlledLRSDwq688G0K8cjnOJXmSW0M2W1N2H0+Kh0CCQ80FeQ15DEno7yl3CTxYg3MTr
AK69KnQb+qqT5YtpJgelJBvQhhlFc60IfN1D9fpM/hr2VKsyhnUdhAFsXxhjGeZ49dZMIpSa2ov/
fMmDskK9riMhFQ9VwuyEGKpAWdBi8jSUsvvMfaUprwVtNCfXbRQT6mWPcW7Hq5gJJ0/si7zgZ6kz
wbIKfVhr3ZyXGfCpWAX4wKuanJYqClA9MHGUpgpjl8dTd93CI+VNpaIc9GmyfTBvvBUQ7TqidEIy
MpEDgcU71OfdMsDghIcnUp/ttKZwIG/gtLjkI4eX+4kDinfKpO+qV3VEpbCDcrrShwZleHhU1GdO
8765GxmlpPSga6p3c7qr4e7lht7tIx1Wb2J6xw3BaI/KQcxEtjjniBK521IamIA+D3OAWinRy5d6
ZPOs2RjISKFFzO28Cton3HBhRntKQWtfj2UFZUXsymqdfCbLtNlsLclvmT6I2eNeObB9WW9J9X0A
B57N3hy5FbU8N+29aqxUFlCsHIVFowCqf2BpzMGJey0B+zTut0tOBcgRHh1ZFgBCVT5zJhgqGemj
0CVvbTr5sGqDFfZjQubBKcWSuRQZ2RjN+o7scfu2/T51h2GaeINX6qBHVWXobGTB7hwmXmBVYMkN
r3vi8qEbSEi63GBGa8yrHMYX9Mln17aF4s4M/0zGAXiL3xLQFF4riJGSyxydCZ7O77UUHaGdALHT
eFjB4Em0BsPv13b8FeequwtMtnWol/uiRedGMmkqx8TmqlYcdvX4jRL6zpk6L7gKT+cXjVxnZC6w
PTi3PSFWzgP7S4o3aVPdtcsKw1EWw5yReZPkXTJKhptGWWirj+RXReEKKSjLICB69km/S7ZRz8oc
qoxcyP6zriOih1IGL+TGzMHRhr25ugMAiyey5XzojzzcLbukgwIvca7rROj2fx/uL26yQbgS5LYK
pnOCg5CjbNrM8ZWDITRX0mjtId0jjZdyrsNftL34cdakUMhxO0mxgkK5LLV0CLdb01HzwDbDVMs0
Toa0WC6SK6bc+2LEG9T1r3QxXioUd+mJa0999ceTShsB+LBgzMGK3ZKkQa/k9I/Xl319dhOTO7xc
XDB0gBOgNgfmYOUZtNjPgUmbJ+7X+cf9mv3pdenFF/uSAfvZRnVuqgXg7jYECf//kEJEJF5FYrCv
++1+VxazGl9yvLu4KvD5YJpxKNh94z5PgfOJk2w0uwBrSf4L42PCSyd9p9nb6Pl9FjPX8z3qiazu
/cTD17dzbb/O/nMlyCJoDog/GuDHOBngpHXXJJ2TNd/I54YwpieUloPGiRdgaqX+X1NoNWdB9sb2
4I3fX4F2OVF1LsDEu6prMqflKHLeCBK1TwAwISa3csPYvrZAJ/9k3/o+/ebgfuL8mY2TqoEDvhD1
TD2BZy4GKDqK+ZhpIKXcMD0zh4lBksjcaFdcFF86NRie3V90+yQ8dXZnbmA/tAQsml9VtmqBx0D+
n49mtpuduknf2VGA1ng7T/z6KYLPFtsfg+EZXdDACRHdwhptKd3gpmQ9+VIBzSMPXKONmlOdNe1g
WdCY4x9j3Nek5WSdOj5oeuWNwVQIrzfkqBA3XRFxyQy5RnaBJ7qvz6mEjc9y8qrFo4O27AQEDrfb
djNDcxf0c+OYz+23z03CrsKXdf5JbS+5vTxOD5QfyYQldHf+5Pirj/aVseUvsAyTCfncawowF6/u
SP1OAe4qKEq+0UlRTn8diCqZ6UWPOzxPKy20V5EyrfpPdxHBrgUgayygdqI/slRnXcc71wPFBVES
W6QvzYP4MfcFzOZqoYavnpZJxcaqUYeyyAEVmxmZzLhuN5b/NUp9U4NQIi8x/F0y9VozmPLhrSPk
wjBxni/w9xDrbJwNwuREhOoK4RMWUb/+xW+2uvfGy3i6AwsAQCOvmwI7ykNAHdBk5r+ormLM9err
OImfYZGLZlDn6TXSGa6yCSdKzoS97h3Lgv4s3m4tn2K9OH98bSDUPbOKxvVkb7Y1O/uCyD2wtkXC
Li1poAKK59dcrTbdRlh5Q9CkXARE64/ZpL6OMgpdtVH3IZUY7sq6tXO+9RSVbQLUfRqnMwMU+hCI
NDbvHGXr8aJ3zebl+FUiIODpJdaJe2Jw/QQFP83oOUyCCtmyF9Fe6dWegsZjdcXab1YmibRFoKDB
V/pBa3o7PoNNgXtd4orp2qyxn3o3bkYsjRI5QchV0C3bBsughE0eqXyKIVTQ0UyzvlhVj3JOP7l1
U2RBQjPEfybxzfQbKEQDEs650bZU6jhmM0IUyk5VFXblbTaVWAV70OvhBEzO0uHZuRYay3VpG+yl
Andl6d3R/sncYwdAsXWG6cqNteF0apS6GhVNsdYRdAlB+tfpXP850396ngiqbs/sYsf96l0AqptX
3UAQv9PdQ/iMuuK8sunDAocC3/OX/Y8/jwtSXbM/ID3mdqfj6Wx/l8GQKSTQ9hxGtRQrbSilAkey
Py3pE1pGoPf8xtnADWp/VQnbbxOqzPtEwbM9IO+HRF9aGVXJk/ckodr1y0H/BFUH2ieweP5oAXe9
NwcBDa+Ydj48YrmQ071ubMH6Uixwih6mSD7yDvDHSfASpfq/ki6VZtoPtiK7wxbJoEF2+haUzGnj
lcmiv+6241g4TgarXCJ1L9TgrpLT4tMadjXGMn0KKC1weEapKo3tMZ85rOPOSy0sHqeG3wosJ/SK
xCEUPv2KiVOGn7qmVjXys+CJsHztgDDpEs1oHu3y0tJigY1gaPMQmKU16itrztOgBbATbnFbJGMj
vWGkofE3IOo0zoSP1gqsKEuyD2zbxCdRI/PvaSU60hWynHyIGpCwDK7mn75uXF0019G9kUcqG9XW
pxClhzRE3Z/iASGeMXE+3IP5601QEOGyEF32SfQFGtwdxAtpO6TYSK6YI+k81+7txxRy0GPz98nd
XWTD8sKufZcpQ7c5SI8awVuwCUuTvASvijyzrdM/N1VQTIZkgBopPcvoYzjo9usQmnMS4ShVqNvH
FjPBGKOtEldUXiu7wwpBii8wiO8CmYoaC0SiPR36+t8kPVUlb8wHo4vFFYI2FwlQhzS5Y1weikIO
xuoQfkAwy3/9L695wwG3CPucMv/NssbXGIqgI1efC+k1Usyx8LhQ9a+TcDqYXckTHrMtQvv0sPQ/
3cXwCVsHNfPJDlOhCmRbbxcy0MUb0KoO4oijSVaU0808XACucD1Z/NedcyOGLfXMtuWmNji+a5nw
MPDPIVCCQdn3dBGb0r06lYfu8rg5jOkXNQ5unQw7bq1UrrT/OzCL4AT4ak3xKhd1NfVIYHWNnP+t
kgRMzfJwbVRkWYWlR5VajItAFDQvQ2DQZ5Xqc0Wrv1rKS5hwzj+BvM+4DbtkiX2h4AVnff6t9TB/
d6rTi1IttJ7rJ1NvxFQ0XE61N6QDPEy+fo4hwl/TaS/7xtbHKQnjYoljROwt2qDGjGcKUp4lCIqt
BTuDLmSNTvO+pWV+MvJuVY/R43CZ7CqBNtAXPM3iMEXFuBywBMAGBL0c7HRtkX0zyanDHnFQkEn/
hwxGEFuKCaB241NiugwV54dvvcD7nZ1FPIwSlXWe4+oQ4uslunMtqb/7aFevz4R2R0tC6W7AYgqF
VYaQ6Yd1+eiQvB/GzFFI8XQNyn1G3vd62B1z3dCk19C4XJf4Upt4c6NIut0Mn2x+bacFIH+TcZFD
SOuQFCY1i4sVk9pEDH5Xz6FvKera2GormnE4sav4Qtb0+yIxASHMHKd7KbJaH6VWzsKsybCa3mUk
vQNsKQbzsPJOuZVOu91SLXqGeNOieKz8AKBf+stkl6FavtJxUaQPol0qz7sgWm1BCkczSfcHVEvA
UsmwPLMVkea3Rm4Dtc3ClhQy8VRDYGfdbO9q+B3yo702vDpowFe0gCBg/A0mNqBTmGzgC7vO7Bjd
6gtd007DuwYvfF3Kn8oT5/wZTjncPj6szs/Kinw0PIWgBZfQKC9+Qz8JLMQkZ5m6bJ6z7RNfMMVL
tw62huCdsz/256UomYpUXmhL8ZgKhN/Z3TzctIB5xFiOs0o+Pv9g3et+P7Mo276gRFXu/37edpSe
osNfp8vypbe+WOI2+Q2SFcwFan/8goiwjXGGOpms9Orwr0Z0f1+DB2tWMIJjn3N7bKJNClYqI73D
iaSIQS2aGTAaR/acRHyTYhHMXs4SbGc58Pf1ScoWnV1HKXE9DgzmaAPQu7oYEqNJ0Nfy+Kg2DPdv
iRc7RY/tj3O0Jv2rhcM2KXDyZ6tE74JTXIuhKsAXf6RhFwfcS6HcCPdFKs54VJ4JEH7Ho7hIGCNB
cbJnLKQUHuT6ysv1F3Y4PBHyugALZ0jPbdgCCLqTjzy9pnOiv0F5fSiIBwlHo7eF+g8jPoLXYuJE
kQaNmG+drKwSbSAi595y3o194+XrJEWULSK+rXBYFNICwQpvG9AovIcrj6lYh94ptTWGr5SOQNuH
aAgQzu0YZYWMG8FIpWYjSrdn52Ti5HqSchZkICfnC0RfCdaXjcJoKvUSzyfQUgilsQE0jhGNEdcE
YO7I5DMaZG885Ck8EwhuKO+qYlvEsZ/osfkiCLC+D1Q14RvgsdWWvpPY0PeVYBPqfz8fV046p7sj
Qlh3t82gG6zypu8AIuCmgThxo39CHUiGXRWk28vSf2X52HXUXKYPZALG4sLdqOxIWXLenqKkp/yd
fh1Su489PAU+Uasyz6zpDq48n5ETw+0/kGHmBRANef2C2Docz2BHWEZm3GtlfIBtnZ8BClY+8EGq
87u6N0A7DGqkHYCvoGyrQhMEpC2HgLavuHyGgOdNLl5UUS8qdsdutmFPJASGKq/ta8aNRb81TTNE
UOUTtGb+xkiWfGV5KfobgOKxk+Tohe/dIzF8iP9CdWnakS0mDysQrNb4ayvTwueC8hSnMkT8Jliw
r7hcvQi94SMHsuH/9tg42qrNsguAY4HuPo6k31gskyugtTcLGV76djbU4m97XBN3q7FW0AY9bHIu
iaX2f2XT8rEpCiC3BxG51TN11mJzMvrlNKBB4w1/OwS4eeswpB6yXR/KWtcBucx396ZpdJAHBCIx
7CSqfDGcJblLH2poAM0sKSoTRWXEJymYY7tKG3UTxoKu2Sr09xA19OmNKG5qxpRW7nOE0RTWk36L
DV0HIyg7nXN1FRFlE4WCu/1u9uEGgG35QBhTLd/YTAILaUkoXXXIhpAZGw8MCi6Lo+deVXQlesz+
NGCYL3MrHwMZOWi09/BHYgxeHzx7mnDraepPPsQZWdXqzugkGTti0bp0NLa8lVYg2mka8umK7Tdy
DJ4FkjH/kVeQdWLgPhi2UILdDn9xHQEE5aFVXB8TqN2f52jDThOvQTV+2KRjf/LniBfTtPhPHU9Z
soFQjFZfV8UTq6OC3B30FwNa279PysshA4m9gR7f/2XLKG7NYMfYM6ckZawDW2UC25urK4bnmX9Y
NbKVFu78wdn+gT+xy5as/DYKpUBCqyJZBEeJwKu4f4qNAx+qIGAu3uRcZ5Wu9JE1ES5m7OroKO35
xoAba9FnmRHEDSHR95AeYvU+WNfkwiUhJIuDf7friltcQmFgyQIIn8NyfkGVlPJWxEkCeGHiV1FA
g0BR3wO+1aRUAjdubd0TAvNiy4VbKFZiabdpW5IogaadsdQKKBiljzO6oHo/g1jnBhDge3x1v/5n
uj/9B27UYLiTTZEfccTNvFSFgFMVunvQDkVIy1jJlO2KnYqnwQvjmGiIihSrjWXFjHP14Fq3+PpK
dvYl8OzB9ZHit7jFAjWqa/qXT6k/rk3/2edgpPGLJazqPIh41QWimSQQsH+i7P559CLpalPntN/G
sNcP+BaymV3JeB5lZy5G5UjGIQE/3ZBqEztTNcrLDNKOIBp43b6EhIjXeziblyt/LAH9dG+ELBHu
+6ZdSbFEYVVF++hYP3ZjrOxwNJNbheEps+eVe9y6FPq/v9PXTQGEfL0zGxoH/vCRlmAFwADxp9/l
XTNN/85ffiLhwXfv0JuHYzwbrQGHntqbB7JR2UeEHpU78jenci31wQmhlqPgQVf61YVOJTO5D+Q3
hxeWytKxQ4SAdm6CXp6ws2cpdBte1ygIg1WQ98smkXqbcpfLVDbSZaPbpizz8gGgePlOnJoioBeL
fmn9rGRDOkbfmJRMpKY//77/IsyY738NBXUMW4jm7Z+pCEs30krGygZdAH7cHF2EcosIENS4GG+F
cKXW2NVRn9YCCqhOIpq5g2/buVKKpLdfibolLejbBz1o+cj1J9DyB6CtyNC5qoAfqLBWYByvrpaw
DMtfarMbSCbsqjo2HMIFti6pykDbGjMDP6E7/4F+/396fwWNTQOB3VhbnEM0e+z1Z96S73O9oj2R
xjO4j1oA0J/obLNhookrqIPJW7Q2ZFqGBfcE8hTfihanBANQQo5PPL+bYY0MYKxJPMRDsHXRKMwO
hp0Ih6BAIgnD2mbj0ekS2NAAAaBqY0MEsmWDDpGZaixH07CKUClMY91Y3T2qqUmbD5kScRfqtWfV
PLZyQkDXCWM0uVVomMkgb9ojluDlA3iidkyaKBSPEQd6AbqQ05jbRZO7ManbZaNQLKmhEUveEBmX
dXTpMz/vsBwXW/YphndZLc8hJy3xWRWsoDdDYEq/7RDxZ7iHz44aWYh7VMIYiEnLyaDd+1KFp8nJ
r2ag2fVo47ZjHwUJT3jMDryZtr8XbuXd41z7gSSk+F4LXxNIEkTis82XYzkzjD9BGfCROGckW66t
kzpe1BLIlHuz+qaKw6r0h/VXnqwhUSTr4ZUmGc2cscaJ22j2AQGOyL4VkcmRc0Igzy/BswUrBwHW
1A3F7WWjSBKHZTV86QiObrcEmR+EDtGq98Ny6EFvhgwcCrI+Gc9Q8CO8f6LwTii/3ur7H5Lb9SDL
5zU+QpOm+ln0sPmaLYDS5NM4Z2abfU8+BFwuT6LisF9subox6uTIHWZxUqJp8G7o2FmF2WhoXKJo
LUJNwRiFTHQuxh4sCvXU7hLam2cdobUNYeuXWJQg0+2z3owNb0nfzWs+00zaYs83ZcfTznL1ICYS
1K7G2qOtk3GOaEM/0tveobI0iNmFylrWDOyJ7xXCkgpDUNBlGAQWqTaCsInNhPCxgLBKiMcW49Yy
GkkRYIcoFuyt2FOKbWsi9Uf+sWwUW4xC3gIuiRDTnfSS/BRRfvhW6mSCcwLOZ2+n5y2qO0dDulht
LPRIDELeVqT/888bqFG6yAINSYocfqIFEpQvRPH7j1aseg8eF8zNOvx6HheoP2dRFJ023rhGxav4
OU9rPgZ/flKEd46K5v+O+VRORUlu1VVh4weO3I6zZQq2lT59czFQOD/Vo3JJNiRCL0FrW1B4tiK9
0mlyp0aBtzkLQuU2clHTTcComWBsNotnHTCqERsgIqUm2o5zeaUkK8LOmNPTTj2deKQhsvepOzta
Z8S8Rq6WW/Ik3TiguLIotor16chItxrheBMw5t5TveE31b6acNeFJ6jDeT8n/dyshcIKY3PPZyyG
xbFFF26yG6zM3eUX8SKY4PQ4cTLqQ4brFU70Kam61G9h+1E2NhdY/Pgva/BrKQ7+pjM8NWTu1qL5
+T4praQ2hl9qHOAUn3Kbzxcn7+oLdcYrF6txxPyrYFl0kUidp4Sk8BiDttjvJxv2N/JaQtKq4qir
JWP/XhcEU1gdsEAjMdZySoxci2B1IAPs8dRe7Eu4j+2xKOmwssBkjbwD5idemfO4BVA7Kq5iILRy
0UO7cYA+JBFDIl2c9/mfwaLXWKBnQTr9pofe6jdZErVksHANXBe20nspJoomJUCaejNHWoEHk0e/
jE2aFJ8uonBlDDENv5+yo+C0eRoEjicka7jWoT9oP1hjbIkK28SK2F45jndl9XR2/5vYleGJX0FU
Qsnz7RN7CnTQWnzehzT2CtKPKtfO0KBEAIVkggviJTwuuER9OH7JmxMK7wjRNzrO7bedqgwJUyRD
uVpJNyf1Lke2i0ssD4aKjW0d8oXPjnNgMyhjqTDRvwmM50uj1lDPPjaDMVR4jOg612m8WmPqlDZa
Jszcg8/tC9kHDCB1kM3tjgxnGRSZo5Gu6lxkOU85/gpbhA3tDztFEcY9vfIhdnJDHSn39Lcqo0Tp
dhzzYkd2ZJBL+kOs7i154IM2y2ZeeyiwNcEoAAb/x13j+RHL9GZn5eepAfvGOQPv2TykZC1gRmN/
6lHGX/AzybxwpBTsaKBVZqeaMG1FjKv/u5M1QLitqoWDOvH8AsEU5cQh7fCcSEnCP2BDlUcQdlHJ
uG+2eG58nz/LiiUgj2+eANayaGSloEt3O2TVsPOz9qgugNWAfsBKBxhcCsnfUoW0w2qT2+BNGt63
JX8yjhpQREG85fZmCLhHpsITkquFAAo9Y+hNE3f0oTo2qlibmaE+2kLNS2s6/WoP5Q1gSCF5RrnC
Xdn7JzepIR6WwrLXS9dXXtQf6cpsiEO67jaz1adGlmjpFhLwxbQhQCORp4fozM/4H+TRszgsoMzc
ENbqaW/hU0jNj2io4D+lyGsZPx2rbzvDLZ8YuLeoihkPXO9QDQgQwMCrg6dIG4aNcQWJn+ci1Nnf
xB2eQd3erEUVMZCS8CN3hd7JthmFaqp+ohNcxjEZ9ZnpArFXcWN61IBf4XKs+HXUYlerz3//vIxO
gkZ5LmMNk4n/9kZsVsa6JajeuNxgoZUIxJrs9J1+bIrKpUNan+tA0KXL8nD01G2OomjKXgHIPNm7
Kt2R+PjesQvELjvy9+e1msTwTSJPOzrMNWXqARvWPvw+wlWp7dgMIZJjn9JyJW1r7lFvAq9E6r+j
MoiZNvrd9dyTGTpcg9rSKp9oxwpUJgpmI0s5EqfVqzfDBoe/EJi0A3WwVDj5ZiVkOgG3G7HdYDtn
3xaQ2GLIHn0/XG10YYDMZWNSBn1E8bsXOwKWidu2waQXXClduOBWnoUZKmDzdmw+rgy4Rq4Q5mGD
i5IcOTLfAocbRvf8hAngfF0/V+oXcWhsQmOVSXmZtABYPtGgahcPcM2fYARTC0m6j+DY3Oa4W/dk
wYYcotW+SfR8ThCg92eV8yxYcqyflP+a0IBl0w97uzlAoh8HSeiIgsMbmVfx5ofwEzq276ohwloW
kDVdJzDI3jGiaH0FujWjNzg6TTj71u1JhtwqaCBUcWOVOoYLbhyxWIeVepPvL0JEciqHu9XJjvoc
aicx4cFq8QNYnbPVi1l1CXP4MIBspUfis/MvEb0PHjIY74C+CfDG/DDMcXAPHIAY32mStk56qEAw
BA9wXfjWmqDy+5IOwIMRRDPnZAXmZ1d8DkzF/9gkQgLsVeSdjEUFU6XRFinhxG+TEY2BWSauyfz3
vWXaOrjmx6rNVa3Q10thzzUrifuOWR71L4yHExayRd8hqgk6mPWv/8qktiwpNz8OjlZ4ASHA/+Uz
4VoHtDYtsZx2VXeA02vvUqcV9qc8CsNoBlOeJcjvGjbXjw1Vu2qdZWWwdPY1Yn4EvQqORuUMvkF9
e2WRy89hIChNBhbCHmSZFqHAN7l0KEYeB3Mj8CJTXRtUaIR0mLITSNIrCYkVjxIReO7oKs1HnKAA
kmOz5z5ka6RNfce7hC9d5/GiDqsqzfh7/fG3NUTZRSptTGhQleRjOtitz9gN+IDH4OLu31KiFiyc
jOrHI/qlHkY+i2yKytDQJruI9sYp+Bz1OlL3LuDaRuPsqdYGcTVVnDqb7CK6NUHxdyhDscfVxk73
4z5+MJ6gnoKzfmnefuirLGdqFO/GjBNeVXImgDaEuz2uVwgylpRDI5K+Z9M8Z1W1fzmcJqGhYKNn
jiDVllVeEFbl8YczAlf3dQc+4raU5s1wPWwPf99R0+3TNatsTQEYYh0axH+16nU2Z3n3C2nrAhvP
yZS2qv1n1o0CHNkYvHPHPxdxItHCScjrAWWY+/h5wiz8nvF56Kwvgs6JmNuzKuOBDNkX+eaEnMW/
+e8T2/Id6gykxQYKt7th+RdzCLHhynwGY5ThI7KVHY7SCI0823yn4jaj2gFGq5fKIAW+p/i2/wqM
d9eGHI3dvm75z8edJq+MdzLcDnHGHi3GSLyckinvcdiphdUfi4mKKAISbcQ9zLgM20aPhag+cvKW
SixatTBx3ElqeerfOuuna8ThkrLaUq1TvGo7ym00hgivteJycdQXEsJUS8d+lBJH63JRaYiLcMSE
42vEZOKj6XDcXfZc6+d4ClxzrD0Xk6xPs3WV3hFNqjfg8VuZMjKFuKQTe4RkMIiGrdyi2bETUdlX
zhT533NkR9pC/H/AT+cEXBCxmgS+FYlMLZCvTWQMh8Rz+aZzJcpeGORIlqoz3OVlribyconWYNZv
6ZGtyUbXiK/8H3SEDpJHoD6I0xtFZnSBQx6UVxbYK/9iA3rKIcHJio2Pu0fOnPGOLiEZNU7O4Glz
UgWmiLX+gu1HMAAqDqhURpdp8009opTPxtwK3X+hFcdZkxs9h85bHo1bj0UKz3jNH4JzhEs6IBhz
uJe0RrqfO4Zumc5cgAkW5mjRDIXIk0FdeB/klXv8KEiWurjjgLo2MyrX/Obm7pcURrW1yFXRfRfi
Ik8724MgPtLlngO/HZm1fgMPpshefnjwEjF2g3A8bpqoQdPXRtkiW7BJR/eqvuevlsvF/tzk/t71
espaXZGXAcHyOxxXM/ryeqEABNHU7sBwBhEP1HGeKy3Fobq3I1pggLMSH6E8aGRF0scPY/f8IEUO
0wjEZgFyKPjOD0RrWy9QMM+WSEBE3yDh4peBugN2BroWezLV5Xb9MufpDOxrvjxUlh8lw+QAeNpQ
gj6qB2NeGpZfTUDHm8Uj6/NRZHeSxLqkdcRp/xHdzYlHygDFRHCbyDoHbgjMcU9OBMlm334Nu+3d
64VKuDMWag5WJ1ibDDIeoXtT9516ER7wJ6fo8IPdIephXAXhOVpkUi+Vm8SsKMy19i/sfFHUcnbO
RT45VUT11Xizy3ToSEienJ3XxM8om/mgdYlvxE9ztUMpunLgOrwOIZfgyhZVGTQYkIg57oTDLEQE
90R5noHjB2LU7MsLYNRXzLg8DiFkCusiI56Ha66ZY11Yk8PHfLb4tkAImh6CCc5wq2BQNmizwj6Y
kNmx3kWeTcqq56H1qixZKkpzUAopxb9ju4bBdbXCu0AT6D1bn9F3s0MwWeBT6oDM9FrnWirNmYuo
rsYuIlx5mb3Yw95peGjxfxvoG8+XS3LHRcFthCaL7j6WbPEnBlig6Oz5+1ihU4eA9TrATNnKBIWL
3AaKtGwnElZ936VPrfef8sfrs7OhdSuPesd7J4WGttwxhJ/GEVYQKNYXpueyos/r8eqRbyTWDRP+
wt96gyEB46CERlmAFlMlv90zYUXkVl/xGydTc8Ybes7SVWma+zZzBo/l03C1vPDz4rTy79OvGhKk
NOXaW4qPDJBQ6vnrdgDoT6UM/zii/dLzDsyvHTxx4vct7+sNllNdIXTT+1pb6uICN4O0dkPFltS+
vS4InYKVptgFsjb8Tr7fHgFjUtj9X4oD9YpXjDVUVh6Mt8lHyiqvnnxPQTv7xLDx43wMgxpi2NTU
u1olcybpM1bXUITPTaa6udgqHRM9IWt3tBomedDhydKBtEvoLqoeBvmN8eP+et4xuZ2kSbpd3VRh
PcjxOiR7Yrt4CFQyK2zogRyFXJcswKWaSc2DOH1tncY5kVAwCwJBWBNiJy5P8gchqJ/vBQp3f4eF
HsGUMU1CIPwm1WOwUAEme+RrJ7c38yVAVAIlmSFnI7+fqgoUlRVUF43rvBMX4n0ARRbYiwoKvPKg
jZsTdumWBHgRKiPF76KCA08mUshFMAVWBodjUQ4px2M9jYvNilgUqboHULybaX0T7GHFQZxmvPt4
vifIv0i7SJFrvaBUgwxBpReKL98ZBlj+51DrcKpoEubOCydjhbNVw/yAM/VGWkpNIOj8OGBhh8mO
EH29meHPY7frZMMXNu8x9+P/sZ+hA9pkuSc3D45HW5Rw/+Hm7iTYvTtu2evVbYY6eMfeUGJjqs2c
DDk+VkWyc9202ny0wxcIDOE1ppDpTp9QzA6v9JQPsLWQST+paMc7V8PqVvj8gqXtqxUAGubbhJ1o
Yjn0SKnv6deJBFD1MAE99yyeiK//Sik4MV357ph8nLfccTLdnHZQ4vb+e8qGAphIpJ5yQuV7ItWU
7TF7hGQmW5rlwxHJclWkcl5ReCqBsa6ZshIstR3l8Lx2ZwyB9RwScGNZs3nWG7l/pOOCstED42Lc
C9EElti9GEtNdtpRvY91kOO818kUlLmnm72lD++3Q9atIbGaVq56y1Yp49ZU6dZii+Qg4DckhGs1
oTR6NCSt/nLvQSKQ/mrLB6l8arDn+MJ7Uqy0bXHx1omNhKDIlJkSWAlWdZ5Kz5ncQve4r2nSHmo9
0lnU8mMd6EkMqY+bVs3NSzu2awyuYBIMrVDpASXmdI2AS3eQGSqlkRVr1rSElVMf2iQsDc7mZt3G
EqV4cs5mgfEzSrTKf0lIO6tiAmvx/W/otyOE8oWJU+7uGrtzTDgnkN2Qsj7M9rqx7VwZzRaeXNBl
DIEVQG5u3wh4n/NOUV9YAaisrSsBpo5bL4ROQpkRaToFX6+hUmecH9TrGrIsU6s3ehMJVtgiIndJ
tR5dymgUMFyAM7mN5hT80BqRRDHQq9YaNTeyHBRZSlp4RnFSkWAxMB750dKHjWaX1PGnVubQbHTh
WPB4+FBUhy+CZPXZY+ryYCct7MGlhjAlHbTueHHi6rLzRU8TvFeqDJrXIq/MbDZWqeOUG044+rqX
nclbjKk+u8ByJYMcDGti6KYf04i45GDFKC/x1W1xznKfXBgmjqzvtGXSWimS9j8iU6hpc3CRgjMK
q9rGSkm3t6oRXcAhRqyUWiJwaqohmFxN2rR0iutuqaZiyUhfWJ8tvwXZwBqGKWWxrru7VU5cq/rJ
3y9OIaBz/27/FGie3kDksc8hpk7cKSWOAg0pWN8guHTSw9zCGHWKXjMc4kqetF6kzElZoJQrn/cQ
cqXZ1no/l3lqdvU0Zc93UyFXerxUM/rNtMc/7N6cGxVtf1nyxbvUaBZdn8ZzFRs4z1Q1+nvYgGN7
QvbDfteYcxI+QV1c0Hzdj+0tLC6/xqWU7N7hifRNqgK44Vl1cp+p8yuf0zIMEsBqVU7QNU/IBUt2
sR9+lOa3syCzoBNVwphRgZimyxqpGA4sDfTlloat76+iusJ7e+hNRwHXrlnem7z3eoLO5dNkVcH8
gRm5thqYoA6LepSNluAK0EBCnNRzaqgx+Fr88M/1pCAHueL/9s35L9E6lK4iBRBD7uUpeLeIisn8
a+4BTNIMqMUbZU1bIA0jpzI3vaw8y7Oi6VKRJ91JEkR+t019J0Uh2GVACBQBJaq2LMfc53k9rCE/
u8eS8JNqYryrykEXzWNbqjvsHhpgTGwusCcyfZxymiFs1yiWKyXrvycjg4d5wjUIkv1gpL7dDVQr
DVrsWZvE7O6daCdjhrUuMi2A66ZlplK+7IK8m+5mQOU812fCJlnghxKpIUXvzEGAJ5qdrQftvYXW
UQzovlMTupJbQJx4qngjodFwcV3VdGKZTGw2qyXlnQXWYbakBPg7YJKVVGijnX3f/azsmoT/826H
ybp7EnB9Yp0UxQWptvW+I8T1WhGXO4zGS008KH1/ZTdcU9L4aTmB5Am/WmoR77nts0fCxgpXSc59
vTYqrRwVJnscfLPPR5Gu9hCyqvDUtrbQvcEbZFhvmRtBbJHGH9LYrSDwDXH6QfPtVnRTvQ5NHmvv
fEACrY7PBzC05278XLCpWFXt2QXZjP2PLeBBU/znqwMPYYPHSYiqSl7lTfBDm9DRDoUgnGmtkw6m
YWC1GRctTTXH9lQixIE+eGhnExWdyNfd17D6+onuV/PQM1k3RM1M6YNQza/PHFGPayIhwIK8XnrB
oBDC2t9g61NCxqkMULhdtN1qOV4ufDhqzUgxxUQbCGqfN4Tmw009EopfmG5x5YGkDbntAfvK5FSi
n0C5545MR4uTL5fkwnKwTC0GgM0q3RipitHWrf9Ze4br6p89kMEXiNpF7Tfm2/C14PZ41fSFUhDK
dEoBdJSxSZAhSRfJDJ6qzavPkJ/JagYchOlxz5JDpE/UO+KJJnlhA8yZxA3UkDzfpyxGjob/bJ4n
LT7MSCW8+uQK0+aWmdiwA07tYSXPIO9pp1AEZ4AUQsPJYICAdokWIZ1GPp31Y/O/Ug1phKt4ppd8
2iYWjzqxdJam3E5gG/wxVpWxSfXOuWxN+oczkVDOm7h6ZwMRCYpMDBwrRc5RTGHsj0JoM8ciuP9K
G/f+ly4aHlNiPFie9XxXYkIWByWaPnLwskpTMa0wjiCHl5IjNvdT0Yvmfi9+SzspyL4XkqJIQKcY
Fcl92zMJNVgUhwjVIc6ofXRKarrFcOgQ9VjPlFw60En5rKea2AHOD1M+iCEGA0L8eIFjXKmFqWpT
xgTpjgstqeq36aLlhDg2izhUmhadQB7yufGe6MFOBbiIovboVAiwf+csBQ19bFGIyPGKL6TKSoO9
1zSDW7H8VNhWE/IpyOH0lOm9CAsLnA9qxwaPfT5mw7CSnPRtgqKmsVm7Ef28qIG/b1GF66xS0P5+
SsUVeMYKRLHCXdl79j5nRHJkREllSpQy56XIQwm9neD8ElwXMwyQykJpGM4bJ4aVYBa8zlh8fz81
6ZUzmn5nrngCd8bTKrXSMgcJekEmhHtB1Mzi3QZfIg3DwhLh8sPuNCgQnLmKA+1bxtMxxXYmjpu8
CJI2n/42GkR+jw8pR3YXB+2N1g/lkxDoaxHP0Ss3Y/PmBU+yDVLa7QNmpAYyJn15UnrFwUdeqgJ2
95wclWyLGnZUugzNabI9g20bqFzITf7jEWwpWqHsLZc7zfAJNTrWV8EQVArw5h60N3RKQmeDXKnT
N7Kiq1GzroTZ83bWlb3vw51i45dCJrTmAgRWbgdZqUKhZPmfqP1dDpAbb4g4UbnhGWQA4nVh4XkO
yeNHfPMY4J9W4gTPUKF59RWf2rVe9e1CoW6AQ7oOmceJg0kVHjTFBp6fl2xpswZ4HNiGy4XuIoor
3gu35BMwJd+UVML+ibUEMQpm2o6IUVl0M0gXO16nmTLje29hxMqkUuJb+QrBmtey+8cQSVLPTGyZ
zKZZdtXW7jYOCyFEGoGD7Uao0BEd6e8XIknwo08AVUHO7/kIiqTPiLGJxHX+v7MBOjRKBrZ7v5bv
mgOeBxbq05cLTFSwBGDLSoJRnCGCCqzTvx62Bk0ArdEqWeU9hOZaTu/WQikW55z9aHBeCUD/066q
Z0K4gOOVpcbAVqNz+wPpHOeOggUK8M4czRn5xLm6rgbs9Z9lWScQ8ICNcGpxUKJJhKmZpcYMPbi9
CbaLw3L06wJBkSEhx2NtFy7Rr9szm+m7pUaFFzkXzG7kpnnAdbuosDi/CH8R2kmbVUMVNys84AhY
sYuSOgHvsxPNtRpqEcaXiB/+clcX9yZ82YeeCL0LBaAotdHiam5K2uAS1hW/9HAFhz5nf+zJvc+w
CgLGnYQ+5Eq8lhu8/HawS1pKgCoMk9L7ARJ9hUpg3WQOpmxFrQPEts/kgZ5mLuM8tdRlI2lXeQsN
xjTw9RNVC96Ul79bm379mjPtOnYLJ/Cnb6amJ+q+R+MlxwtDihsLzAQHoKbG4fGrbZkUG2hOtG5e
/20JXNJNLgMlS/lght6toh5TajBcTS2vnhuepSShGCnW/mfDTz2zYrRD8X6w3sdX7JeAD9EHIC2x
W3wcpjKMVzbqmDsOshnDMBFW5vCXQLHQzLn5Y5G7cL4/8r0wtn2ZM1C0P2rr9JrJYcMrKE0wcC/5
gDa3qEXmXfP8OOaPiuuXOGc8jAJVrAt6n+1hMMTtfjCfX+aEaZU+W8LDS1CSramUd01yh8uvhXiB
vwiT5t+TxvpOb9I+eXfFRykLDv1UiiI2NRmRFYLLLNG3aFm+idscGxOeyzEXh7hjLRtCeH3lmp2p
a8n56tSmh7qwiH1UMG3UrPohZA0cYEOKGP/H59bI3RFbOHVR08Mv34xjqX4eu1qHFuqiAS2Y8IP0
A4u+xH7dcfNvX6LVfx8RZ7FM2TFfEf60uTSqHjMrerUqLTjKSVroaXEryvpS3vVkWT2kr4J5eKpy
3uBx0y+OSgOVh/bt3aDuBbSqW2YXDzQVITH2jzRuUS14fyUPPSJwllGm3l9blX64+koKkGsNiL5W
4XOqt0EDkM+mDJ5OGPYTHk2NYQAvGFcH3p2MysoEUD9AeOXrlM3ptvUIBMZW9HL+AWWCtlKm8cH3
DAdqoyBGTEkqWlQAmc8vxZ7Vh7MC8kWiTpL1YzWhbP7vRP6JnuI0AALN477d+pVbeB8GTJwNRPrj
Mpi0NvC8YM2aiZvCNftXhrXjLNql+TmzeFFGG/nmrkHJ+eEX1MCKwttXLlHCYcpGkavf2b5THtP7
KnCDvOfOwK34Mc66UvXq+fa6XFJRAN43zcUS+bqRVsnEXS6Kk6hXcUPFrLk/G6Cq8qWW6SGUR3Zt
EciKlUdCf6fh0u+mZdYNZDA3lxdvCBatKEVf2tenj0f8bJALs6utrgRjW3ie2Jmgbf4ENoNgPSKw
VAne3MnMvqRO2jH++1m59pMvyURSizFYzfZnAda9zP2lv68axHT4omUS79UyI8JTBjQEYfqVhbAn
Dl+mJj+MCyaRBtqHR8LEIRWJj6LlY7BbkjgTUyFURNYirjPuHgeID431I4oqOuOjKqbqkkl++5q6
Ljiiqwh93287SyCUQSjRtNj+T2VVb46O6mnPmg+31oDem5FxgOK46WQr7cg/IARAu3BBlwul/LGk
IP08S5YpoFQwJkc4o3Kre4U1ElG0uWDNZeyi1sBLYUUm2UvFjnE8ROuVDjzOevIMtWc5ykiwzkez
I4ne0dKlmzatBkUER7hW1y8/jRRfcuS9Oc8WBEXd8Ca3YJvzxS6/qPYjnEsu3h9q6WRajRKvjCwq
KusRoSciH21deWlxorNyvn/JpdbNSNBJ/C3RrsBc5oI61wwxVfwMbkfBYAG0qtHtfxdKIqII9Z4a
LcxyuEGT7TBcayBXfGyruggHwx0HF0nP/Swuez4Nna89QjJm7FA5wp+F6RagB08BIgRBnib8GqTL
JP4EcBeHx9zL3HWi4TvqTN3qn3d8SoGaQOdwkDZilWRFdcofA5Iuze8ohNr0BLdrjRB6PqHNzmgb
StHHPpIMxVw+Yf6gEC7pTDoBOp6nej8dttNpkP+UHFjQ9kDRBwFEgE5XeecOP6u7fNtnX0MoUqXI
79rhtyzoJ9wv4ClNXDKJCsDZQ4TzanXpze+xKbfaAA/L6gHj7hPo/impl6pcLQJKfjVWY/jbsDZp
PiDHrH7EEgx7LN5NC8PRrQZDXvR9PtOBe7wf4DTxjx9lvYpI3XXqBMtkOCme4BuUxOez1KzR0H9M
pX72bdbBoXjIPRxjlvyJj9BjM4tEARxPbZ1Tw9pEIKHqjX1qMllrh7R92Xpgtg0V2bW6YWcvFgxf
INORzVGlCKfV9FowxPqTTzsuo2T+WFZjEsHhMfXx0MfVcLFvy5PIu7hnI0SHcRYqlI/yvD2wAQ8Q
6XOQcSH5lMrsAxtJubosz8EB2SN+ZZB1CDn4wnOKi1ek4Sza9xSEeAaOHZctpdW7TyTuULa8woTU
CrFnNIFQ+1uJvW0nzH5e9Ke5RNjSjgT+boTy/hpOZ6xLdZFj05ggfeVJjVAdJZmV7cMANEqYyek2
xJNNLic1u+eNkkUpRtiOgcBZOzS8JACXdQzpdDUZFtT1gCf71ZPN6Mm+BT1+v571J53YKAbTNC/C
kfAqYFis5Kv0njNQToNUg6mBH+gM03RuZMG3Sk7tp4NMDw190CRUwTw6dg/oRN6BLo/RJFrhgOoF
zZuhvMBAVRS9jaHVGwU6SuBcMtPWFMXrBUiwZP6hUdOFEU0ByME8CZV6rY1QB1bkmaDhLzyHXZx5
Rigg2wQ9mCdaAY+zlQwfmmEWJ61P2usad9FDeiHCVuKjCxu4DYrh4lo+xqai+vtRVtSUZU4iIvWL
psRBfeyAuOe/2jKyh9uhOyRAUh+65AUDsB30E2XY0F8v/osV2JHo7jG3bkryHKFJF2kAdmrVa+bd
aiJOjppyKhKNDHKd0unwXxQxBsi0CimTZk14UppPpivaulbJXfVi0iwtCaiqskwI0eezhAW6Mc0F
SXytAveC7KmLP6grz64lm9b3s99M31QEgmCVUdEAzLUTpfwt/SA72kFdubBb5yzb8ZQ7yjvXrZ3k
JkWl7hYY9bW+a+xzQSkJ1sAsIpu0y5Qe0JWNeuFrDadM5DbzI0r4B5cYFdZQfD7enCgEci0BN08g
yaAQ4dFyBDae2PPghBx+TEKKmIhkdDgr6wzEr4pxzojuYAMr9W/9HgHaPYfJ1d6HyYp9X3yVABp7
GbfOudaQYpG/WGoBg8o43pl1Rt/dPPAveg7wLJNHi2q7wSMvylr7xjMQPECIMi9qLlfHjicuMgSC
TOpl6X8pmZlHeJmnZMqpC72aM4Q7DG8fTlF6voXm1RU5Ye4z2+I+Dnwyn7sTijd6woTAl7RCLOcx
WNiRkL0whrCVmwjrEZ1D8DQGtK3afTm1gOT6eU3LnA0a+6Bjm+3mgjCnuL6TUjwY1747DKJwNH/d
h2Az6gASM8f4V2SOvi9dp3jvNUAJHEGGP3h0d9OP2aNCdZ6P/ndf+d3hs3dWQ//0oDvYoUIkKxE/
s8UXS6ZrTYCPYGXQNaviWpN1uvf+CE3uUfj6GUKckB91Q7vV5RCw7bbBJc180c8wMfECVEOcmViQ
7Z5UpvE9Fc9HEFUwDi00knh4jEFoYRCXT3iW8sg6U2Msefz10F8yI8lYEjOCyknRZfO6zpvywc2Q
kVVT/w1eFDtSuryGsgW+3dYR/E4JFNFVVPqjsRj6zataakNmKqjgeQTr8MdkVAaiS1t4VTdJrLIJ
hL8kgHHrOYWuXUEA99gBVp/jsjcEZRsNRVjvaz/LnliVQGexTICaL4TBDiVYMJ6eNhcMixlwRQ5+
VjUy8e+5iuhHzRRTnyBHAo5ORgWWnwiH4o/e39lx+KB7hpJ/+svHZEJwf9sSVIG+qesynn7EcSHY
P1jBAWyUX9pf2oOK98FpxyOcKz1Cboussz8SxZPYLbB3JSa8nchYdFZlvyyS9ZnmfAiIt2pyY4B2
S8BeBfTHQixmO6LZJnoITOTvj8pS043AdUM54kJAsa+vPz1vMi7132zeX3C7rC4vgz5NywhXo25f
+dI2G7a03yR+aQ7LbvLqDMxn5rhKcWYSd89KhAputG98gL1Gg3hap6DE7KL7GdZIrW7oZAl3Tt/T
Hs6keOP8Sl6DVCulXfpeZq/RRnQkosd6kE8vDDZtgMOLLkgMiEWTghf1QtbD2rhUe+uKvcK5Xn2E
mjMDAo1gvr1SGHmROOJiwhZr2llSYAKadjvodW99Rzzq1IIYdYoBEuiv88DNPy+rzZixPENmBwZ8
56tkPLxmXJMDlmqB1bgpLb0N9s/fm575zttltKJ1oyq5t8scbe2yeLyiwmZMpI++HhuCiQ9Wtn1u
8MKnOXCmsRjo4upb/fLZgEI/ErR98GRsxZrCT1vGRxDD9dJl7G1C/zC/sGSQGNSbzI+J2yEmyMuG
JOU01/zVYX1HmQwqUM3C6e5m/pyLOtUFeUcXt0q5TFP18fdqXR+RmkN5jGTfooVB9/EA8OAAdwp+
iM5ljgRGPLNVxW+ZTd0Aw8cgUDTgK6kYwcIyDTIQGi5YXScHWSgKR7qhD6JVO+KSkt1rTRKWGhsG
JivC2TzXghWwvv+VRposoowagNKtKpkpE6F84ZfajeHrnA5cC17+6dkDann6Q8wuZl/JIRnzFiwn
92Mwuep+c1enUjNR77pu4XB5CRQDhVzATRJ7y5YBO7Hf8Fo3UMrfArMmBH3yz0NquSRIhGvJsZ3K
itWnTUWc7n4XPlUmXueijdcJFl8nyHItO0JDy/PEgoDFvnCCf5kEobKcOZTgEXT6ugZDQT3gcM8o
cxrw3aojDnS3Gi/gV79aZR1mipCPqXgrtnPn9hRkkCTaU3sbYFhoeVNhq0MoUbW3L3gRPnXQL37V
sTD51SqySsV02vLe/P2wGBP3Jy70nkNx+HTZ07ZQO+0EVKW/Elcfsq1/6ktcYtginGdG3eFDqipE
P2ghMnIQBLpai64l6kisoIpjqqFfrWX91JUDJSN/tH0gFRpWCqNuByUDsqLkyMaFbTiYidgTK5Cz
frvpywqc65u7/jtaswQQkI0ci1DWj2/gd8PRv8WkhvWwDTFPtpNXpdqbVZTUzLwFc0zz8Upx38lu
imG6AvHP6FAnWwTBNqigpaonfsykEW13DDMi9YZvsplOacnfHUDKGO3uf0rUqP5fOds8hE6eCrSN
kEsI2+Ahq0NtJiEJHvJSdAR45ksE1auIsmY1fEVVb5rAI8bKB15ABmYkUegKxrJIDyoFyv9Je4G1
+cMg0fMYGvlA/5PFcivZzM6Mp1xRipHwgQMOJFqJtCAMuWlYxX/EGwf6cL/eBUvsVOuQpoYNrvOt
xNTOM3aD8jTBD2rbknpxHmTOnAAGEDEE6z7GEPdYmzlYCl7d+KXZ0Lcw23fJS5GCxDoxNG8FZFO6
Gepd0lheBoQOlw==
`protect end_protected

