

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N0hMcXbI5hCFMXvbzZaWNMXky7Cb78UlPrOh26mC4IyomLPXkDt4pohvBi74RwhMjj/Bp6A1/EjU
BW4AL9d6yw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O4cgU289ETKimPPpC1lQoWfngvpNmR5tUZAEw+00K8UK2gEeqXn1hb3g7AZENGEwMii7hns4XQy8
DXQ5xw0Yp1Lt5kPvabj5mKM1bMdX8dvR9NHP3g1Qjd7okAVBl07/JG0NTnpHDOfWPgdIKiG5gomz
/inOtmJ9dyw3SQwornQ=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DU+IJVy0UCp9Ru4O1AHH4hAsURQvG4KWjfdJuBdXBn/Aw7vf76lLrDggWEsh/tDsD2w8gcTI1KZj
gte8Qz0RBjJA/tV/Q7C3IGP9sKs04WbpHeToWiLkJhGVSOi1cfBwcXqun7kk3rw8tbtRvnn4LLnQ
VVSnOUM0P3u3t9b+354=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VU2OWBPAFdMWY9YsdLW9vHBQultKfSyqJgSm8GFxf210g4AV7503RY1sTzcwbpKduWx2mEapVrlR
2+Drhdzv1Rts/cH1vI36ZrlUVzIXAPfly2Vw/ZI3vZ8ecksIx4K68q0S13FJLdHLryPXLuFGokYw
gCOZnAxTuOQQMCgsJA0iDJVXFdmLXzqwRYBXguqf1r+OMVPXs57gcwlgVB8r2wrtRxBvH0uRcmEd
9XDbIcnUXETCLhyRgVVpblWBh8bZbcQBY/zZZ/sbyAPD6J7Rp8CEPhLVVCsK4EjNey5PsDgo/izg
h4bUKLC5eF2W7tVckgp7jyOfw3DgIr/wn7RxeQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V2G0fgDEE2OFe05Cx8OR1KsgdINzVEXBIBadpSnPXIoTc7xRwAe4/VP6V+6MXz0QrLZuQHVAj7G3
9F/ijf7v4vM07B7zCCzqKWXPOd8bPZE51/A2H7Mt+ilGqjbh/VKLmxGs4hilsENWISKVXeBdKnPY
gj2HGvaphMJpBpJwjPAKBmbUyTX5Sd9nNIMzcSRJNulwiaiEOrABFlrZOI+c7bZY5sHmVeOtg9CQ
vhwpJiZDt2xEUYZdJ+nAzC0+NS9jg6KFWoyyUeNOwHZC9//fhh1MCUzJ0nZg2R4hBpRaxLZstp3w
PM0at5MBtCkDuhRItVUmq9A0HtCUCEmB412P1w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RN/6I+vbSUSbgQKZutSOM516q9s9JryaK6V/qqxo3gcYd+gU9W/srRAx8TWXTu0WbgzNnJ4y7Myb
hqdFZXcfJ/PxMgXPrrBTM9dc9q6Om0xxWrgSNxYalV3KY2vgAYOZai6mnccqhDfT+ZicibnnsYmh
yf5l9IBMwTbxQ9cpGytJTrr0jtjFG8izeH9CEj3vxYZQ4tA0TFJhsFvQhk2xXEnWnEBhTQbSX/B3
CADhGzXitOUqpBt3ylEkYkNM5wRAzze9LtBQhOCFWc4AJq4+3/P22qqco2g+VSDFNt7Sbc/BGwyj
q/3tdC0FZkEZB5DXnSDvgc9OVq2Fggic0aDyNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
ZD842BQwol5M6XdsOj/OdDZsYkB0ipsAKlCXkrbCaPGw+/PyZr3Y/OISZjZAxhM2kclxsQ6UBVT4
oNNO8jnithmViXSd92a4Z0TyqLVWD9zbXVErGIn6y7ZJcZnWbSmbNcTuXY+FVa1CVEHEkOULbBk9
ro0P8j8vrztMC4kdEGznoY/iP3Pf971W0nWBw98P6473vqY3BsnM6NZNFofKyfFF5M+Cr7TKTDwV
mB9cmgob0mqfKfk/S6po48nGguQqY3NoTTskhEMVbj89mDefe6tLZGqovp2jW/uqKXMJ4g2BkPTU
6V1ThQLV0OxzDZcQo1sqKeby0bDZr0c/7DPAkropG6DIO3MrKkK10YpNb49MRv+f9MJaUpON0Bcb
bcDE6TbCnFycfO7xe2wSY0oYt0H6MFmvtJDTPRKv7QXDCVwGbeeFyjkc8IW6W7xl9AHH+OgMM+QS
bkr3qY+ZB7O4LuDX4xwHZrErBJjtVeIcrvnfJ2PLdX9MzpHLWUypzoke03vc/5yjw0TgommWDsqY
3OVVy8TwUPH3mzp3fletVKxNasYabDPRmwD/NPF93795SAyO5AQt6Z4zQthH8CWVpxV4DkjXD7hO
G8rmiAM/p5McSZYDMOsdzz/Iid53R7Yf/tQpA/TMnVQWKNRLlIa7jqGThyLW9YYlYaQaifdy2wdx
CUjpnPBThulRRnAOGoFJpqMDlCdEB/ruV4GRPX//5pWV5A4D7zpbDOnMUWdzov5uroGFNr21/dg/
mQRWXwkBO0UVBNUt66hPf8KndGE0HN4HdbooN1oGH7Ljd3cjGVWjWTiEw7bB5oK5SfGfzq4LAumh
oH7kKAxvYLqpQbeF4METthN/lb3LjimYg3lu88MmeXO46DWsYj12ZJV7hAIp7LczU6ptJ3i7vGb5
x/96MPEzQCKpGu/JJ6MpphE7FuaOgsJrfqIPkZkAWQ9yCH/80IoDOsdftLNpPQv0Ft82WKTzpi4H
hWJIgLQGeyrpJVtLvoDx7VNEIiGC3PQSgNZpyvLpOAmUpyXZ/zK5neuJ10+uN57Dv8+8RP5sbn/n
j2vUOB1RF/otpESN+iAwbVWPGZt7lLBnXE4TA4lgIJAdgtYGIebDR8Wk63WA0bGRAy3itJAMv1Rg
Ger6aoNtJRvH0F11MaMOzKCuqRBrC5XeanEkKyaVfuAYz/xfyftBs+5QGWmL3VvLpZyQmc2BoM3S
QX3AiHj+TzDrhEXSntYArfzKQgE6n1OC6VD6Etp9mcIs5KH1aP1G1AIM6/NX9axs7qZ2/s7QeDqK
1V/cRJ2GhCQQz+lFIKp257O5ml2seLjndRqVy14elK4gyvNo17yDhBjzCrRddSU1fh+Eji8tLpYc
XtTcos616LbeMCwFOxshvnPnA0i3pHuDKmQpDide8LPAJFEC4vtdoHtI0ez5saxD47l55CN6r+YW
FpD3XaL5oqfYmiBHkq5vw+KTZ6GpcmNEX9n0ctK/tk1/6l4BliQFPXhozGoB+ywKuEX7C9PIsQBE
1FIKKvW2bwsk28poXhaSFF2oAEfD7mj+d2VzmGcZK9qQpKynBk6MMTFkRcbqSj49EfUnaJqMcaZc
4sB4k0BKnL5Ya75cR+wPeuLtf8HxjamWFxJQQDTfnnTU9RQzuLpx7NiBLNUzC7ByznpgOZLl9a7e
8mviCO10jEDq7WU/PtvO3UfA0xsYibRpM1YJXgQJVsAPDis05panPw/YqK73s8AsYLb6z1QE68Pe
8RMnfYyiUD+g3El9B1e9o4YSOPsOC2rOZaKQjhvGmneca5QW5mVwutg3fmlMnYTZng2XOr1ue61m
djifjb4uyF5AFkbmOCPxopAvVge6TlxkuO9JPNXO7IuIIZaIkEpQgyYmImeRtvsU1dgx/TmuDmA/
/KMUR9KSNjTVZPUJLQWbXFq1qR1Cw4A2gfH6cIpcNC38SKyu7QKrT9rSQtIh1rtAdAvZaLbLPM8V
/WmcRJF8+kcDpZG21lsVC/0C0Dz2A9NjtHnNcIZzmXpie3szWZDM7HZMUAGNuUFahztl0nk+VKyr
ptEpBZpZve9gpFqjaewlCnLohBNt9j5h41ngDuf7bRU73ChXBWeQfWzVt+2D8GCH+ThPwNOY3/6Y
68RlKqiL3FtZBiuz1wDcIe65BDgS4wkolZrCN27YQxeQmR4stX64FS4X1j6G4NLYJ4X2wanU33ls
RiRoiPvQz5MpoPWbVfO/fkdEexgJQc+xKpaLT7VQkdgdSBJVH/k36t51RBYSyS/YPEv3EAvSKte4
qME1Sm3feTzEI30LlbXdhfoUSPsXZNFxQYUvde6A9+M+g7UOe+Ec4o/t9o7ufd70kIeHTCZanUrZ
ns8lJQfPdpVXk1mZUjDP+BJ5r66y4IY9QwsTVucKX9ATEsco8KQbAOrx0AWGLtOJgyGzyCG6aEJ/
1RtlXJTAmCAE4vx/CPdWVIAVqdvy1KqEPZ2TcKfhgPg0z/NAIAlIZzEFmCpZ/f4AKMyTLFnJiZ2T
kAM2mrkv1qCa0ejZ+HX0D1PT8LIpMwLkRSsAfI9yVn7ir29r20MYbng4uM8M3agjKvxpvtqvR/lq
EMK4rqUzaxfXlM1yBEvyAEov9Hg6MFXTIE2qexWLvs56aF2R/moMaHLahsxfEt5GvGtd/SeW8CQo
8SMh1WD7MZQS5bzMmtBIj4uRSlj66cKwsAk2BI3rHZGOP3MJHzMR2fRfAwtSwYo7LuTomPeWhjQp
VgTM8J4MGJKUNaqHq6d8CYRzjuxlDUooRocmsKefMgSZEbud1Cxxv+sUbUF22s3fkJRxxoABrYT4
7KeD1bogbZ0rd1JjAHeghc6Jj8HhHeY4raI4WPTm/CmtUztBRywA6YYP4s/oFPvD3taxOTU53m9Y
i+IYpjRRuXzxJZI4IKILlVVKxBxf6f12bcSd6kh9VT633RgBK5rbFq39MmbBCMcsTv59QyRmHtNd
hOtp1tBliVHZIIFF6Ovg+BB6BEn1oDnLCa8hAihHE+u93c+mk7KGACjxgZlv//2JYQqHHPFhzrbC
3pywsZwueJcaM4diYUCZIdKq7ka6S8AwIl/ILWgjKtWHtL4yp699kcYRHWBgf01LisCkFVZEORIn
P8S3Hfmlf15xmDNKbVjKT3jjm5ZOt9z3vBNBaM9YJEtC0nv7kv7swdEL5Rmjs3s1R1bH/0gZQ9ZE
Nkr2djhbxe+cnUAKHzkAAQHpef1GOq0jE9xGIgCAZZLV87nJmCWErM1BPoE5VKIThUXUXqqibzKO
2vuniYTzoXGuKRWRo7yEKi5XKz0d5AhSI/K3mEb2Izv2vDo1qiuZiDBpaBWPgGOv5bxx+GYhrtAW
4d/uB08/kcW3YuenPhJeQSAJuvo7Uhde0D11KfEZFZ9LvgvX+PKNNeuTGe9liEZMOtM2zVjUPruh
WB1sJIGqIhGN+0BIf5S4/O8aH2nulPZcuH+OFqYffgHM3ZMGm6O/q1JW2q7IfIk5KxbvhYhtgilI
PEL0+m2iIeX+sKELrl62uBr+qb3g3tzTVcxu96264MwFYqPP6GipFWJ5SJNry2r8s1R1zEJw/jeQ
eAdelKVvumk6sJMVE1fYQYBfMm67IJYwICW1knDDViJT5dqsTO4/Z08gXJvW5JRItpcVRE8xcAYU
SDjEF2zkCRKPR9OjErPJQDLwUWxPPInZms8arKVF9udQ26EOTo5JmfOWxI+sJ3uXf8lgNY+B+F5n
wz/zIdJJAF6qbtw+16CbkLIsBtfkDFtimUaUBNK3y8TZGjzFx5m+kWnz5YiX2dXPC+/JbtQ9DQGQ
7Mcfgi9stapo2evBuxXStzEf2zeYCD2c7Cb4ArrDsKmjf7Nzgu8tWuOeHdhFJlqrBm9BD8IxFLx5
eWNzvaQOUTk2RMX+58Ip/K6ah50ToU99FKxClcox0SEzfl2ZBWIdoP1zrGh1dd2MrJEeXCaR7wvT
Y7FEqzrP6Z3E6hL8x3hyhN94IDhH5lER2zj/JCWj14QvllwwPNGuV4jdrhPFQdNmqY5pqNyYdgrc
l0NiseMe0ru4V20yR1eL+bsJlvJh9pVPUBpA5uNpSXa4u2HK4o+I4u0Ac0pT8YLN3FH00aehMD8I
RJ6SmHYbFad4LzLOpW57hbiL9LFhREa/Yl96a9UajEoTBmRFAGs/JB/KZXu/0erkC51fZJtnFjGr
RzN8C35fgr9DSOxBuXq75rXhk10tcdviSk2h1wrnMCoIZRYAgK328QWhjbWrGObIko1YdRMG91d2
/J8OdBMqvISniDd+bETDVuzggY0XaEnNuGs4J4nQQX8S4zTjSG3dINr+ASRNUyYXIz9uy94Kx4Dv
AO4HfS6IavF9I0DLGFlFQHrSpgMkPhuzuMd6rQc2yuen6ZrdRIraktaDXxw7D4TnJzHmo6qpTcME
IG+q5N19rk90Y35Tk8Bi8g3O8Fu5CYeqSelpV9ULWpytEoXnUIebEsHpIygIStx51OWxPQsIKfWm
BUNkJvMv8PeEPyayU/UuBX3AjjqSPwUsP9BF2HvYbHo4Hoj7F7VkQKRPFu+HCTQiPBtcBvUhEuOB
Tg+6LmC5nTN/9Cf2+R+7oy9L1viYIWHW3SJ0uEpcn/bGKBUYbnUIk5nuUjQrnVuR02mokJIm6iv/
muhVvvpF02tIzOs+FaH2aDbA4qGWrV6sRWSKvqneRwQFnHKx0cZ6FP7AwtdHVG3jXRpUvQKxQjS1
gc6C8rX/bTeKze1r9gi3lMUexuFJdjLzXDwe9KaeMauS+0C4FOFPydX1wnsK5q/Efs4J+DqM4Grs
RGdPkbdZU7S+WkBRpjKM6AqY6IbFZQXVCB50zGrvV1dSWpOfmbHHV1tAkIV6fnJiVIo8JGdnsTuv
ziGh0mMNCDjAudhQawAgw9NerJIWyDAcEb3HLaSmUmZ3WUlGyHARcgRUqUYslvFIaJ4Gt8CAU2bg
ZwN+QAFmQYO3J2xLyNQK3oS8mDpMg3tJhEUXB+xgA7mrflH8QFQpwYgVgxtuhDwSacJVcFhWz5B/
Fq22qcJUOrlGXdApZxMt0XDg3SKz09YAmRwVo1RAAinBb/UPjJ8lFY+f0lft+VoSQxPM/BsUxcy1
awbyw7jQkb7TcW9Y4JKp1BvSjeQVRdh7ZogC6mb5Kt3xLnYOBd74y2YPz90suXSLJVPB1nYF6ylv
T44V1Si/4Pju+6PBWEYDei7GrB28DU7yDOFz5LVunT3cJhYtjT9vamtBZRwHF5kkc2vuNrkYGmhs
FNEvXkP2lV+R+gofpEK4YNSyudXyrTYyTzkvTbaH/Mf8rdN4oeasEeJx43QAAaCClmN/ZWJuTWIO
X4NhYS1ZRfTpT1wwS/yqJSSo6u3ZxxUh1fvSAdyfQsde3SHEECuB1dvLq6apRUpQC07bFYUFnywz
e+7MAiJBCPTczNRKXX0SHEaRmbw/4aNwsEj25HHJuzURa0iOZdV7WoctfzuV9ZRDv732Kff1Gkse
+sKxvaCLe+xTCZvxXNpA/P8z5AY8mYQXGzLW/Z087nJf8Qy3bo6rNaT+Gs33E/DorKWBFeEJI46p
JZGipsX3WMW6Xv8s0Nx1LnfuTh9fpvsgoouQYwVRL8joszOU/kispxxEa1ebsCW+wQol08CjQrvP
rprA5TGKyuHysWW20D2gX+Alnc/3mWl7z+pE9JOjlzuhRJy6N0Gx9jz2SUfJdJQSix+zl/2KSUED
IALYf/SDiHftKyN/U8C9+zjR1SRbFk3ick9d5pLVHppX7hyhZ9gJLgz74DsVMHWw+/CBvBCbg0hs
1lR0hVJKOaQl3q4ZgLVAda8FN2A24uhfpydx0dE9ppGd12ZLwwfcIcWKr/9mOIs3QLC6Q7qHtsvX
uppue8Fa1QEk2QFJtEL6r0VPiJxxQk7iaNL/pVlFoBLmLYwvCOrMQOIWu8T65C20fwi6O0Hdu9oS
q21oShOkMYPtIq3mj3U59C59GYm4v//BjS96KzDvO/ZEgUsPaoZwm3AktCD43PyivigoqyMqInHJ
yyvkj6Np9ayl7FCRPbU5PnfeLDdfbacZ8/MIZVnA/lSyzH2ISVKFQWjs3l+uqd4rWlY1mOChmPM7
b1Oki20yrvp9EfjAgRwis0nsaKRVQndqLdAOCBJNkIQ0lP3uaMRDDi6WZjeV3/DNCkn3waT/p7z8
WjFPu7xsXXfnOQYs7PwQrwy7AhUhPE3p6BSWAjDJaJumA5obZ6hXmSJN3KuRsTJ0Iu4Eh39niH69
cgrH5ziiBu2G7HOyCqjZ+5/m5Yx5DQ7XRBNRLdfXgs/dIW5tMXo+r3YuD0J8Z0MoUlrPbBh0KKHg
CQQsAt+qkwzdxNdhoKGN3wpziIoCn1zRWLrEDtaJ35wtbeCFne641nZtwBJT34wa/j3P4Wwqxg27
NywW0L9wkDSorc6vhTtVObgpGBy34nXUta0cFlij7jXot8wG4oGOESJdbCmFgbL9GL1pXnuHTtcx
OVpHzM3ExxaJgYzeNBe7UC+7PjK9iuYGUP9N9FbiMMV9MkT7d9otggFlbDkDrMIUSFwR4qstHcH9
cd3RQRs/WQl5301+XyqiDUq/8VM31NPeATWwUlJeuX6ADQRzgiQZ0WkfXrcxl9bCvqpol3OrEaGB
3l3O0yHvWyjWNurqECCipoLguLLPnfv3u6RpdsWDaQyMs6IBvYxdjjdZgAsFewOF5ooNnaKVHD8Y
VbHFttmTmMYSc6BWPMsgLJC+g5vcymNVES2aEffHHprEo+dYDj4mQuzGr2d8YNF4WYI6ZpH0zvhg
Oz1yDPZ/KVwdvFK1QvutouH7okg2EAqUQOgiEjMSHUrKrjsYaTb6ZZZzq9qV58ODbMBy2DKbfMBO
3UliXoNOUi/UEfNQvmkPGY2r6UC63ah1l9fwwtKm/rCCps9+Z4BqT3KHHdBfuV048RzZaKa0eMof
1vB0aDxlCPdyqw/LagFEI4F3k6lSIi3OBojilPvCe3jvjDqTYZSNHUNdTcU5w0vXTGcgz4uQ2CEt
8XdLsTixTcoGk0VkvsbSvfZ/JG8etdg0n5yaIuoY8TcycOTwzNUTiTkojYOiXyj2Owl4H46xhzU9
dOfaHr3z+0EmQ0sJ69KNA1Bf8hTGtX7nt8VEoKiMv3QY7qfLeZ9ECqSmBPRnOe/8DEGwU4DVQMFo
rgi+S6KcuohUUjQZiPUd+xYI+QUP4fvubdkGxWKhYepdGbYQOKjmPRKvGlxtRW4Y0VLM4PcHwjXF
0wAQJMIcCY7S9E6KJ+ul3hFaL7IKp4a+6sUFl/OoFLRwHQfouSH2P7TlagGC9VDCIvfEiHRB1bXt
dUyMYozxzKswN9MsjRmENHhXyMT88Y6Uf4SMYgsP0UKpVXawf8BGwygvUmOWRjsooB1BwwmJaVtj
8/e5O7uAOZynsKPYqBL0Q3E2K9W6Sb5eHlWqw/j98EXS5Q1LsCRiZx0/hCfl5RJ/tCvXQiet8lxn
IQjndWKpJY70U05Z1OzBYUOMiZQj692QTJWsRnsPWM1m1TFTUecF/l3Oo+KnQ9uUakIqGd6RFejK
4ENxk3Xj0m4yQw+deSbBSWfsPhZIl2ZJGAdCB1j+lJjCA6LcL+lh9nj5cRJ+FuFQDXzxCMHhkR/l
xYigdfQ6/8ybFm7rSVVhwBwfFKrit1jXmqRSR0ubdjL4eYFJl1lFnUcyHLvayCCpXAauY5R8wa0P
JAkpIOWKLWjJOW3yzQk3XnMsUvI8uAUKu6T8ptb5cxrbOu3a714RqykFAOGhxmo9xm8TOpC19v6H
xZ42+fAYgNuWQIPQqtFXi/L87XuaQcZ9H4iIi9dOmOjUst0BlDhtwKkZ+kCfjGhKyi3XaM1eFiHZ
OmDcGgzeskcWRQehdXvlmnEYwr2grZWBwrGkikHzQ5JznJxJS82DykZO0eCj3BHPlLh3jCigvhTo
/jAabWOru1KmU6I2GkdImYZV8QWxb7LY1tBqGml+ZR1M3OmsexsnmCGqRAjxpG+bU1omSoxhxXE0
6lPnfr0lbJRjVJ20MqOqg2g3vaujzql80TpUQijPCv/4yC77bzAJC3dTVol8vP2kSYxujgGq7roi
FytWLqsvVEO9nsvTX9ksp8Tk/8B2IjNttXOH8HomEBqx42Le4jH7dZuHLR5sxuSQUAsYBUle6CVG
PO3rddbO0oJNpWf4RtMwAxeWCZHPUde4BXEQMPLaAIuYchQ2AaKUfxzGxt46mmgezCJRSk7enKJo
fKO8cGdQfi7ogoPjheKsiV4N2dTIRf/q43NiwfEmRkl7Qds7VXx5TQu75IjD4sz935z9DrXX76GY
EBGtY0nVNpVoQRSBi+8sWCWVCjsEMqjtArxs+ymg76WbdXr+RTZxFshvo4wD/PFKDPyOHcuGgCVH
GukW0ym4zTDigJPKJ3FdvWp8rG/1fu4BGF68YZTW8oIYzVObayJK86LMW/9/MolRZUmo2vUtFuI7
/YBzEAfuUHiYsmVU8S4t9noaXQgYHjtqeUSdtGG1/0yAruRrumnnc22Dua7/Aga+260nq/JO8Okg
fH43PPygJKB9XQuVEtzjQeUFXLUa1wKDuAtpkdEPGsRhKKVbjC3sm2gm+5nJOI1W1k7FU+wN6AMN
5B8nofJqmoAZCKRtReWiUnR+Y/Kod/HgJC8E5QzdaSflpsqkAbaMLfkBi0V157FyjvIhvBRXr9x6
esPyH3DKpjp5/2Y/TNmr9J7f4knkgQ5fqBSI7av2ms7RReDuASDkR2P6HKtdpN2opHIgRLvHzFhc
kLgYaTYx6O1Kp/pcgwfdiE5CqLHDVG5nTyOHGxIlTkFGIWBqn3fNTW5DZmm9LkPLUoNVczam4MU0
U+IdJckv+RjZ5mxJq1H32oUVvbcvgf1DB7JOflf+TysLzkMGNmh1iL68D7WsQLvZQAOhTtFOPz+p
PDzzdN4U/WKoA/7Tv4qQZ9o/Tv2U3bZOaGUI0tNvGfBO3ZtMmc0AHLEdLq9UWfJor/e1SRZE6Zeq
fy5qoBMp+VnQbjyPXsjvCvS0sgTtF1CCgBEflY114ncMTmJkAuEn2nWm2I4d1Qm+fBk5lOvgWHcs
gIxkT/BbLgD50ep6YLw+G+olezzBSYFQEkS9i2M0gD9MRP829125ifmyqkVa84dpBgBgWz8UHl4p
unhPbPQzKT0G6k4n5RVrBvFv6OmYvTwOF8QbrQA+H0WD8tR6Hs7VP+v3y0UMhzHRMF1IY62yBDrV
jT8C/LFu07pqkvczZe8CfG01DzprwOwqrnDuvK04xZEXfOrV9DD/j3ugKyN2MbeYj5M3Fm7aBjlI
t99H2EOHA0Q1pmKzJrYb+A/qAbBo6K/xZr/6sj+GAWHBHkOTk3VAzGt5Tnto3PeHcTGGl5OrAGmM
MgWIRy1q/+Zs/mVUsv6qJj0wnO7PrR1E8//zQAYIO3FmmCE1bioQzURNkf+WiiZRekkSlgFnhb0V
tuU1Anp7LClhXB+hSS/bdOKtJSHGggrcz75Vw5V2ZHjMkL6A1s1WOpy5FV0Z1NtVcg63bxBYSasP
5YD6N3A493dSk4n5kFLR20CPv1vM9c4XoLdvgk9p8sLXgKC7zwwrZbRX5DH2eOsqSP4pjhHvWGUX
p9xT4tIvBe0FxSnZ0J7eXtbXg8M5TWmRFLuJad77CBWSCHS5E9zXHmetYiltyo7Va/gOv3YvGI0F
LLw2rtfh1T270qdHxgnaB3inXfQpX0fBzyFu43kWGd9l5EsTAsAZUhQrjNmdaW8gcNhhYPwQQX04
qH5NQV8dZrTjKbMUyfnJptO+CL1YtlNJ2ShOQyx+AVUd+WoWf8CqSYDl66iMyXCgghvBAOKNnVRt
OPy/PE0aPVOFGo0m3PZh5dsXaeVETKa2S6YJ5XGnENj9YjAvz46HSdIhIhXNKVflk7cnXqfzhnrU
FJOnR3wx81kh9fV9V0+SQbncYe2024T2VGpBgCYN5ArOO+2nwsFGvQ5vbl8ozWw78JPPuCK0GMmv
C1iORMTy2clv9VhtcOJnPi3E94bWue4e0V+VkznJzDPT9egBxcwGFK5dE/sJYuBNbhMhsN22yZh0
QdNa9ekJPXdYERS3zdKPoyZABhRw3MVnj3eSZCNZgo6mx3oJ578gtWthsTNrdX0XjN64oP9okRrz
5QoEvJUQAetKTTzD36ZVvejjKPsMgFVC7GfhVgymQmzNeMp/qUjK/oBPlpgFp2k6KHqxmBLfX9x6
EgaAkK+GkYhLonbbkLw5Oj29F6OCB2m5AdWJDt3+OHe0EHyrgwPk9mqcTzQlM30s0Vl6Zw/h6RvD
ANGa79+1ZH+yngq9gNkTMaxzTJmWIP609bWH7L6XqlnI6eZZoMqg17p5v/AtDIjV/pQS4lsV/G+B
R3FGTrCYYOh1gRO/inr36sC+lBrkLOtkcoxyl0rXsndxupJ9SCpCVE4hb4hoZfd18UEQiR70+WAK
EJGhWo1Kdtzpd2aJRUtD3xNz3Ljq3BJhcJ2+m303oqUwlvV7v1/r4rYzMN7YnFHBO5yX/Pyn7tyc
DI/DT5nvEIEbWk1AvFV09O+VqeBy65ZhHdFVMZ+oJVS6/nnlrouuRwijLjZhO10qLZ0Vi1cL62vl
f7VcFhU6hPu5HHdP/+05f5CqcNO2kdlvBBFF6pMB5rcth3is5mR6Qdk9UU5TEY7EM6DLtzXhwAzq
XqAeDHyMAtP4d+7g3avZ7Vf6oJBpFufI371Z1cCmLwI0klpOOk9LQxjAECCHPdkOlGNxsvH7BOyw
wwACHPmdqvFhonZroFC59KDHM1HujDVeiP2jEIQBaty4RETZgQa6B8GlIer/hSUuHggsva6WScfJ
ZmblMwsx+oizeG3/+QdsDdz2rYV4KdajLklhFtLBf9op8DxdE+DntnrY3aVtC9izKse2Kz2mQmOM
5q3H+Fqwtnp6YHrjX+qCU1ggZBIqdKE900vUSKmc+I/HwfR4mi1WDnKmS4WzQFCVGnkgNwtZ+3Ae
KzCdp0Yu27taM6PXG9WkUttGj639HYrQl6Ut3uvv97fKpOoaLOXPBSBEWXNAD0jj7SWoWdiTQEDX
Bla6gKi+lpyEc5vr3DUa4TMFgzW3HncxBGZ0/QTSzJKJr08puKoFQNTAsi+5NN8eVb5ssNK9bK0W
4YOzLRmjZ4VlekA5MVciotj+ZLT8xEYvwKTkL/GCUX5Vn7No+w0sML92JX3ZPf4KkaVm2cDXoQju
THMudBnwOevt9mmvwSFGE97YnX1k3kQzj8xWdyCARN4NclOUpl6HmVOLc3E33xyzLb4SdFgL1iNI
08iFiY0TCTkYCjSOMhTNLNUaGShIOQGn/7L7LD8Q6U29xgqAxunnG3DV2L8nmcjuBMfc3H/UpuFn
g0RsomeKFw6ao/bKWl5GFeT4KcGTorcSlFu4V/mwe4/xCmC3vIn0v+eidOs0wb810TwyJWcOuCB8
a0JVhdx+CtubIZmbay+jPiADuTPSyTBOxxwL+f8h4U9N0TCZbTjlf6BnIB/kRXIlfix+WcORrydA
3Nm5rCYZgp5H9ySLuBspCpuYNO7ThxcCFaVPQlsz1dPqlVtiuOqVs+gSusayH295B2M5vv93uLN7
9xkFGb6fk1Fxb2I2p7jKBJ1DWooeshEwKzRgdNdsKSMjR5QOYRku5erRxqagPYp6PrGZBDowK5zg
DuIAZGYst8tL+ZnxVKYJqxPX/jIGrdu79EEgq3GT6ebQM3ofgG0CDQaApejVPYNl1l8OTddhvLqI
7QhpI4Xmt4GvkvwTHFReDNW0uVMYsN7mu3LZSUpI4eUc85cUdv2qn6zpUQVP2TpxXi9d34FUFnOh
qwKxDn65GH5H4wFohol/08gNh0pwkSiHaKv6SxRIy3LTWTVHi3jjSQJ2qPabrOJBrclwBbY+BNyJ
3EeYj4Fx89vcMHrMyXNUapfsJhashBsynoEvz7kYhsZw88A+kegasw7A58EpJ2WABHRabFed08pM
uzG7KcKKzpEq/Oda+uZ8kyz7x0pqUdlxY6YF46JLeJYISw7Ux8sbGoSm9oEUryGDhOEFiVGzU3eJ
aIYev8nd21TOIrm6KxlvJcHmlM7EJXIVm5nON+pL7cp1A+N5fEDsFcefzaDnooiEaWwsBmFz90Ap
3+wGbnJCTOTCmMkwfKdD1dnliVAx1475KRepylk+6caAu9jHwQGKrd7CvQ4n6l5aiDNQ6McFpmKc
ZhpJ1vhqv/WAo2G0TaAa9FPCaTzihGLx6NfaEFKXTzDMow7U5PWEQGfrXdoYDscTVrqj2VNY3DjF
vgEerQf/XDAs1C9a/Qsl8AVXjLHWLye8pW4+u0rmqU0cIA8QYlJiOWQm9HD9fYwRqZOBe6auIL8i
mbQG4x1M0eooGxvzjN7eEdbV/p/SaRysltxXcdXLgRXGFybNKdNhDuhbK+PLt0t5QEVcPJZjgJ3D
Vu2BwXOe0tOmYKFgRTjTsYPsDT91WV35XAfSHECoFhwqzE2GIKIfLDl2u6ZP/C8ArFvCEQc7FliG
wOPTXIx9HAyuufVNJbFH+r9goSEDF4ztTNFaOJ2M9XJQcHzqrWCLbBQsUGKXS28Us9EHpppwZ1uJ
jRRk4+wKvTp/Iq/ZemwMsctsH7cwDc42E+8ICcwVcM3KGK5xCE3bRnSIBx651XBrYukc8imMf4yX
gLGKiBibTDnzb4bOhRVvLGmonNUgvcagW+Fgq4qC5eZTUTCeNQEEYIw9jJzYDoBkDRHHygTA1DQk
dMmGmHk/0AXlgscbv6RrcHIc66qP+TygMZaoJhjjPBqFpJ/1Oxgpu810empGUy0HVwblWr6a9q/8
FS0Ffr/WzYmgZveApD/ep/5u3lbNOV4ASKdhB0DaAMDp2/nHW9BWzs5kekhK5qd1eg9qfy29m4e1
EMu2WU0+gzkiiMo896wwNc25t9S8XCc1M+82F4dNEjIazqax9ZTRD9WiZ+uWDZX/jbVWLQa4AQqi
Vy/07ssQiRrkWO3rH9RIt+TvZdYP6+9sO/TBHpJVuuUYmJsLm3uG70/DgNwWW9jVQ2D2rBR10tY8
XVXJSwy1aVa91QPRiv1fyMtubu3D+mWoeSTBGx2N1fih/ElrAO77goU+5irDRgVzngcl6pIyr4kU
rEqGsLEgXxf6OBENIejJGfDGOUr7mVmygkcqqH7006jBcmwMEYe84J+qcqjgoh1r6EPZ6lnCihW7
4w0XHkGae1o5rwfdv/zFsuSSgPPZykAo4MfMWfnA82HL6qoRI/rg6nSRhWyBZ0Q0W6RvBZMSHMDy
mdmGC7vpYWyV2e5BvOgZMairU0Q8ma94U/rTNCPA2z2bEsRHBNPqSOKDNHH7Oo2VN3+UnAhLzvz2
uOUEfr+wcEvne03E/FKkhrE2zgEe4uk7K8jX+m0fNDhLJRRQLqt9GzkI7OB8BrWMJqksV3rLQFWq
jOf+Ep8CfhKT35moSfw7jSuPEURQW4vPrVjGfs9gZSKmHipDFamEXRVtfKFaOO6APc4mG/Ayhn9T
+Xq1mqMcgkOGmMs2py3P/88liGK5LC3nmSy01RzC3pvu9Tlj/kHiFwik/An2XdN/ldDehOrzMewe
ynbrYK3lTmmUxzxO6uPYmJzvLafFXBIDKGJ+eQ1tnA62olVxr3yIKzEFpUb/EqCWK4lU2lABk5Jc
MoOAMDGNzJbRWkONT01psdbt7mDYwJyXHwc/0JUkGNXA3NSYEp7zgSXBgRhVmgzvPL4Si82U1mMl
zV4hzjopRT6xEdDel16gZqWSmcGyxV8g/VH99K5tO1Hb+C7pFAC/KGfM36uDTYy5tFQ3n0xsbA6P
T0T0vS2n0gHje1OI9T3BURYcJduN2fqbdFJ2dkWr2i71n/hG8jX0X6EXfgZDe9NErh0ciVVET3ht
JOXuG0cmpYuY1l0Jls8zXzHgH+3TEnTB7oRHAFld7mYIpSj1Nh8xMPHUd2HPCorM1XTKhCDpXJcQ
jObwqgGAW7lm5B+vJcQuCHY6hqiEtIK8pFTXP4nEdBxyUnDHRXdsbpV2KN6QLhEn4foUjUEsIc7d
sU3wDrWBKOtdg5TE/ApmIwwDDTCXZ79wxEmW1jtoQNFxdxAcADMcRcsoctKO/0iC8ou4jONayslF
fnWUAPIvTGkW17UWcmo1ksz6VtEB6zRitTZ8tGeF/g7vAkdfHthR5T/OK9tsy3DR21vaO3UKascB
KIj+NH3ECze+NbpCNsNV73X4vj4GGbzuY08GmZ3HyQLA/zg5zVxMEgq2DzVbguJlGyCFL8eVjv8J
KEbfylCG1roSRUA3D/nRWtWAWReSNhLAB1e5cmYFSFcB5ub7axyWKBlzo16d976k1RaoP7NFBPky
zTxANtookdZrE2AEtsm7jTVXL6x+lwpxIgcNh2GFMs+eW3wR/h5Nk1q/qz19mRIbEA56nka0BAMx
VL78twsM4JMZCq1GDeyMPxBIiBjj2Ib/nFCNDraj/c9DUScHWXB2e4+IZs8yatNRe0DIvo2owdV7
tLP2jbheX0hmG4+UjxO6WAngt5uumAMvXA8yyVVX+6fIeiYdawaBv8pmjh+0TkG0hvz0MXu+atFQ
z9PL6gwhDJMq12DbxeuV+1lF0ZEkeMZP4ELDSBV+VdyjtwPP+JYGtP+Czeqv8dYRm6owaTXajuyl
t5biCeFkz3wzQPpbhvjsuWby6vIEi6gf1mciG8ED3Bfn3Oxjb6198hm9wAvI1fVL6MdsFUwbLzzi
NfMrM0Unl/2duSm4XqD6fTu8CeZ2bGuUIGGYJb/DSK7MFwyhKLbhOLUF1BiSDv8rI+FsyzLlIBgS
H8wzHTIbLKYSocFAN7Ui6PaCyn7PErvnF9u6Kk1gYM2O8dUU+GLFUtSOJ+cbdPw2lUmoKNvuyH/s
AmX2Swe/QsI3b0oQh/FyVlJCiE7i4mQy5yMk2Z9BvPVEZua3Mwa5TaGrNulMEwJRLqu28wRV6kd0
CjtiQ4XRZQAtoXD9ZVZeiMPXm2bXsNe8dyK/+yZL7MYL/qJEW7MlDacnjGfKste73cGkP+7PFj3F
sJw8fil5VnpgvyHK2l7C2rSOkCVXHXE3GOMdrIBHHe84ruwduhUl1GnqEzAacOnvpWiQByfQk3/F
8Qx1EFM/hcMhbXdvWKkltltsm4duZSZeVjShb5nUbArk/c7o3YqGP8/dxG6OnHJpzGakXaVCy91c
Ws7iKCxJ8yePLkR7StP3PLCVsTeDYsGTnWAQ4+Mdh92u2AeJD2zjpHub9qOxGFZZlcjT27wlGWQQ
nNOuTM2cA0lOpc/ScMFlrAOpgTQr6sKnv61T96wLl4CpjNIj13NykLiaHmOqEd0QyvNvqc9ofzxe
+45CYD5pWLnfSYEt68bpbqlcQGAEIrqFdn93DGWfUALbPq50g0XG7Pd4xXZKIywRmdIc1oCQcu21
ymuH3M3S+mIFSP78VOTY9r1kXIH7YTJwa3QGs+g6tgHT1NdwI9ep+CcrVYzUgt18Qk+HxKuQ4Rk+
dH4lzW9zSe5forSp+EFjbWcf8rXZ/3NMhU7pSU9SKVOqpWiW4I47q3tgf9qufqQcwVqrZB8a8a+b
KkTdqXcHWJKTGQ9zAd3H1fdyAPzQS30AqGP9wsYNCBSP4ZjFegJpfEBXCU1EB46KD7CSuEBazYgn
oIIPA8xu+4rzJmccTzqY3IlrRa77nmCKbaIBcCGqs3g054xB1vIDYhQjPAE+Lj0WB5JTFNaLl3Km
Jlr8SlOfRQTCSogzDqsH4bRU9nQeIwQQNNYc1QcKJoK/h7wkGvBWQRKb3lhZGDKzTRIXMxtNBqmL
poO1/lhGf45qeU2BCy66KQUOhIBVGmcd53kGBp+cFtVcs283iwn1Wx391mENwfkqySIcDJhtc5M3
knhsh0nMt/sOC+WpiD/yTVxAIfcwoRDsAJt0qciRnRFWySQG98gr/ST55oxXDexUYsPbphWzmCne
Ro4qYbdOi/0xss3aQAXUxOnFE86lE5dslCpUVBIDtnT3bc1fTghAflevlAdoYAxpexT0Qtqpxf6z
aXhgsuutZWA9Eth9HoLgT47Bl3zjwoBYXfKQjWwdbPMWHcVymXwXvtUwTc4uIw7vRLQ9bv8S4pl7
hqb7wKDQhuegKy3hMgWNUxZbk/v2r9h0U7ohERs145tOwwH708Yx7ws61ibgYFy95bWADUJF9ZbT
xl+m8rr6Zd+5ZIVMr4WRUiXNuVJKW9H8tFGsThDHwFceYfPs9Lhl/vXZbSOTu7vPdgLdOGwWF0p7
GSrOBpYjsmIl0GLyOI0BJqZwG0e5tdf3sfawcN7J9QBAfFJD/fg2mmB35CCgqJtieRBBcfdH13z6
I5XoKYl2LiaH/WYrljWvFTsxf4LoRS1EtZgGTE/0JM6Ea5+C7Dy4rm3GWWAjjHYq7+63gNatr1iD
DqD+s7SfYMt5a1An7gmwwJpaX7Jr+c0o7ZL/bv5X4THDz7ZqlaOUnToUYGmPGkHai+R9pO/xENVw
a5lhwXxscM26DF7g+3ER2ZQ9r6QNd5bV2s2d2Q3jhMJYzkmuwRQLwGMMfjkgNr/J+PZ4RVhC1anH
9Fo/O7PZ9z4N/VnKPnKW+4tmUUzJCzg1syZqXbxfOWh46kaRhIhrohB3UkrBQxgKXe7p2mbCfHa8
NVT8ggvGxQsjRu36ksfvjj2aWCcsfEYW69HaIOYApdAAo9SVQDaZODgvf6cZu7aDTMT4UHfO1K5n
g1/Yy2huRcqAwG35SzLiZwAqJMGQGIDUmocf1Q9brpMBFJRy7IBJUZlQ5BXNzSt8yMfDqCauuRp6
9COlDaDSW37YwAHy1jzGKYNqxwTsia/1kj9UDdVkFmM7x45VF7bLi1zZcHtxieP/ALYSscwlYNqh
BhDW1YEgdu0SqYmC7A+4PfvLHJRb0ZBH+PyQp/On9mWBH8+qxOC9iVkQQnzsL/sPsQF9CB3tdiyo
ABnTHDtPM+nwCQ5JNlnN4bGUjTYmhbNt1GnsXFnfHwdaO6zmZgAeR2FGQQxi1ZdRhjsqo66bPLbK
Qp6/DoXMij7dzuCTT/pePlEtPEScrrvOOCz4mDyh/NWX1vkTSnjxalxfd26LBNFiOmdfhPJHcjDa
sg6xlAhf+JIsTUi43pGTSdFuuV2JFpwEw/pdeg2zCX2PPqTsdtodzpjKJAxlObrW/a6eKF9g+UMG
9en3KONHnrqUb5digwZ44VsKuoyFAnp3dh7Y7eQdZVMirRzabNWc113mnIHtZug6PSIXBLY9BkpV
VbKVuq/5E7TrDWcSJ8qaY8pBA1G2kh8szKuFrh+dKVly035OqkOEC/J86heTzB9NxR7OlmADjUCZ
xIxwA0bGu57iLk39L8hhAVzFRVpr4CNNe6lx3pKPV5i0w2pVwuRo8OgQYs3IaSkkZ6Ez3spI+mvb
eBkP55arc4kT5dtMCgZrp6mfi2hpEcr14Z24H7fF03zqDO3Z/kN/tV8WiT/101muDS9n2SRs0ec0
ll0/iF44XAHqQtXtbK8s+AIbDyiGepFjaqGy4eMP3xeb8KCyifNIzMOL2upSMiu+qPfAdqD1zaqt
hr9iHR+UIRtQPQs3vjog8WhGSsOzEiFak1PEvc0+A3DigF/n/7wn63I6I9/KXHPGCpVR/vU9XkBy
Iu2+hBwrj8ADT4iDLkwdW/UFvy1qyByMfyxf0aKHmC8uyk1la7WfAOgAnrPjCADdEariQjaaiIZa
PblTo8IWr5Gb+QHFYg7Rb+GRCMo4dspqdMp14zoKuPN6xNVGsABvgnX2CkDjRf1k4XbriZrVXG38
4JoDxBPX3/UzQIMkl5+vCOG1YOCbzW0fE4DNNhcHl+cPqEr0KaZ3lvAJN/PDipVxpwl5Jt066Zl/
2jY835rBu2P9WfhPwtnRQ7PR07Wqyw/WbN4li2WTU6bo0E0lOmsjBhFtyGX3yEoSK2Ih060E+l6k
y6b60gCB8p8e/SJtLuXefD/+gD7Uu/aiS7EgfPXD6XG8q4kcvJ9my9wkZpxvSqPe+AGcfyOLFLT2
XkeIOMao1S6sK89opfBsagwkLxYd6iaEjTp7WZ1cRSJBSiomjmj1kHhhaW8dZICWGOBjKbItD1tt
6qL1QybBTymo1kwuylmqhwYy0xoXQuOMbfAdXBpUeLpwz7TgfeO34PL4ViDfbhWq+nvZUoj6nMvA
aGg2zdw7ImNRk93/zw3iIj76IFsrRzWEJCzIdMEJ/TfS9G+hHZEgkxjCiwnCvrKJ5y1/vQfvoOL/
TIQqXsocLm6CsUBvI6fu8VJaCQ/cxkL0JMbdnDDZ/LqQD+1o7FXdly9aYoa0rzt3yifTPXLvOSw/
ck0TtnLidvQgQRVkH8q/n4b2kwPfZ7q6qGZKt12mOWqN/V9Du2clbO+cgArpf3fm2HUUTKWPTjn/
SyI5MOBC7x0nkAyLIbS95drBUe0MpEjKl54XKn4vaNYVz7yw2+v54JOowMtu9TLsozMvhkGJc1L8
uXD45druNR2H1KTEgPqiTZZRTBQX4w+9ezKdfWACg21w+/g/C3JeY0LNAywQjIcWQDZi90QNgAS8
om/tQ7OKHpvztIb2QP6Wqo470655e4VZPUQqMm/Gz9N+wbZ/ZLzCBF1McnOyll3Duz7ep/r/jnHw
uX8PPv4JKmeGaXmV8JROHCu2UhiHY6HsSJX1Npyw/7yqgUA00YkCch1Oh0zlB5lRe7qpWZsK1KnP
YGpLK1RqoV2ZYg7f/ruecIMjRV5rSg7PWj1gfrXkxmcAXlM343Gv7AipT7D5FmZzXFpsnnfcKrg4
9kRWW9EZ8uzTcSodQjgfrpMD3T9jinXva8f2U/C08IofNQhHyM9A6a6YWEXJSUz+x9cy2NXahua0
aBO6bhGOdUzVXsrKuSzX8z9zogK5Vx26dJf0z8yF9ICYNII/jBHoOOS/iLR0Qp/qB4CIuh2EOdY/
7452vmle7PMRD8h9Y6WiM4hAUzl7It8pE41Z6ajseQZfuS8xx8mfaYvWGfg5o6RYrKu/7ivORXn3
NCrZRZ7z0W+KRYWehiWNiz9ZuSmAZMHazMzfcIOgfVWBCIPxKN/+wS5XwgvMXYhIYvFJ+L8zUXBw
7pXbHfrxuQ4uzNxrKTLE0EmEIpKs2fB8ZM235HOip5lpMsQi6e4Cw4Jr93E75cm2CmCxDOTeuSKl
d3tz5bgTBF0yj6c4Wr4fOc1wtYasEul+/m0BCMV/q2+Rc1OOZXfJS0HTbkGyznQdxGFsgvCy+da7
plhYVT4nkhFWoiCafcVnXxmlmLlPzqDz1X+6CXIkqV8IpOhv0qWV1wRTK0qH0KpdqyB0zCYcF6CP
mBzdEri2MLXm8duujxjrv4I0wp6lyoQXUB9ZWCVdIBmZ3mwPtq1NV/TrFd37zJnBcOFscgRalMFd
ygwXhAtKhr+syIxudiisVOMARDue7fh6LNtc1QlV6hGBOJQ+gSpUGQPJ+wn8IvwgGsR1jrQ5d4vG
tONqIXnzbaaiGTwGpWL3KTRkHC7JDYa1tEF2v0lEf5m+FKOIwvp4Y9GltgGvnbOik1uQjFST/1Ly
pTte0H7GlbQY37MCL9Rdv03R7Lxdw7xsb43zdGUCGFtm6HX/c8kgXDzRiuFxGMnRTmoBn3Qx/agR
CYryaaBqt+H5RiaW86MmWLBxoQyK4b3NRlvWcQEiM7gX5Qcm4aX5qhbdbVnMkhnFc//lzG8UIa1N
ql3oWZ4x8K0GIZLOi2I7UhHJ96/uAYyGyHhhU8jOb1C1MImXXbdCw/aD1YtDEx97s6HV+XqO245H
c59RZfasdI2dQIcOnBpqYeyeRtLBv9DqNUsNZTnOy2S14Dxj/KFlwJdyUQ5fa21Az6odFJeMaaoD
+rCaHBnNJnOzLhukMafnZf5NSULFXyMns9OXH0G9tbmEHzbhdO51y3hXPei8NV5SpYlK2Ltdx29o
fk/fzGXHeD91PKG5uuRMkWDrFRYL9v2Vk8ubmwAX+zJvs70Axm1VEXuSJIC+rpwky+45jeUc6KxV
L4FokrpDq8TqfaiNmBMOKCIc8irDsf8ulxoxp+GgJSHx9QkY4HJlrZUtOq3sjZUJppUitf7FH5xm
IiI/1YhH1Xcunv9+mspduDQZch3BQhWlvLVCJzev0AylqSo0sRSEaEbUUJ0zFCEFpI9nd4bEPdLm
momAuYDAejPp0u4b1/YpR8ds2u3U9efrZv3LpBkjZkoaP6zzsZqKnCd/GXO0/UD+s60eU58jOc67
fZw9HAwJaZ0nnzaYGXYLS0wtaJwBeLLiHLQgoE4zkbAFOWySZL/4j4/BSsA1ktyeIo+QbiD0LovY
DGPMj6WCpV6tNuK4pX8+8KHtXMK/49arnyT8Rh3SA+OsW0TfwO1xtKNVbGLO3Z3KdU7bjFmiaNCF
BkTXbLII4Xg4AopRrdDK6nrl9e0vFWglHSCpBHUZG7496FxpNnyBcb3K3Hd0Hz5ZY7aQ8+nZmZWV
KgENWvEivH5P7qyGTiAvGWVx7Ij8gH/RPSTYJR10/v59FZLiSxDkz31u7qjqJoeX+Bz1BE7lPqye
8F0K1GgJJd7ipaPQpyc1PibRNXlzacgevYoWf3AaDGFt2yHpyzYCOp1VNMFG71wClHrh8/6bYZlw
nNZY0R6NLPSowaw2+U9WejYpDET2+e7sy+cEdcK5+DcZZZYKLBL28/U20x2D6Jlz5c8WgfzxeK1n
UCDQgjSU0St9JR7xXKKgYQu2v3cXkh3jQwY5jPw5FHhRH6WfiA83LTMMDMHj5H17ywIt6qJ8//Zw
riR46WByCtsKo1heCGYrf2g2No8jK1Ny4RgqZp8xR1YYeSR72cFv22gpmlLK7HnSIi8Dqqv84pCt
OeOK/xb2l1qoZ6v5ANLq1XYEXsvgDd3S5H2fUmr0YYmHOS4rkIK2KHT0JFzjU+mwcODStRLLa30a
awTwsohLfi1jVk8sxLoudiSlY4mnfuWR0EDbO7CbS4CF0xB55hk/X6NYJqAMhuX5dIvHzj72DsdY
+KWRZGK6BHIghVoY7ybUosRFO7xHuq8n2wQmnEeVkBZa9tOP7yKEBpM1he55mDmiCwiG0IP/NNyS
gf+H/nvXv3qKPqzAwHDJ9kKleyfxTEm+5/+KkiQilU5zJhbc2THu1An9Af0I8AqraFzlp+/3jRhi
sQu90LA/HzKMIuMTqzTG5H3DCbBew/jBIrE7lx5zO0KaYiFprMYVzeYE4srTWcHPP/pkUfN86ZZd
aeCCiHPeHgW8pWYeTjKu0zV9JjStlN2brAFkWWYb7T0H88wLkGvVIrw13yE01Bpl0uym4MzGunUd
XwQlYD8AAuxh4rHZp73O4o+TidYf/O5AIbVmsyQVgf1s0J3iinbC/Ij+/lVM/Tp77D0qwTV1vXgA
8zBou2hHVRkTaaGL8I37iSsU1lIW+cK5/uAxbYzDMttKMOmCeAGjUgg2F5aI2phAwpo8xJihhMwf
2PypQQiizKyU8RYjHAjeMubUYIJ7GjbXCWufKusLCMh5+1vt0LTHbOCqIu2+bStSfmZL3CG+3otZ
DM3P//Iv+H2JAOXJS6vaZjhv+j11gN7Dz4BfjyD40uiABZJV9w8evMeo0Wk/b0Zatu68xgFotEzA
FOkuQv5Vkguz0aDuh3SiThbsGEV0Tho+UsvdYm2CwrbLttwSKhz5g3AOAgE6+/rTOR8y9V7/wZS8
IgWP5EWyaEF/MrTEQWhwO8PWwIu9z8fjmucBjIePKnM79GRPC8XTwCG5sCBpYucs5f0bxk2alVp1
JTgo/9eYT8qBfOMELMu59RvBM60uftxUnXtKQAYeuw0bZCuQHDG3eDlYgOqBqUHAPcHWPtWtvUHj
VdJtOq14k7HcncKuCjKDnTdb9IJgxKKI4j5zx87GocwgPcyvGVs87KK0EjSnypTEZakIaHQHPfRL
vxPHog8lzwbdQL6mYoOArG21Zoa8Lf+ioNl+GUpxapb2kw6nNtKCqvQbNGtvv4L88KLRVyNz6yEA
VbVDqaUjwMHXZLi6EUPY70OUATzPYOn3tDHuNjT/gkaLS47hu+cQ9vOZt5gHjlY0zUEOHINOpW+d
UnsIDhj+8laRFC9/T8FiItXDyJeGKnKDRD8lNQbhn9XHoImsuS3BzbbZE4lRx4f/h36baOV/uFjA
j6FgTwQNGRIShqMxhrTpB7BCwIQ9MIxCdpd6tfVjlzH+M1V7N+Vq2gSu7plCn0hpyYMULCutnc4h
0BuxURrOpxNho62DAaub2b+a/QLjysJx4gew5JVDDteGzBOfa3Le2hoYJkogdZv22N/YYruo1NwQ
cdT/cBUc2dpRfFqsliwE2j2XxoAPhHmT1LBQlupxF+j5wIfcuCDUwNRPGXyfL8sOvfx0nXUs5TWt
RUEP1ztmOQcnPpITBXCE10d61lWApz7UGWgKK00/l+ATdLvfHDSiKhbEVffp89vuwahQjQ7KkcR3
JS9Fnr3piEIWLregp/M797KmPUomS8p1g4xK8GHHu6BQafIgaaPk+Xr12uQ7VtCuxsFEi1T8Pvla
NkGYocAtT/1nbtiSmQmVbV1UKw7BO65x1hhwdg0cZ77eYDnHSPXaIyDVREBmGu3Y8g1iGC2LiL8V
h1bz57jfWK4pCm9RirHVeBK01NDZF/fGVbGkAUXj0LtLkRkxdiHisXU2m5bBymA3Cygb4h2N5sjl
IHEsfC5hgcTRaiXgJ+8jDsfmgZ6B10MUsroHUdbNHpBaL0LoWq0R9Rn7W7GWwIHz+yvDB1Ayix/9
U9+jcV3m2gpdf6QTcutSwcSji5MopnlSAQOzbYA6zoh06VSm9HD7Yo/OIK7dwvsNJbic8c2sifdq
u0ii3zEETtV1WtOM0SYb84/SGHpMrTdDl8FLbirfRXXzhMqVPrEslK/yZC4ivugYP1YDttRAvZgc
gPzDVZxImUSrODjOTR7GTAUijsqdw4HmH2HYjuj/fw52rWAGeBk5ijKwsn/nzdoY/pDBzQV/H7XY
ppWsW3lY/KMO37q4A2mLOZj1Txalp7nC/iQXDAbV3xlNhheSxc6/zjm03Lcnoql/m9sFvn0s/4dc
dAGoBj+aPgJt/FEyH8NznLEBARkgPCTZlU2X2femUBX6qCS8lHVA1mUQaZ6QW7meyD0OXHzyVrwf
/QWL7DKi4+D9E89PorbO0qq3o0/WtCByiXPXExCXnJVxzFp0TsWlq/AOtQ5qToS0WWIDhWOB1S/D
ln4Cl3qfpg9DJUtr+U8pWC4DIF6VU5FH0aoZlZ38WixgGBE1JPXoAHQ5CM/op+MxnTgKSHCHiqCx
9/AfpX9fHLlaUXpPZ7Xe+KnQdwti0O5Jk9H7JFnWwwU94svstn5bhT6+D3wxmwk1LM7pf1IoZOsI
wwSQWV2Ii3PS/WFFgBSiJM54tbWE8WRYI01j09AHxK6+s3nHrrv6mQXYqWJecQLKqY797pD75TtV
ybQuGg69DMKdCFN59YH8i+3paeoHJSrjv6edw1r3gI5M9alPmwGXwHJqrskCKYK2ZQFs1CuekxbC
y5CGcMwzh9mW+wGRWCfGMpna5NdxhNChUKlHZiLRZZGE9ahuYJhXb44c7xpA8VBAf4vf4o0aNmZD
cpvq0OD9UWgdjlGrQZm6DxT+Oxso38Cx/zswlnqrP18apd1BHEZv2vlZluHpjJMKv2fhcUkC25fy
hqUHeaAax51ojrpenOseqyRAE0B51rs/LZRFeBAlRA679fW9XQn/01LHxRbEWbBrfqZImpWYMgMG
D9jSG02TGxmkl329EQSD3wA2jSwFsZUckP/GIuAoo0yqow0R8uPqfTG+muEknIMuQbZ77V07iOyy
qpPB6VePRRp8+69lzuScllulOvZ5qEMnWgqNnmWDwG1Co0dfp7Y1wc6UEzOG6d9ww/jtBGWtrmY+
uJq3I7Ti0q7ZJhsV8+Zy2k4J2pKXjXJ0r87kBCM/vBqAplmHjW8am3FZPziV+ZpjcKzltqcrAphW
la0P353wnhOS/Cue8kHFOsonuyTxOsFmCYmd6roa7Tu9wRjdUqJjYGCIA3vbOfQg2mhIHrIrpb1R
RQNbRNDtwNWhUzXo+59W/ImBM60Tl3+8/eUtk3Eva8vCim7aGK+AzLZ9P+3Hg5FnHtBbyPWLdzN7
nEhYkGXe+aIV8ORNf91t3fjeCo744n0qCBrMwib6tqGkWqXoxLeLt3+Gp2K7fCljeaYcjnKE7Zut
DZllGAIPs1+hLFiUEPax10zZNRlC6HfUEedWSArmVkeHtljy55lQpTBjbvAWTCPDFO6X6yXNhEHT
+KBtXDps9b5Tzmr89TREuLkU2QW6RGyMyQS9FbvViuwOLkld7ChxPmhm2zBmbYODt5Gmo9iT9cxh
YlTKRU4UYftQq3eRRG6AywLl6d3iTsuJpz4aA0+L1/MVrqHBzDJ0T/7s46OiED07+cmGsjp2iMJv
E1pY91Y73+HjhdXwms+zZKq9HkwSZ9ZxnRPShBPF3ki6sIccovIFA4HufRfa63ovYBB5phlDs3nx
HDs2iYpbDSz4ESVArFHt4XpU0nSuLKfArCdZJAj2w7FRhPiEhYT+HxQBY9iCOu5uekxkb+zCsaKG
b4Q1UklsPJhRzpFHPk2xavRFUfJi+fPiRVzyS3HvHgu+ZSvf4KspGzPRgB3xouXWSHth9eUkobG+
12kd83YLhvDkmbNx3CJSA9Patx8cSc3PAGwSE7+Mplc47g04+qVxZ+Qc8YO21aJ4d0FgOvs+yuEX
yLBnS1PoTLZtnLHYg+NF9/j3Dx23/BrvGuqxUSUZcBTldp2aaTDlY0G2nNpkgiKA6KL8aXisxPEp
ztPwniaf/jgMDOs0437krF7otz8QH2m6TD7CeGIynwA2wa2qim3sZZiGa3nEWcLhb4IgeyzMZPwy
5fH9MM1xWALEbn0m/tXN7SLukBKE2flXT6jHJ2nO6FgdXt7Grf0WLm/qH3QVa+5lTkmRIv6/TrNE
6ouCfA4oyk4s5QsjC4lJckxR+q+qAGr4xui0bswQt65uxdflWtCxvB52KOa990SprIh0XN8WBOzX
W4M8T6Z33pqREB4k6WJbjHHpEPN85ZFRw9DfWJr2oBbAW52PzSpBu+H9oyyEW7ut4S0G05UA4+Ub
qgy9Qk+RBOSz2axXCmg3R5lbGepzTigaWwAg2/xc2mkHI8tAmo2f00xBckqRNM2HL+iZ+idiNhOr
Ml3ta/9LeB3diy96qdrYr8jW98SlayQKsmCj2lhlaAUmDJPEeJYl/b2NgpXIKPkGBsws4k1rF/LT
uMJKwFmo+jfb9OXimpKyrPcuYEWXbbErEyp5pGFZpngCZbWcErYPuoIooFg/GOPoHZfEf2g40qXj
mXXJ8wK8xfSdKYOO3Inc9RLxTOeyuENpuyt2la0k8O7sqrl0rVNoNLBiWxMhW0qxipl51VBSbXwH
sGaiIefgEnPLYQWkR3HOPrvuqPPTSaiORso7y61EpK0GbpoY2rZeuffV1Z6zjDlbnA6AKSVSh7KW
IvXjUT9oFd0eTdTlpsS3n8KFnVtazO8IlgXq29Mo21GPDnGpGiDIZ9EEXDIKFsDb7dJZomAuN9i5
4LwE31oPgzqUAFJ3Dd8vKgD8OwvTlv4FvnWe5mM6/8v7U9NZx39nhWTzov/rWe3MAIx+FS/rH1Xa
L5t1ngk60HzrAzL2z7RW5B/YC2Il9qZJC8cRX3qaftWX1njysRLNhb+VCyeX05o3BN2nHu3DKdQB
f3r656t/8s7XRKb0prj1jxK/IfVkTcGpfqQYNMUQh1I+flXNeO64xqx/BK+Q98Y+IHEDrh9fODiB
xA8LfUeIo2qg5eO5ZjOl8MVKo2lHlWNUJvORntUttG+UH9+RApRsMymR9UZNUXLHkBFhCBcw4njQ
lpeMKns30a56bIkGBK01pz91lxzJLj6tsc2nTwoDXVbaS4yhcMYMymiZjMHjrzOPrEFQ5EOldvJo
xfTrC8cdFRx0NjBTStmDpGl6UNEWchr2959gzNMMzZ/hUFO6Nvv69JF24Ib9GU/Mk6T8x8j+MEGw
dzSKUaD0cFIMMhuNG/DURNY8SJ/EVOTH0nZz+z2ND6OSUVBjsAMYkZWKS6cce3nNjJxhsFRWnMs/
1HG7snP0R665tyDXuzIzS6cUqCH33uuaann+AdakUY1HTqjbBIHOb84UQ/hbGQFOsWJx+tdc7Pi1
aWdDJCe+6U09if1prF/zV4j6ve9CGQOsRVqZoTPZSLm0K+M96rmJkP5tguEqj+a5JX99bVufDgn1
l5imFH7aar55XcHZNQqC9hDcmLOGWDnCB10NM1E47y4HWg66RNsHTLRHveOOvovRqo0omMwWMjNe
Kvk5hzn3Xm4kmNNoWUBWCWVDzPxqprEzoc4yvFHUzNQCqCnM2XFIlfASqTxG3D4kKYcEJMKfle+Q
EMDT1ZfcsK1CQ2NZa/wat70euLJmhex74iStMpUK+RAMsIdIi0pVtBDny+CeCKOzfXiEwnJFsjZD
QiVZKzDznGZu4vqpGBitielHILMifA+Do9ykh9LMM/BeprM3Cbxu0JNHh/aTjEL8Rhe+qjkiyheM
VUaQX331FUJvGSbWpQRuHTYjpNYPCGBXrF0jzubkZabLXCzEEA95FTGxZ+wZKA/CdsuvbS0FoqSl
tp4rNWUDstmrfb10MrS22okrplyrXN4bz6Kv5pWHgkEDB2JwH6Y2eirM+pYHEwIOI0c5W6C9gm6J
4pgb1ReZOnI5joi/3+ltlSz4XJb8PKEk7NA7ysAN6+fuy/YBHjwkIzOgfJCHL19IO8M7LKaY5jM4
yW3JWyQbPke+mvx1lruCfAjn4h4UUSk1HemKgsORjgHPVovKXDGvINT9Oofv1JL5dM01Enh2ltuj
AOp5G7M9QKC0zsRylF6Mcnu44isb3tnT8Akzu8hkI1AjxndgRVpZdxDidTp4OwhicJuYX1j5uTTC
X4YT2td6zw==
`protect end_protected

